module alu4_2 (
	i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, 
	i_8_, i_9_, i_10_, i_11_, i_12_, i_13_, o_0_, o_1_, o_2_, o_3_, 
	o_4_, o_5_, o_6_, o_7_);

input i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, i_8_, i_9_, i_10_, i_11_, i_12_, i_13_;

output o_0_, o_1_, o_2_, o_3_, o_4_, o_5_, o_6_, o_7_;

wire n1, n2, n3, n5, n8, n9, n10, n11, n12, n14, n16, n18, n19, n21, n20, n24, n23, n26, n33, n31, n32, n30, n35, n36, n34, n38, n39, n40, n37, n42, n43, n41, n46, n45, n44, n50, n47, n53, n51, n57, n56, n61, n58, n63, n62, n65, n69, n73, n74, n72, n77, n78, n76, n79, n83, n84, n85, n87, n88, n82, n91, n90, n89, n93, n94, n92, n96, n95, n99, n98, n97, n104, n101, n102, n100, n106, n107, n108, n105, n110, n111, n109, n113, n114, n112, n116, n118, n115, n119, n124, n125, n123, n127, n132, n133, n134, n135, n136, n138, n139, n131, n140, n146, n147, n144, n145, n143, n149, n151, n148, n152, n157, n158, n159, n160, n161, n162, n156, n166, n167, n164, n165, n163, n168, n170, n171, n169, n173, n174, n172, n175, n178, n179, n177, n181, n180, n185, n186, n182, n190, n191, n188, n189, n187, n193, n194, n192, n196, n197, n195, n201, n202, n199, n198, n206, n204, n205, n203, n210, n211, n209, n207, n214, n212, n217, n216, n215, n218, n220, n219, n223, n222, n221, n224, n226, n225, n229, n230, n228, n227, n231, n234, n233, n232, n236, n235, n238, n239, n237, n242, n241, n240, n243, n248, n249, n247, n246, n250, n251, n252, n255, n253, n257, n256, n259, n260, n258, n261, n264, n268, n267, n271, n270, n276, n275, n280, n279, n287, n283, n288, n296, n292, n297, n302, n303, n301, n306, n307, n304, n308, n311, n309, n313, n312, n315, n314, n317, n318, n316, n320, n323, n322, n326, n324, n327, n330, n331, n328, n332, n333, n335, n334, n339, n337, n338, n336, n341, n340, n344, n342, n346, n345, n349, n348, n347, n352, n351, n350, n353, n354, n357, n362, n360, n365, n364, n363, n367, n366, n370, n371, n372, n369, n376, n373, n377, n380, n381, n379, n384, n383, n382, n387, n388, n389, n390, n391, n385, n393, n394, n392, n396, n397, n398, n395, n399, n402, n403, n401, n406, n404, n409, n408, n411, n412, n415, n410, n417, n416, n421, n419, n424, n422, n426, n425, n428, n429, n433, n430, n434, n437, n445, n448, n451, n449, n455, n453, n454, n452, n457, n458, n460, n461, n462, n456, n463, n467, n468, n466, n470, n471, n469, n472, n476, n479, n478, n481, n480, n485, n483, n482, n486, n488, n487, n490, n489, n492, n493, n491, n494, n495, n497, n496, n499, n498, n500, n502, n506, n504, n508, n507, n513, n514, n511, n517, n518, n515, n519, n521, n520, n522, n524, n523, n525, n529, n528, n532, n533, n534, n535, n537, n538, n531, n539, n541, n540, n542, n543, n548, n547, n551, n552, n550, n553, n556, n554, n557, n559, n558, n561, n565, n564, n568, n567, n570, n569, n572, n573, n571, n575, n574, n578, n577, n584, n582, n581, n585, n588, n591, n592, n596, n597, n599, n600, n601, n602, n604, n603, n607, n608, n606, n609, n610, n612, n613, n614, n615, n616, n617, n611, n620, n619, n618, n622, n621, n624, n623, n626, n625, n628, n629, n630, n631, n627, n633, n632, n635, n637, n638, n639, n636, n641, n640, n647, n646, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n677, n680, n681, n682, n683, n684, n685, n686, n687, n688, n690, n691, n692, n693, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n707, n708, n709, n710, n711, n712, n713, n714, n716, n717, n718, n719, n722, n720, n725, n723, n727, n726, n728, n730, n733, n732, n736, n734, n738, n740, n742, n743, n744, n745, n746, n747, n748, n749, n751, n750, n752, n753, n754, n755, n757, n758, n759, n761, n762, n764, n763, n766, n765, n768, n767, n769, n770, n772, n771, n773, n775, n777, n776, n779, n778, n781, n780, n782, n785, n783, n788, n789, n790, n791, n792, n794, n796, n795, n797, n799, n798, n802, n803, n805, n804, n806, n808, n807, n810, n809, n812, n813, n814, n816, n818, n817, n819, n821, n822, n820, n823, n824, n825, n826, n827, n828, n829, n830, n832, n834, n833, n835, n838, n837, n841, n840, n844, n843, n845, n846, n847, n848, n849, n851, n852, n854, n857, n856, n858, n863, n862, n861, n867, n865, n870, n869, n871, n873, n872, n874, n876, n878, n879, n882, n884, n886, n885, n890, n891, n893, n895, n894, n896, n898, n899, n901, n900, n903, n902, n904, n905, n906, n908, n909, n910, n911, n912, n914, n915, n916, n920, n921, n922, n923, n927, n930, n932, n933, n934, n935, n937, n941, n940, n942, n943, n944, n945, n946, n951;

assign o_0_ = ( (~ n19) ) ;
 assign o_1_ = ( (~ n636) ) ;
 assign o_2_ = ( (~ n627) ) ;
 assign o_3_ = ( (~ n611) ) ;
 assign o_4_ = ( (~ n18) ) ;
 assign o_5_ = ( n10 ) | ( n11 ) | ( n12 ) | ( n14 ) | ( n16 ) | ( (~ n817) ) | ( (~ n819) ) | ( (~ n820) ) ;
 assign o_6_ = ( (~ n9) ) ;
 assign o_7_ = ( n1 ) | ( n2 ) | ( n3 ) | ( n5 ) | ( n8 ) | ( (~ n717) ) | ( (~ n791) ) | ( (~ n792) ) ;
 assign n1 = ( (~ i_9_)  &  (~ n177) ) | ( (~ i_9_)  &  n180 ) | ( (~ i_9_)  &  n182 ) ;
 assign n2 = ( n50  &  n522  &  i_9_ ) ;
 assign n3 = ( (~ i_5_)  &  (~ n776) ) | ( (~ i_5_)  &  (~ n264)  &  n296 ) ;
 assign n5 = ( i_9_  &  n47 ) | ( i_9_  &  (~ n771) ) | ( i_9_  &  (~ n773) ) ;
 assign n8 = ( n267 ) | ( n270 ) | ( n275 ) | ( n279 ) | ( n283 ) | ( n288 ) | ( (~ n782) ) | ( (~ n783) ) ;
 assign n9 = ( (~ i_2_)  &  n332  &  n333 ) | ( n328  &  n332  &  n333 ) ;
 assign n10 = ( i_11_  &  (~ n807) ) | ( i_11_  &  (~ n317)  &  n445 ) ;
 assign n11 = ( n448  &  n326  &  i_2_ ) ;
 assign n12 = ( (~ n61)  &  (~ n666) ) ;
 assign n14 = ( (~ n701)  &  (~ n806) ) | ( (~ i_13_)  &  (~ n666)  &  (~ n701) ) ;
 assign n16 = ( (~ i_4_)  &  (~ n804) ) | ( (~ i_4_)  &  (~ n42)  &  (~ n334) ) ;
 assign n18 = ( (~ n574)  &  (~ n577)  &  (~ n585)  &  n596  &  n597  &  n599  &  n600  &  n601 ) ;
 assign n19 = ( (~ i_0_)  &  (~ n23)  &  n641 ) | ( (~ n23)  &  n641  &  n640 ) ;
 assign n21 = ( (~ i_1_) ) | ( (~ i_3_) ) ;
 assign n20 = ( (~ i_5_) ) | ( n21 ) ;
 assign n24 = ( (~ i_8_)  &  i_10_ ) ;
 assign n23 = ( i_3_  &  n24 ) | ( i_3_  &  (~ n542) ) ;
 assign n26 = ( (~ i_6_)  &  (~ n53) ) | ( (~ i_10_)  &  (~ n53) ) ;
 assign n33 = ( n39  &  n655 ) | ( n125  &  n655 ) | ( n39  &  n35 ) | ( n125  &  n35 ) ;
 assign n31 = ( i_1_ ) | ( n557 ) ;
 assign n32 = ( i_11_ ) | ( n118 ) ;
 assign n30 = ( n33  &  n31 ) | ( n33  &  n32 ) ;
 assign n35 = ( i_12_ ) | ( n118 ) ;
 assign n36 = ( i_0_ ) | ( n247 ) ;
 assign n34 = ( n31  &  i_11_ ) | ( n35  &  i_11_ ) | ( n31  &  n36 ) | ( n35  &  n36 ) ;
 assign n38 = ( (~ i_6_) ) | ( i_7_ ) ;
 assign n39 = ( i_0_ ) | ( n233 ) ;
 assign n40 = ( i_0_ ) | ( i_1_ ) | ( (~ i_2_) ) ;
 assign n37 = ( n38  &  i_6_ ) | ( n39  &  i_6_ ) | ( n38  &  n40 ) | ( n39  &  n40 ) ;
 assign n42 = ( (~ i_3_) ) | ( n247 ) ;
 assign n43 = ( (~ i_3_) ) | ( n557 ) ;
 assign n41 = ( (~ i_5_)  &  (~ i_6_) ) | ( (~ i_6_)  &  n42 ) | ( (~ i_5_)  &  n43 ) | ( n42  &  n43 ) ;
 assign n46 = ( i_0_ ) | ( n45 ) ;
 assign n45 = ( i_3_ ) | ( i_2_ ) ;
 assign n44 = ( (~ i_5_)  &  n46 ) | ( n46  &  n45 ) ;
 assign n50 = ( (~ i_12_)  &  i_13_ ) ;
 assign n47 = ( n50  &  (~ n763) ) | ( i_8_  &  n50  &  (~ n471) ) ;
 assign n53 = ( i_6_  &  n653 ) ;
 assign n51 = ( (~ n174)  &  (~ n765) ) | ( n53  &  (~ n174)  &  (~ n497) ) ;
 assign n57 = ( i_6_  &  i_7_ ) | ( n46  &  i_7_ ) | ( i_6_  &  n223 ) | ( n46  &  n223 ) ;
 assign n56 = ( n57  &  i_8_ ) | ( n57  &  n39 ) ;
 assign n61 = ( (~ i_12_) ) | ( n118 ) ;
 assign n58 = ( (~ i_1_)  &  (~ i_6_) ) | ( (~ i_6_)  &  n61 ) | ( (~ i_1_)  &  (~ n421) ) | ( n61  &  (~ n421) ) ;
 assign n63 = ( (~ i_1_)  &  i_6_ ) ;
 assign n62 = ( (~ i_0_)  &  (~ i_1_) ) | ( (~ i_0_)  &  i_5_ ) | ( (~ i_1_)  &  n63 ) | ( i_5_  &  n63 ) ;
 assign n65 = ( (~ i_9_)  &  (~ n73)  &  (~ n364) ) ;
 assign n69 = ( i_3_  &  n65 ) | ( i_3_  &  (~ n61)  &  (~ n99) ) ;
 assign n73 = ( (~ i_11_) ) | ( n118 ) ;
 assign n74 = ( i_8_ ) | ( i_6_ ) ;
 assign n72 = ( (~ i_2_) ) | ( i_9_ ) | ( n73 ) | ( n74 ) ;
 assign n77 = ( (~ i_0_) ) | ( n45 ) ;
 assign n78 = ( (~ i_0_) ) | ( n216 ) ;
 assign n76 = ( i_6_  &  i_7_ ) | ( n77  &  i_7_ ) | ( i_6_  &  n78 ) | ( n77  &  n78 ) ;
 assign n79 = ( i_0_  &  n69 ) | ( i_0_  &  (~ n72) ) | ( i_0_  &  (~ n778) ) ;
 assign n83 = ( i_3_ ) | ( (~ i_11_) ) | ( n39 ) | ( (~ n421) ) ;
 assign n84 = ( (~ i_3_) ) | ( i_9_ ) | ( n118 ) | ( n497 ) ;
 assign n85 = ( (~ i_5_) ) | ( n58 ) | ( n197 ) ;
 assign n87 = ( n196 ) | ( (~ n406) ) | ( n650 ) ;
 assign n88 = ( n656 ) | ( n73 ) | ( i_9_ ) | ( n62 ) ;
 assign n82 = ( (~ n79)  &  n83  &  n84  &  n85  &  n87  &  n88 ) ;
 assign n91 = ( n144  &  n98 ) | ( n655  &  n98 ) | ( n144  &  n173 ) | ( n655  &  n173 ) ;
 assign n90 = ( (~ i_6_) ) | ( n656 ) ;
 assign n89 = ( n91  &  n90 ) | ( n91  &  n31 ) ;
 assign n93 = ( (~ n53)  &  (~ n101) ) | ( (~ n101)  &  n173 ) | ( (~ n53)  &  n655 ) | ( n173  &  n655 ) ;
 assign n94 = ( n654  &  n652 ) | ( n497  &  n652 ) | ( n654  &  n31 ) | ( n497  &  n31 ) ;
 assign n92 = ( n93  &  n94 ) ;
 assign n96 = ( n36  &  (~ n102) ) | ( (~ n102)  &  n108 ) | ( n36  &  n144 ) | ( n108  &  n144 ) ;
 assign n95 = ( n96  &  n40 ) | ( n96  &  n90 ) ;
 assign n99 = ( (~ i_6_) ) | ( n326 ) ;
 assign n98 = ( (~ i_6_) ) | ( (~ i_7_) ) | ( i_8_ ) ;
 assign n97 = ( n99  &  n95  &  n98 ) | ( n99  &  n95  &  n39 ) ;
 assign n104 = ( i_5_  &  n453 ) ;
 assign n101 = ( (~ i_6_)  &  n653 ) ;
 assign n102 = ( (~ i_0_)  &  i_1_  &  (~ i_2_) ) ;
 assign n100 = ( n104  &  (~ n757) ) | ( n104  &  n101  &  n102 ) ;
 assign n106 = ( i_11_ ) | ( (~ n185) ) ;
 assign n107 = ( i_10_ ) | ( n364 ) ;
 assign n108 = ( i_6_ ) | ( n656 ) ;
 assign n105 = ( n106  &  n108 ) | ( n107  &  n108 ) | ( n106  &  n32 ) | ( n107  &  n32 ) ;
 assign n110 = ( i_12_ ) | ( n114 ) ;
 assign n111 = ( i_11_ ) | ( n114 ) ;
 assign n109 = ( (~ n53)  &  n98 ) | ( n98  &  n110 ) | ( (~ n53)  &  n111 ) | ( n110  &  n111 ) ;
 assign n113 = ( i_11_ ) | ( i_12_ ) ;
 assign n114 = ( i_9_ ) | ( i_13_ ) ;
 assign n112 = ( n113 ) | ( n114 ) | ( i_3_ ) | ( i_10_ ) ;
 assign n116 = ( i_5_ ) | ( n376 ) ;
 assign n118 = ( i_10_ ) | ( i_13_ ) ;
 assign n115 = ( (~ i_10_)  &  n118 ) | ( n116  &  n118 ) | ( (~ i_10_)  &  (~ n181) ) | ( n116  &  (~ n181) ) ;
 assign n119 = ( i_13_  &  (~ n749) ) | ( i_13_  &  (~ n684)  &  (~ n685) ) ;
 assign n124 = ( i_5_ ) | ( n649 ) ;
 assign n125 = ( i_12_ ) | ( (~ n406) ) ;
 assign n123 = ( n124  &  (~ n181) ) | ( n125  &  (~ n181) ) | ( n124  &  (~ n268) ) | ( n125  &  (~ n268) ) ;
 assign n127 = ( n50  &  (~ n748) ) | ( (~ i_3_)  &  (~ i_11_)  &  n50 ) ;
 assign n132 = ( n652 ) | ( n692 ) | ( n693 ) ;
 assign n133 = ( n144 ) | ( n690 ) | ( n691 ) ;
 assign n134 = ( n220 ) | ( (~ n287) ) | ( n656 ) ;
 assign n135 = ( (~ n53) ) | ( (~ n104) ) | ( (~ n421) ) ;
 assign n136 = ( n108 ) | ( (~ n406) ) | ( n565 ) ;
 assign n138 = ( n98 ) | ( (~ n383) ) | ( n658 ) ;
 assign n139 = ( n123  &  n681 ) | ( n654  &  n681 ) | ( n123  &  n683 ) | ( n654  &  n683 ) ;
 assign n131 = ( (~ n127)  &  n132  &  n133  &  n134  &  n135  &  n136  &  n138  &  n139 ) ;
 assign n140 = ( n90  &  n108 ) | ( n108  &  (~ n499) ) | ( n90  &  (~ n522) ) | ( (~ n499)  &  (~ n522) ) ;
 assign n146 = ( n164  &  n188 ) | ( n688  &  n188 ) | ( n164  &  n165 ) | ( n688  &  n165 ) ;
 assign n147 = ( n746  &  n747  &  n682 ) | ( n746  &  n747  &  n687 ) ;
 assign n144 = ( (~ i_7_) ) | ( n74 ) ;
 assign n145 = ( (~ n104) ) | ( (~ n268) ) ;
 assign n143 = ( n146  &  n147  &  n144 ) | ( n146  &  n147  &  n145 ) ;
 assign n149 = ( (~ i_0_) ) | ( (~ i_1_) ) | ( i_4_ ) ;
 assign n151 = ( i_4_ ) | ( n557 ) ;
 assign n148 = ( (~ i_6_)  &  (~ i_7_) ) | ( (~ i_6_)  &  n149 ) | ( (~ i_7_)  &  n151 ) | ( n149  &  n151 ) ;
 assign n152 = ( i_2_  &  (~ i_8_)  &  (~ n241)  &  (~ n658) ) ;
 assign n157 = ( n683 ) | ( n686 ) ;
 assign n158 = ( n108 ) | ( n174 ) | ( n179 ) ;
 assign n159 = ( (~ n101) ) | ( n692 ) | ( n693 ) ;
 assign n160 = ( n90 ) | ( n690 ) | ( n691 ) ;
 assign n161 = ( n220  &  n217 ) | ( n688  &  n217 ) | ( n220  &  n165 ) | ( n688  &  n165 ) ;
 assign n162 = ( n684  &  n144 ) | ( n687  &  n144 ) | ( n684  &  n680 ) | ( n687  &  n680 ) ;
 assign n156 = ( n157  &  n158  &  n159  &  n160  &  n161  &  n162 ) ;
 assign n166 = ( n98  &  n188 ) | ( n680  &  n188 ) | ( n98  &  n688 ) | ( n680  &  n688 ) ;
 assign n167 = ( n744  &  n745  &  n682 ) | ( n744  &  n745  &  n686 ) ;
 assign n164 = ( (~ i_5_) ) | ( n222 ) ;
 assign n165 = ( (~ n50) ) | ( (~ n315) ) ;
 assign n163 = ( n166  &  n167  &  n164 ) | ( n166  &  n167  &  n165 ) ;
 assign n168 = ( n90  &  n98 ) | ( n90  &  (~ n499) ) | ( n98  &  (~ n522) ) | ( (~ n499)  &  (~ n522) ) ;
 assign n170 = ( n189  &  n681 ) | ( n220  &  n681 ) | ( n189  &  n684 ) | ( n220  &  n684 ) ;
 assign n171 = ( n742  &  n743  &  n677 ) | ( n742  &  n743  &  n683 ) ;
 assign n169 = ( n170  &  n171  &  n90 ) | ( n170  &  n171  &  n145 ) ;
 assign n173 = ( (~ i_0_) ) | ( n233 ) ;
 assign n174 = ( (~ i_5_) ) | ( n376 ) ;
 assign n172 = ( n173 ) | ( n144 ) | ( n174 ) ;
 assign n175 = ( n98 ) | ( (~ n102) ) | ( n116 ) ;
 assign n178 = ( i_2_ ) | ( n376 ) ;
 assign n179 = ( (~ i_10_) ) | ( (~ n383) ) ;
 assign n177 = ( (~ i_5_) ) | ( n90 ) | ( n178 ) | ( n179 ) ;
 assign n181 = ( i_3_  &  i_4_  &  (~ i_5_) ) ;
 assign n180 = ( i_1_  &  (~ i_7_)  &  (~ n73)  &  n181 ) ;
 assign n185 = ( (~ i_12_)  &  (~ i_13_) ) ;
 assign n186 = ( i_10_  &  i_11_ ) ;
 assign n182 = ( (~ n172)  &  n185  &  n186 ) | ( (~ n175)  &  n185  &  n186 ) ;
 assign n190 = ( n675  &  n677 ) | ( n164  &  n677 ) | ( n675  &  n682 ) | ( n164  &  n682 ) ;
 assign n191 = ( n108  &  (~ n559) ) | ( n145  &  (~ n559) ) | ( n108  &  n681 ) | ( n145  &  n681 ) ;
 assign n188 = ( i_3_ ) | ( n673 ) ;
 assign n189 = ( (~ n50) ) | ( (~ n548) ) ;
 assign n187 = ( n190  &  n191  &  n188 ) | ( n190  &  n191  &  n189 ) ;
 assign n193 = ( n188  &  (~ n559) ) | ( (~ n559)  &  n675 ) | ( n188  &  n677 ) | ( n675  &  n677 ) ;
 assign n194 = ( n90  &  n681 ) | ( n680  &  n681 ) | ( n90  &  n682 ) | ( n680  &  n682 ) ;
 assign n192 = ( n193  &  n194  &  n189 ) | ( n193  &  n194  &  n164 ) ;
 assign n196 = ( i_10_ ) | ( n656 ) ;
 assign n197 = ( (~ i_8_) ) | ( n326 ) ;
 assign n195 = ( n196  &  n197 ) ;
 assign n201 = ( n195  &  (~ n578) ) | ( (~ n578)  &  (~ n582) ) | ( n195  &  n738 ) | ( (~ n582)  &  n738 ) ;
 assign n202 = ( n740  &  n667 ) | ( n740  &  n39 ) ;
 assign n199 = ( n107  &  n99 ) ;
 assign n198 = ( n201  &  n202  &  n199 ) | ( n201  &  n202  &  (~ n481) ) ;
 assign n206 = ( n107  &  (~ n409) ) | ( (~ n409)  &  n565 ) | ( n107  &  n669 ) | ( n565  &  n669 ) ;
 assign n204 = ( i_8_ ) | ( n668 ) ;
 assign n205 = ( (~ i_4_) ) | ( n233 ) ;
 assign n203 = ( n206  &  n204 ) | ( n206  &  n205 ) ;
 assign n210 = ( n402  &  (~ n670) ) | ( n402  &  n671 ) | ( (~ n670)  &  n672 ) | ( n671  &  n672 ) ;
 assign n211 = ( n99  &  n205 ) | ( (~ n104)  &  n205 ) | ( n99  &  n602 ) | ( (~ n104)  &  n602 ) ;
 assign n209 = ( (~ i_5_) ) | ( n326 ) ;
 assign n207 = ( n210  &  n211  &  n209 ) | ( n210  &  n211  &  (~ n409) ) ;
 assign n214 = ( n654  &  n652 ) | ( n173  &  n652 ) | ( n654  &  n655 ) | ( n173  &  n655 ) ;
 assign n212 = ( n31  &  n214 ) | ( (~ n101)  &  n214 ) ;
 assign n217 = ( i_3_ ) | ( n236 ) ;
 assign n216 = ( i_1_ ) | ( i_3_ ) ;
 assign n215 = ( (~ i_5_)  &  n217 ) | ( n217  &  n216 ) ;
 assign n218 = ( i_0_ ) | ( i_3_ ) | ( (~ i_6_) ) ;
 assign n220 = ( i_3_ ) | ( n650 ) ;
 assign n219 = ( n220  &  i_5_ ) | ( n220  &  n216 ) ;
 assign n223 = ( i_0_ ) | ( n216 ) ;
 assign n222 = ( i_3_ ) | ( i_6_ ) ;
 assign n221 = ( n223  &  n219  &  i_0_ ) | ( n223  &  n219  &  n222 ) ;
 assign n224 = ( (~ i_0_) ) | ( (~ i_3_) ) | ( (~ i_6_) ) ;
 assign n226 = ( i_1_  &  (~ i_6_) ) ;
 assign n225 = ( i_2_  &  (~ i_7_) ) | ( (~ i_6_)  &  (~ i_7_) ) | ( i_2_  &  n226 ) | ( (~ i_6_)  &  n226 ) ;
 assign n229 = ( i_6_ ) | ( n945 ) | ( n651 ) ;
 assign n230 = ( i_1_ ) | ( i_7_ ) | ( n651 ) ;
 assign n228 = ( i_11_ ) | ( n542 ) ;
 assign n227 = ( n229  &  n230  &  n225 ) | ( n229  &  n230  &  n228 ) ;
 assign n231 = ( i_5_ ) | ( n45 ) ;
 assign n234 = ( i_2_ ) | ( n650 ) ;
 assign n233 = ( i_1_ ) | ( i_2_ ) ;
 assign n232 = ( n234  &  i_5_ ) | ( n234  &  n233 ) ;
 assign n236 = ( (~ i_5_) ) | ( (~ i_6_) ) ;
 assign n235 = ( i_2_  &  (~ i_5_) ) | ( i_2_  &  n233 ) | ( (~ i_5_)  &  n236 ) | ( n233  &  n236 ) ;
 assign n238 = ( (~ i_2_)  &  (~ i_5_) ) | ( (~ i_5_)  &  n236 ) | ( (~ i_2_)  &  n247 ) | ( n236  &  n247 ) ;
 assign n239 = ( (~ i_6_) ) | ( n557 ) ;
 assign n237 = ( n238  &  n239 ) ;
 assign n242 = ( (~ i_1_) ) | ( (~ i_5_) ) | ( (~ i_7_) ) ;
 assign n241 = ( (~ i_1_)  &  (~ i_6_) ) ;
 assign n240 = ( (~ i_0_)  &  n242 ) | ( (~ i_7_)  &  n242 ) | ( n242  &  n241 ) ;
 assign n243 = ( i_10_  &  (~ n237)  &  (~ n542) ) | ( i_10_  &  (~ n240)  &  (~ n542) ) ;
 assign n248 = ( (~ i_2_) ) | ( n650 ) ;
 assign n249 = ( i_6_ ) | ( n557 ) ;
 assign n247 = ( (~ i_1_) ) | ( (~ i_2_) ) ;
 assign n246 = ( n248  &  n249  &  i_5_ ) | ( n248  &  n249  &  n247 ) ;
 assign n250 = ( n246  &  i_7_ ) | ( n246  &  n62 ) ;
 assign n251 = ( (~ i_0_)  &  (~ i_1_) ) | ( (~ i_0_)  &  i_5_ ) | ( (~ i_1_)  &  i_6_ ) | ( i_5_  &  i_6_ ) ;
 assign n252 = ( i_7_  &  i_6_ ) | ( n149  &  i_6_ ) | ( i_7_  &  n151 ) | ( n149  &  n151 ) ;
 assign n255 = ( (~ i_2_) ) | ( (~ i_8_) ) | ( n63 ) | ( n124 ) ;
 assign n253 = ( n252  &  n255 ) | ( n255  &  (~ n604) ) ;
 assign n257 = ( n36  &  (~ n102) ) | ( (~ n53)  &  (~ n102) ) | ( n36  &  n652 ) | ( (~ n53)  &  n652 ) ;
 assign n256 = ( n40  &  n257 ) | ( (~ n101)  &  n257 ) ;
 assign n259 = ( (~ i_4_) ) | ( n247 ) ;
 assign n260 = ( (~ i_4_) ) | ( n696 ) ;
 assign n258 = ( i_8_  &  i_6_ ) | ( n259  &  i_6_ ) | ( i_8_  &  n260 ) | ( n259  &  n260 ) ;
 assign n261 = ( i_4_  &  (~ n775) ) | ( (~ i_1_)  &  i_4_  &  (~ n196) ) ;
 assign n264 = ( i_6_  &  (~ n261) ) | ( i_10_  &  (~ n261) ) | ( (~ n261)  &  (~ n670) ) ;
 assign n268 = ( (~ i_9_)  &  n406 ) ;
 assign n267 = ( n181  &  (~ n256)  &  n268 ) ;
 assign n271 = ( (~ i_10_)  &  (~ i_13_)  &  n506 ) ;
 assign n270 = ( (~ n124)  &  (~ n720) ) | ( (~ n89)  &  (~ n124)  &  n271 ) ;
 assign n276 = ( (~ i_3_)  &  (~ i_8_) ) ;
 assign n275 = ( n152  &  (~ n659) ) | ( (~ n148)  &  n276  &  (~ n659) ) ;
 assign n280 = ( (~ i_9_)  &  (~ i_13_)  &  n479 ) ;
 assign n279 = ( (~ n658)  &  (~ n723) ) | ( (~ n212)  &  n280  &  (~ n658) ) ;
 assign n287 = ( (~ i_11_)  &  i_13_ ) ;
 assign n283 = ( n287  &  (~ n726) ) | ( (~ n248)  &  n287  &  (~ n662) ) ;
 assign n288 = ( n50  &  (~ n730) ) | ( n50  &  (~ n732) ) | ( n50  &  (~ n734) ) ;
 assign n296 = ( n406  &  i_12_ ) ;
 assign n292 = ( (~ n198)  &  n296 ) | ( (~ n203)  &  n296 ) | ( (~ n207)  &  n296 ) ;
 assign n297 = ( (~ n61)  &  (~ n759) ) | ( (~ n61)  &  (~ n761) ) | ( (~ n61)  &  (~ n762) ) ;
 assign n302 = ( i_4_  &  (~ n287) ) | ( (~ i_8_)  &  (~ n287) ) | ( (~ n287)  &  (~ n506) ) ;
 assign n303 = ( (~ i_3_)  &  (~ n406) ) | ( n228  &  (~ n406) ) | ( (~ i_3_)  &  n667 ) | ( n228  &  n667 ) ;
 assign n301 = ( n125  &  n302  &  n303 ) | ( n302  &  n303  &  (~ n604) ) ;
 assign n306 = ( (~ i_7_) ) | ( i_10_ ) ;
 assign n307 = ( i_4_ ) | ( (~ n479) ) ;
 assign n304 = ( (~ i_7_)  &  n306 ) | ( n306  &  n307 ) | ( (~ i_7_)  &  (~ n384) ) | ( n307  &  (~ n384) ) ;
 assign n308 = ( i_7_  &  n24 ) ;
 assign n311 = ( i_8_  &  (~ n308) ) | ( n304  &  (~ n308) ) | ( i_8_  &  n698 ) | ( n304  &  n698 ) ;
 assign n309 = ( i_7_  &  n311  &  (~ n915) ) | ( n301  &  n311  &  (~ n915) ) ;
 assign n313 = ( (~ i_7_) ) | ( (~ i_9_) ) ;
 assign n312 = ( i_7_  &  n313 ) | ( (~ i_10_)  &  n313 ) ;
 assign n315 = ( (~ i_7_)  &  i_8_  &  i_10_ ) ;
 assign n314 = ( i_12_  &  n315 ) | ( i_12_  &  (~ n685) ) ;
 assign n317 = ( (~ i_10_) ) | ( n656 ) ;
 assign n318 = ( i_8_ ) | ( n313 ) ;
 assign n316 = ( (~ i_11_)  &  (~ n314) ) | ( (~ n314)  &  n317  &  n318 ) ;
 assign n320 = ( n110  &  n111 ) | ( n110  &  (~ n276) ) | ( n111  &  (~ n604) ) | ( (~ n276)  &  (~ n604) ) ;
 assign n323 = ( (~ i_4_) ) | ( n118 ) ;
 assign n322 = ( (~ i_8_)  &  n323 ) | ( n35  &  n323 ) ;
 assign n326 = ( (~ i_7_) ) | ( i_9_ ) ;
 assign n324 = ( (~ i_4_) ) | ( n326 ) ;
 assign n327 = ( i_13_  &  i_7_ ) | ( n324  &  i_7_ ) | ( i_13_  &  n322 ) | ( n324  &  n322 ) ;
 assign n330 = ( n339  &  i_4_ ) | ( n339  &  n316 ) ;
 assign n331 = ( n695  &  n794  &  i_3_ ) | ( n695  &  n794  &  n327 ) ;
 assign n328 = ( (~ i_13_)  &  n330  &  n331 ) | ( n312  &  n330  &  n331 ) ;
 assign n332 = ( n685  &  (~ n946) ) | ( n698  &  (~ n946) ) ;
 assign n333 = ( n802  &  n803  &  i_2_ ) | ( n802  &  n803  &  n309 ) ;
 assign n335 = ( (~ i_6_) ) | ( (~ i_9_) ) ;
 assign n334 = ( i_6_  &  n335 ) | ( (~ i_10_)  &  n335 ) ;
 assign n339 = ( n398 ) | ( n118 ) ;
 assign n337 = ( (~ i_7_)  &  n657 ) | ( i_7_  &  n920 ) | ( n657  &  n920 ) ;
 assign n338 = ( i_2_ ) | ( i_13_ ) ;
 assign n336 = ( n339  &  n337 ) | ( n339  &  n338 ) ;
 assign n341 = ( i_10_ ) | ( i_7_ ) ;
 assign n340 = ( i_11_ ) | ( n341 ) ;
 assign n344 = ( i_11_ ) | ( i_13_ ) ;
 assign n342 = ( (~ n185)  &  n196 ) | ( n196  &  n340 ) | ( (~ n185)  &  n344 ) | ( n340  &  n344 ) ;
 assign n346 = ( i_8_ ) | ( n326 ) ;
 assign n345 = ( (~ n185)  &  n344 ) | ( n197  &  n344 ) | ( (~ n185)  &  n346 ) | ( n197  &  n346 ) ;
 assign n349 = ( (~ i_6_)  &  n342 ) | ( i_6_  &  n345 ) | ( n342  &  n345 ) ;
 assign n348 = ( (~ i_8_)  &  n657 ) | ( i_8_  &  n920 ) | ( n657  &  n920 ) ;
 assign n347 = ( n349  &  i_13_ ) | ( n349  &  n348 ) ;
 assign n352 = ( i_7_  &  n704 ) | ( (~ i_7_)  &  n705 ) | ( n704  &  n705 ) ;
 assign n351 = ( i_7_ ) | ( n542 ) ;
 assign n350 = ( (~ i_6_)  &  n352 ) | ( (~ i_11_)  &  n352 ) | ( n352  &  n351 ) ;
 assign n353 = ( n340  &  i_12_ ) | ( n340  &  n306 ) ;
 assign n354 = ( (~ i_2_)  &  i_6_  &  (~ n951) ) | ( (~ i_2_)  &  (~ n353)  &  (~ n951) ) ;
 assign n357 = ( (~ i_4_)  &  (~ n354) ) | ( (~ n354)  &  (~ n719) ) ;
 assign n362 = ( i_2_ ) | ( (~ i_4_) ) | ( n738 ) ;
 assign n360 = ( n199  &  n357  &  n362 ) | ( n357  &  n362  &  (~ n453) ) ;
 assign n365 = ( (~ i_7_) ) | ( n335 ) ;
 assign n364 = ( i_6_ ) | ( i_7_ ) ;
 assign n363 = ( (~ i_10_)  &  n365 ) | ( (~ i_9_)  &  n365  &  n364 ) ;
 assign n367 = ( (~ i_6_)  &  (~ n317) ) | ( i_6_  &  (~ n674) ) | ( (~ n317)  &  (~ n674) ) ;
 assign n366 = ( (~ i_4_)  &  (~ n718) ) | ( (~ i_4_)  &  i_11_  &  n367 ) ;
 assign n370 = ( (~ i_3_)  &  n347 ) | ( i_3_  &  n350 ) | ( n347  &  n350 ) ;
 assign n371 = ( i_13_  &  n334 ) | ( (~ i_13_)  &  n360 ) | ( n334  &  n360 ) ;
 assign n372 = ( (~ i_2_)  &  (~ n366)  &  n816 ) | ( n363  &  (~ n366)  &  n816 ) ;
 assign n369 = ( n370  &  n336  &  n371  &  n372 ) ;
 assign n376 = ( (~ i_3_) ) | ( i_4_ ) ;
 assign n373 = ( n338  &  n376 ) | ( n376  &  (~ n479) ) | ( n338  &  (~ n506) ) | ( (~ n479)  &  (~ n506) ) ;
 assign n377 = ( i_3_  &  (~ i_4_) ) | ( (~ i_4_)  &  n125 ) | ( i_3_  &  (~ n406) ) | ( n125  &  (~ n406) ) ;
 assign n380 = ( (~ i_3_)  &  (~ n287) ) | ( (~ n287)  &  (~ n506) ) | ( (~ n287)  &  n685 ) ;
 assign n381 = ( (~ i_2_)  &  (~ i_7_) ) | ( (~ i_2_)  &  n373 ) | ( (~ i_7_)  &  n664 ) | ( n373  &  n664 ) ;
 assign n379 = ( n380  &  n381  &  n377 ) | ( n380  &  n381  &  n197 ) ;
 assign n384 = ( i_4_  &  n421 ) ;
 assign n383 = ( (~ i_11_)  &  n421 ) ;
 assign n382 = ( (~ n196)  &  n384 ) | ( (~ i_3_)  &  (~ n196)  &  n383 ) ;
 assign n387 = ( (~ i_2_) ) | ( i_7_ ) | ( (~ n499) ) ;
 assign n388 = ( (~ n383) ) | ( n702 ) ;
 assign n389 = ( (~ i_3_) ) | ( n317 ) | ( (~ n479) ) ;
 assign n390 = ( (~ i_2_) ) | ( i_8_ ) | ( n307 ) ;
 assign n391 = ( i_7_  &  (~ n50) ) | ( (~ n50)  &  n376 ) | ( (~ n50)  &  (~ n479) ) ;
 assign n385 = ( (~ n382)  &  n387  &  n388  &  n389  &  n390  &  n391 ) ;
 assign n393 = ( i_11_ ) | ( (~ n626) ) | ( n697 ) | ( (~ n702) ) ;
 assign n394 = ( (~ i_6_)  &  n379 ) | ( i_6_  &  n385 ) | ( n379  &  n385 ) ;
 assign n392 = ( n393  &  n394  &  n90 ) | ( n393  &  n394  &  n307 ) ;
 assign n396 = ( (~ i_11_) ) | ( n648 ) ;
 assign n397 = ( (~ n185) ) | ( (~ n604) ) ;
 assign n398 = ( (~ i_4_) ) | ( i_9_ ) ;
 assign n395 = ( n396  &  n398 ) | ( n397  &  n398 ) | ( n396  &  n73 ) | ( n397  &  n73 ) ;
 assign n399 = ( i_3_  &  i_12_  &  (~ n651) ) ;
 assign n402 = ( i_1_ ) | ( n45 ) ;
 assign n403 = ( (~ i_11_) ) | ( (~ n185) ) ;
 assign n401 = ( n205  &  n402 ) | ( (~ n268)  &  n402 ) | ( n205  &  n403 ) | ( (~ n268)  &  n403 ) ;
 assign n406 = ( i_11_  &  (~ i_13_) ) ;
 assign n404 = ( i_4_  &  (~ n809) ) | ( i_4_  &  (~ n402)  &  n406 ) ;
 assign n409 = ( (~ i_1_)  &  n453 ) ;
 assign n408 = ( i_7_  &  n399 ) | ( i_7_  &  n409  &  n268 ) ;
 assign n411 = ( (~ i_8_)  &  n921 ) | ( n401  &  n921 ) ;
 assign n412 = ( n500  &  n228 ) | ( n433  &  n228 ) | ( n500  &  n700 ) | ( n433  &  n700 ) ;
 assign n415 = ( (~ n24)  &  n651 ) | ( n42  &  n651 ) | ( (~ n24)  &  n696 ) | ( n42  &  n696 ) ;
 assign n410 = ( n395  &  (~ n404)  &  (~ n408)  &  n411  &  n412  &  n415 ) ;
 assign n417 = ( (~ i_2_) ) | ( i_12_ ) ;
 assign n416 = ( (~ i_8_)  &  n417 ) | ( n42  &  n417 ) | ( (~ i_8_)  &  (~ n488) ) | ( n42  &  (~ n488) ) ;
 assign n421 = ( i_12_  &  (~ i_13_) ) ;
 assign n419 = ( n421  &  (~ n813) ) | ( i_4_  &  (~ n402)  &  n421 ) ;
 assign n424 = ( i_8_  &  n814 ) | ( (~ n499)  &  n814 ) | ( n700  &  n814 ) ;
 assign n422 = ( (~ i_9_)  &  (~ n419)  &  n424 ) | ( n416  &  (~ n419)  &  n424 ) ;
 assign n426 = ( (~ i_8_) ) | ( i_9_ ) ;
 assign n425 = ( n205  &  (~ n312) ) | ( n205  &  (~ n409) ) | ( (~ n312)  &  n426 ) | ( (~ n409)  &  n426 ) ;
 assign n428 = ( i_10_ ) | ( n74 ) ;
 assign n429 = ( (~ i_6_) ) | ( n426 ) ;
 assign n433 = ( (~ i_1_) ) | ( n376 ) ;
 assign n430 = ( (~ n308)  &  n365 ) | ( (~ n308)  &  n433 ) | ( n365  &  (~ n445) ) | ( n433  &  (~ n445) ) ;
 assign n434 = ( (~ i_4_)  &  (~ n713) ) | ( i_13_  &  (~ n713) ) | ( (~ n626)  &  (~ n713) ) ;
 assign n437 = ( i_6_  &  (~ n647) ) | ( i_11_  &  (~ n647) ) ;
 assign n445 = ( i_3_  &  n226 ) ;
 assign n448 = ( (~ i_6_)  &  n522 ) ;
 assign n451 = ( (~ i_9_) ) | ( (~ i_11_) ) ;
 assign n449 = ( (~ i_12_) ) | ( n451 ) ;
 assign n455 = ( (~ i_4_) ) | ( n114 ) ;
 assign n453 = ( (~ i_3_)  &  i_4_ ) ;
 assign n454 = ( (~ i_9_) ) | ( (~ i_12_) ) ;
 assign n452 = ( n455  &  n453 ) | ( n455  &  n454 ) ;
 assign n457 = ( i_9_  &  (~ i_13_) ) | ( (~ i_9_)  &  n712 ) | ( (~ i_13_)  &  n712 ) ;
 assign n458 = ( i_3_ ) | ( n109 ) ;
 assign n460 = ( i_2_ ) | ( n99 ) | ( (~ n185) ) ;
 assign n461 = ( (~ i_1_)  &  n449 ) | ( n335  &  n449 ) | ( (~ i_1_)  &  (~ n488) ) | ( n335  &  (~ n488) ) ;
 assign n462 = ( i_4_  &  (~ n53) ) | ( (~ n53)  &  n449 ) | ( i_4_  &  n452 ) | ( n449  &  n452 ) ;
 assign n456 = ( n457  &  n458  &  n460  &  n461  &  n462  &  (~ n927) ) ;
 assign n463 = ( (~ i_4_)  &  (~ n703) ) | ( (~ i_4_)  &  (~ n108)  &  n186 ) ;
 assign n467 = ( (~ i_10_)  &  (~ n923) ) | ( (~ i_13_)  &  (~ n226)  &  (~ n923) ) ;
 assign n468 = ( n108  &  (~ n463)  &  n852 ) | ( n323  &  (~ n463)  &  n852 ) ;
 assign n466 = ( n467  &  n468  &  i_3_ ) | ( n467  &  n468  &  n105 ) ;
 assign n470 = ( i_7_ ) | ( n650 ) ;
 assign n471 = ( (~ i_7_) ) | ( n236 ) ;
 assign n469 = ( n470  &  n114 ) | ( n118  &  n114 ) | ( n470  &  n471 ) | ( n118  &  n471 ) ;
 assign n472 = ( (~ i_2_)  &  (~ n851) ) | ( (~ i_2_)  &  (~ n323)  &  (~ n552) ) ;
 assign n476 = ( i_3_  &  (~ i_8_)  &  (~ n36) ) ;
 assign n479 = ( i_11_  &  (~ i_12_) ) ;
 assign n478 = ( (~ i_0_)  &  i_2_  &  i_10_  &  n479 ) ;
 assign n481 = ( (~ i_0_)  &  n453 ) ;
 assign n480 = ( (~ i_6_)  &  n478 ) | ( (~ i_6_)  &  (~ n61)  &  n481 ) ;
 assign n485 = ( n36  &  n39 ) | ( n36  &  (~ n383) ) | ( n39  &  (~ n499) ) | ( (~ n383)  &  (~ n499) ) ;
 assign n483 = ( i_0_ ) | ( n21 ) ;
 assign n482 = ( n307  &  (~ n480)  &  n485 ) | ( (~ n480)  &  n485  &  n483 ) ;
 assign n486 = ( (~ i_6_)  &  (~ i_7_) ) | ( (~ i_7_)  &  n77 ) | ( (~ i_6_)  &  n78 ) | ( n77  &  n78 ) ;
 assign n488 = ( i_8_  &  i_3_ ) ;
 assign n487 = ( i_7_  &  (~ n497) ) | ( n488  &  (~ n497) ) ;
 assign n490 = ( (~ i_3_)  &  (~ n271) ) | ( i_3_  &  n691 ) | ( (~ n271)  &  n691 ) ;
 assign n489 = ( (~ i_4_)  &  n307  &  n490 ) | ( n61  &  n307  &  n490 ) ;
 assign n492 = ( (~ i_12_) ) | ( n712 ) ;
 assign n493 = ( i_2_  &  (~ n50) ) | ( (~ n50)  &  n107 ) | ( (~ n50)  &  (~ n383) ) ;
 assign n491 = ( n492  &  n493  &  n489 ) | ( n492  &  n493  &  n108 ) ;
 assign n494 = ( (~ i_7_) ) | ( n451 ) ;
 assign n495 = ( n226  &  i_2_ ) | ( n197  &  i_2_ ) | ( n226  &  n429 ) | ( n197  &  n429 ) ;
 assign n497 = ( (~ i_1_) ) | ( n557 ) ;
 assign n496 = ( (~ i_6_)  &  (~ i_8_) ) | ( (~ i_8_)  &  n43 ) | ( (~ i_6_)  &  n497 ) | ( n43  &  n497 ) ;
 assign n499 = ( i_10_  &  (~ i_12_) ) ;
 assign n498 = ( n476  &  n499 ) | ( (~ i_0_)  &  n226  &  n499 ) ;
 assign n500 = ( i_7_ ) | ( (~ n186) ) ;
 assign n502 = ( n186  &  (~ n901) ) | ( (~ i_8_)  &  n186  &  (~ n497) ) ;
 assign n506 = ( (~ i_11_)  &  i_12_ ) ;
 assign n504 = ( n506  &  (~ n835) ) | ( i_8_  &  (~ n36)  &  n506 ) ;
 assign n508 = ( (~ i_0_) ) | ( n21 ) ;
 assign n507 = ( n500  &  (~ n502)  &  (~ n504) ) | ( (~ n502)  &  (~ n504)  &  n508 ) ;
 assign n513 = ( (~ i_1_)  &  (~ n287) ) | ( i_11_  &  (~ n287) ) | ( (~ n287)  &  n335 ) ;
 assign n514 = ( (~ n53)  &  n834 ) | ( (~ n529)  &  n834  &  n833 ) ;
 assign n511 = ( (~ n63)  &  n513  &  n514 ) | ( n403  &  n513  &  n514 ) ;
 assign n517 = ( (~ i_6_) ) | ( (~ n268) ) | ( (~ n481) ) ;
 assign n518 = ( (~ i_11_) ) | ( n39 ) | ( (~ n185) ) ;
 assign n515 = ( n223  &  n517  &  n518 ) | ( n517  &  n518  &  (~ n529) ) ;
 assign n519 = ( (~ i_4_)  &  n264 ) | ( i_6_  &  n264 ) | ( n196  &  n264 ) ;
 assign n521 = ( (~ i_7_)  &  n522 ) ;
 assign n520 = ( i_2_  &  i_12_  &  n521 ) ;
 assign n522 = ( i_10_  &  (~ i_11_) ) ;
 assign n524 = ( (~ i_4_) ) | ( i_8_ ) | ( n118 ) ;
 assign n523 = ( n32  &  n524 ) | ( (~ n276)  &  n524 ) ;
 assign n525 = ( (~ n36)  &  (~ n664) ) | ( i_3_  &  (~ n36)  &  (~ n228) ) ;
 assign n529 = ( i_4_  &  n268 ) ;
 assign n528 = ( i_6_  &  n520 ) | ( i_6_  &  (~ n46)  &  n529 ) ;
 assign n532 = ( i_4_  &  n651 ) | ( n507  &  n651 ) | ( i_4_  &  n42 ) | ( n507  &  n42 ) ;
 assign n533 = ( i_0_  &  (~ i_7_) ) | ( (~ i_7_)  &  n511 ) | ( i_0_  &  n515 ) | ( n511  &  n515 ) ;
 assign n534 = ( n76  &  (~ n406) ) | ( n322  &  (~ n406) ) | ( n76  &  n519 ) | ( n322  &  n519 ) ;
 assign n535 = ( (~ i_1_)  &  (~ n529) ) | ( (~ n448)  &  (~ n529) ) | ( (~ i_1_)  &  n832 ) | ( (~ n448)  &  n832 ) ;
 assign n537 = ( n173  &  n497 ) | ( n497  &  n523 ) | ( n173  &  (~ n830) ) | ( n523  &  (~ n830) ) ;
 assign n538 = ( n39  &  (~ n525) ) | ( n125  &  (~ n525) ) | ( (~ n525)  &  (~ n604) ) ;
 assign n531 = ( n395  &  (~ n528)  &  n532  &  n533  &  n534  &  n535  &  n537  &  n538 ) ;
 assign n539 = ( (~ i_4_)  &  n198 ) | ( i_10_  &  n198 ) | ( n56  &  n198 ) ;
 assign n541 = ( i_9_ ) | ( i_11_ ) | ( i_7_ ) ;
 assign n540 = ( n207  &  n235 ) | ( n207  &  n541 ) ;
 assign n542 = ( (~ i_8_) ) | ( (~ i_9_) ) ;
 assign n543 = ( i_5_  &  (~ n674)  &  (~ n697) ) | ( i_5_  &  (~ n697)  &  (~ n708) ) ;
 assign n548 = ( i_10_  &  n653 ) ;
 assign n547 = ( (~ i_4_)  &  n548  &  (~ n673) ) | ( (~ i_4_)  &  (~ n673)  &  (~ n708) ) ;
 assign n551 = ( (~ i_8_) ) | ( n236 ) ;
 assign n552 = ( i_8_ ) | ( n650 ) ;
 assign n550 = ( (~ n186)  &  n454 ) | ( (~ n186)  &  n551 ) | ( n454  &  n552 ) | ( n551  &  n552 ) ;
 assign n553 = ( (~ i_12_)  &  (~ n174) ) | ( (~ i_12_)  &  n521 ) | ( (~ i_12_)  &  (~ n664) ) ;
 assign n556 = ( (~ i_3_) ) | ( n113 ) | ( n542 ) ;
 assign n554 = ( i_11_  &  (~ n553)  &  n556 ) | ( n116  &  (~ n553)  &  n556 ) ;
 assign n557 = ( (~ i_0_) ) | ( (~ i_2_) ) ;
 assign n559 = ( i_3_  &  i_5_  &  (~ i_6_) ) ;
 assign n558 = ( n479  &  (~ n848) ) | ( (~ i_7_)  &  n479  &  n559 ) ;
 assign n561 = ( n506  &  (~ n849) ) | ( i_7_  &  n506  &  (~ n682) ) ;
 assign n565 = ( i_5_ ) | ( (~ n453) ) ;
 assign n564 = ( (~ n104)  &  (~ n406) ) | ( (~ n406)  &  (~ n421) ) | ( (~ n104)  &  n565 ) | ( (~ n421)  &  n565 ) ;
 assign n568 = ( i_5_ ) | ( n656 ) ;
 assign n567 = ( n78  &  n77 ) | ( n568  &  n77 ) | ( n78  &  n552 ) | ( n568  &  n552 ) ;
 assign n570 = ( (~ i_5_) ) | ( (~ n653) ) ;
 assign n569 = ( n551  &  n570 ) | ( n77  &  n570 ) | ( n551  &  n78 ) | ( n77  &  n78 ) ;
 assign n572 = ( n149  &  n508 ) ;
 assign n573 = ( (~ i_0_) ) | ( n376 ) ;
 assign n571 = ( n572  &  n471 ) | ( n570  &  n471 ) | ( n572  &  n573 ) | ( n570  &  n573 ) ;
 assign n575 = ( i_0_  &  i_3_  &  (~ i_5_) ) ;
 assign n574 = ( n186  &  (~ n823) ) | ( (~ n108)  &  n186  &  n575 ) ;
 assign n578 = ( (~ i_0_)  &  (~ i_2_)  &  i_4_ ) ;
 assign n577 = ( (~ n709)  &  (~ n824) ) | ( n268  &  n578  &  (~ n709) ) ;
 assign n584 = ( (~ i_5_)  &  n653 ) ;
 assign n582 = ( (~ i_0_)  &  (~ i_1_)  &  i_4_ ) ;
 assign n581 = ( n584  &  (~ n825) ) | ( n268  &  n584  &  n582 ) ;
 assign n585 = ( (~ n710)  &  (~ n826) ) | ( (~ n61)  &  n582  &  (~ n710) ) ;
 assign n588 = ( (~ n711)  &  (~ n827) ) | ( (~ n61)  &  n578  &  (~ n711) ) ;
 assign n591 = ( n506  &  n547 ) | ( n308  &  n506  &  (~ n682) ) ;
 assign n592 = ( n479  &  n543 ) | ( (~ n351)  &  n479  &  n559 ) ;
 assign n596 = ( n550  &  n564 ) | ( n43  &  n564 ) | ( n550  &  n39 ) | ( n43  &  n39 ) ;
 assign n597 = ( (~ i_9_)  &  (~ n581) ) | ( n174  &  (~ n581) ) | ( n497  &  (~ n581) ) ;
 assign n599 = ( n874  &  n872  &  n567 ) | ( n874  &  n872  &  n32 ) ;
 assign n600 = ( n871  &  n869  &  n571 ) | ( n871  &  n869  &  n454 ) ;
 assign n601 = ( n876  &  n878  &  n879  &  n882  &  n884  &  n885  &  (~ n932)  &  (~ n933) ) ;
 assign n602 = ( (~ i_5_) ) | ( n426 ) ;
 assign n604 = ( (~ i_3_)  &  i_8_ ) ;
 assign n603 = ( i_7_  &  (~ n39) ) | ( (~ n39)  &  n604 ) ;
 assign n607 = ( n736  &  i_1_ ) | ( n197  &  i_1_ ) | ( n736  &  n671 ) | ( n197  &  n671 ) ;
 assign n608 = ( n402  &  (~ n603)  &  n896 ) | ( n602  &  (~ n603)  &  n896 ) ;
 assign n606 = ( i_0_  &  n607  &  n608 ) | ( (~ i_5_)  &  n607  &  n608 ) ;
 assign n609 = ( (~ i_7_)  &  (~ n39) ) | ( (~ n39)  &  n276 ) ;
 assign n610 = ( n357  &  i_1_ ) | ( n357  &  n437 ) ;
 assign n612 = ( n942  &  i_5_ ) | ( n942  &  n519 ) ;
 assign n613 = ( n203  &  i_3_ ) | ( n203  &  n348 ) ;
 assign n614 = ( i_12_  &  n39 ) | ( i_12_  &  (~ n453) ) | ( n39  &  n606 ) | ( (~ n453)  &  n606 ) ;
 assign n615 = ( n235  &  n232 ) | ( n714  &  n232 ) | ( n235  &  n353 ) | ( n714  &  n353 ) ;
 assign n616 = ( n898  &  i_1_ ) | ( n898  &  n437 ) | ( n898  &  n668 ) ;
 assign n617 = ( n899  &  i_11_ ) | ( n899  &  n894  &  n891 ) ;
 assign n611 = ( n539  &  n540  &  n612  &  n613  &  n614  &  n615  &  n616  &  n617 ) ;
 assign n620 = ( (~ i_7_) ) | ( n454 ) ;
 assign n619 = ( (~ i_10_) ) | ( (~ i_12_) ) ;
 assign n618 = ( i_7_  &  n620  &  (~ n626) ) | ( n620  &  n619  &  (~ n626) ) ;
 assign n622 = ( (~ i_5_)  &  n943 ) | ( i_5_  &  n944 ) | ( n943  &  n944 ) ;
 assign n621 = ( (~ i_0_)  &  n622 ) | ( n334  &  n622 ) ;
 assign n624 = ( i_8_ ) | ( (~ i_11_) ) ;
 assign n623 = ( (~ i_3_)  &  n312  &  n624  &  (~ n626) ) ;
 assign n626 = ( i_8_  &  i_12_ ) ;
 assign n625 = ( (~ n240)  &  n626 ) | ( (~ n471)  &  n626 ) ;
 assign n628 = ( (~ i_1_)  &  n237 ) | ( (~ i_1_)  &  n618 ) | ( n237  &  n621 ) | ( n618  &  n621 ) ;
 assign n629 = ( (~ i_12_)  &  n909 ) | ( n41  &  n905  &  n909 ) ;
 assign n630 = ( (~ i_11_)  &  n908 ) | ( n900  &  n904  &  n908 ) ;
 assign n631 = ( n906  &  n624 ) | ( n906  &  n250  &  n470 ) ;
 assign n627 = ( n628  &  n629  &  n630  &  n631 ) ;
 assign n633 = ( i_12_ ) | ( (~ n604) ) ;
 assign n632 = ( i_11_  &  (~ n23)  &  n633 ) | ( (~ n23)  &  (~ n276)  &  n633 ) ;
 assign n635 = ( n114  &  (~ n276) ) | ( n114  &  (~ n406) ) | ( (~ n276)  &  (~ n488) ) | ( (~ n406)  &  (~ n488) ) ;
 assign n637 = ( (~ n50)  &  (~ n276) ) | ( (~ n50)  &  (~ n287) ) | ( (~ n276)  &  (~ n604) ) | ( (~ n287)  &  (~ n604) ) ;
 assign n638 = ( (~ i_4_)  &  n632 ) | ( i_4_  &  n635 ) | ( n632  &  n635 ) ;
 assign n639 = ( (~ i_13_)  &  n910  &  n911 ) | ( (~ n23)  &  n910  &  n911 ) ;
 assign n636 = ( n637  &  n638  &  n639 ) ;
 assign n641 = ( (~ i_1_)  &  (~ i_2_) ) | ( (~ i_1_)  &  n312 ) | ( (~ i_2_)  &  n334 ) | ( n312  &  n334 ) ;
 assign n640 = ( i_5_  &  (~ i_9_) ) | ( (~ i_5_)  &  (~ i_10_) ) | ( (~ i_9_)  &  (~ i_10_) ) ;
 assign n647 = ( i_6_  &  (~ i_12_) ) ;
 assign n646 = ( i_9_  &  n487 ) | ( i_9_  &  n647  &  i_1_ ) ;
 assign n648 = ( i_9_ ) | ( i_10_ ) ;
 assign n649 = ( i_3_ ) | ( i_4_ ) ;
 assign n650 = ( i_5_ ) | ( i_6_ ) ;
 assign n651 = ( i_8_ ) | ( (~ n522) ) ;
 assign n652 = ( (~ i_8_) ) | ( n38 ) ;
 assign n653 = ( i_8_  &  i_7_ ) ;
 assign n654 = ( (~ i_8_) ) | ( n364 ) ;
 assign n655 = ( (~ i_0_) ) | ( (~ i_1_) ) | ( i_2_ ) ;
 assign n656 = ( i_8_ ) | ( i_7_ ) ;
 assign n657 = ( i_11_ ) | ( n648 ) ;
 assign n658 = ( (~ i_5_) ) | ( n649 ) ;
 assign n659 = ( (~ n421) ) | ( n657 ) ;
 assign n660 = ( (~ i_9_) ) | ( (~ i_10_) ) ;
 assign n661 = ( i_7_ ) | ( n660 ) ;
 assign n662 = ( (~ i_3_) ) | ( n660 ) ;
 assign n663 = ( (~ i_7_) ) | ( n660 ) ;
 assign n664 = ( i_11_ ) | ( n313 ) ;
 assign n665 = ( (~ i_3_) ) | ( (~ i_4_) ) | ( (~ i_5_) ) ;
 assign n666 = ( (~ i_6_) ) | ( n398 ) ;
 assign n667 = ( (~ i_8_) ) | ( n398 ) ;
 assign n668 = ( i_5_ ) | ( i_10_ ) ;
 assign n669 = ( i_7_ ) | ( n668 ) ;
 assign n670 = ( (~ i_2_)  &  n453 ) ;
 assign n671 = ( i_9_ ) | ( n236 ) ;
 assign n672 = ( (~ i_5_) ) | ( n398 ) ;
 assign n673 = ( i_5_ ) | ( (~ i_6_) ) ;
 assign n674 = ( (~ i_9_) ) | ( n656 ) ;
 assign n675 = ( (~ n287) ) | ( n674 ) ;
 assign n677 = ( (~ n50) ) | ( (~ n308) ) ;
 assign n680 = ( (~ n268) ) | ( n565 ) ;
 assign n681 = ( (~ n287) ) | ( n351 ) ;
 assign n682 = ( (~ i_3_) ) | ( n673 ) ;
 assign n683 = ( (~ i_3_) ) | ( n650 ) ;
 assign n684 = ( (~ i_3_) ) | ( n236 ) ;
 assign n685 = ( (~ i_7_) ) | ( n542 ) ;
 assign n686 = ( (~ n287) ) | ( n685 ) ;
 assign n687 = ( (~ n50) ) | ( n317 ) ;
 assign n688 = ( (~ n287) ) | ( n318 ) ;
 assign n690 = ( i_13_ ) | ( n116 ) ;
 assign n691 = ( (~ i_11_) ) | ( (~ n499) ) ;
 assign n692 = ( i_13_ ) | ( n174 ) ;
 assign n693 = ( (~ i_9_) ) | ( (~ n506) ) ;
 assign n695 = ( n112  &  n662 ) ;
 assign n696 = ( (~ i_2_) ) | ( (~ i_3_) ) ;
 assign n697 = ( i_4_ ) | ( i_6_ ) ;
 assign n698 = ( (~ i_3_) ) | ( i_12_ ) ;
 assign n699 = ( i_4_ ) | ( n247 ) ;
 assign n700 = ( i_1_ ) | ( n696 ) ;
 assign n701 = ( (~ i_1_) ) | ( n45 ) ;
 assign n702 = ( i_7_ ) | ( i_2_ ) ;
 assign n703 = ( (~ i_11_) ) | ( n619 ) ;
 assign n704 = ( (~ i_9_) ) | ( n619 ) ;
 assign n705 = ( (~ i_9_) ) | ( (~ n186) ) ;
 assign n707 = ( (~ i_8_) ) | ( n341 ) ;
 assign n708 = ( i_0_ ) | ( n696 ) ;
 assign n709 = ( (~ i_8_) ) | ( n673 ) ;
 assign n710 = ( (~ i_5_) ) | ( n656 ) ;
 assign n711 = ( (~ i_5_) ) | ( n74 ) ;
 assign n712 = ( (~ n241) ) | ( n344 ) ;
 assign n713 = ( n276  &  n383 ) ;
 assign n714 = ( i_12_ ) | ( n326 ) ;
 assign n716 = ( i_5_  &  n499 ) | ( (~ i_5_)  &  n522 ) | ( n499  &  n522 ) ;
 assign n717 = ( i_4_  &  n82 ) | ( (~ i_4_)  &  n912 ) | ( n82  &  n912 ) ;
 assign n718 = ( i_6_  &  n449 ) | ( (~ i_6_)  &  n703 ) | ( n449  &  n703 ) ;
 assign n719 = ( (~ i_6_)  &  (~ n196) ) | ( i_6_  &  (~ n197) ) | ( (~ n196)  &  (~ n197) ) ;
 assign n722 = ( i_10_ ) | ( i_13_ ) | ( (~ n479) ) | ( n654 ) ;
 assign n720 = ( n256  &  n722 ) | ( (~ n280)  &  n722 ) ;
 assign n725 = ( i_9_ ) | ( i_13_ ) | ( n98 ) | ( (~ n506) ) ;
 assign n723 = ( n95  &  n725 ) | ( (~ n271)  &  n725 ) ;
 assign n727 = ( (~ i_3_) ) | ( n251 ) | ( n661 ) ;
 assign n726 = ( n727  &  i_8_ ) | ( n727  &  n250 ) | ( n727  &  n660 ) ;
 assign n728 = ( n231  &  n232 ) | ( n232  &  (~ n448) ) | ( n231  &  n651 ) | ( (~ n448)  &  n651 ) ;
 assign n730 = ( n228  &  (~ n243)  &  n728 ) | ( n235  &  (~ n243)  &  n728 ) ;
 assign n733 = ( n20  &  n224  &  n508  &  n684 ) ;
 assign n732 = ( i_0_  &  n733 ) | ( n227  &  n733 ) | ( i_0_  &  n663 ) | ( n227  &  n663 ) ;
 assign n736 = ( n223  &  n218  &  n215 ) ;
 assign n734 = ( n221  &  n664 ) | ( (~ n521)  &  n664 ) | ( n221  &  n736 ) | ( (~ n521)  &  n736 ) ;
 assign n738 = ( n429  &  n428 ) ;
 assign n740 = ( n46  &  n324 ) | ( n666  &  n324 ) | ( n46  &  n223 ) | ( n666  &  n223 ) ;
 assign n742 = ( n675 ) | ( n217 ) ;
 assign n743 = ( n168 ) | ( n174 ) | ( n114 ) ;
 assign n744 = ( n108 ) | ( n174 ) | ( (~ n499) ) ;
 assign n745 = ( (~ n559) ) | ( n687 ) ;
 assign n746 = ( (~ n559) ) | ( n686 ) ;
 assign n747 = ( n140 ) | ( n174 ) | ( n114 ) ;
 assign n748 = ( n217  &  (~ n308) ) | ( (~ n308)  &  (~ n653) ) | ( n217  &  n684 ) | ( (~ n653)  &  n684 ) ;
 assign n749 = ( n662  &  n683 ) | ( n662  &  n317 ) ;
 assign n751 = ( (~ n53) ) | ( n114 ) | ( n665 ) ;
 assign n750 = ( n751  &  n115 ) | ( n751  &  n108 ) ;
 assign n752 = ( n220  &  n98 ) | ( n165  &  n98 ) | ( n220  &  n145 ) | ( n165  &  n145 ) ;
 assign n753 = ( n750  &  n752  &  n217 ) | ( n750  &  n752  &  n688 ) ;
 assign n754 = ( n109  &  n105 ) | ( n658  &  n105 ) | ( n109  &  n124 ) | ( n658  &  n124 ) ;
 assign n755 = ( i_4_  &  (~ n119)  &  n754 ) | ( (~ n119)  &  n695  &  n754 ) ;
 assign n757 = ( n36  &  n652 ) | ( n654  &  n652 ) | ( n36  &  n40 ) | ( n654  &  n40 ) ;
 assign n758 = ( n89  &  n92 ) | ( n92  &  (~ n181) ) | ( n89  &  n565 ) | ( (~ n181)  &  n565 ) ;
 assign n759 = ( n97  &  (~ n100)  &  n758 ) | ( (~ n100)  &  n665  &  n758 ) ;
 assign n761 = ( n602  &  n671 ) | ( n259  &  n671 ) | ( n602  &  n260 ) | ( n259  &  n260 ) ;
 assign n762 = ( n672  &  n324 ) | ( n42  &  n324 ) | ( n672  &  n508 ) | ( n42  &  n508 ) ;
 assign n764 = ( (~ i_6_) ) | ( i_11_ ) | ( n44 ) ;
 assign n763 = ( (~ i_10_)  &  n764 ) | ( n41  &  n764 ) ;
 assign n766 = ( i_10_ ) | ( (~ n102) ) | ( (~ n383) ) | ( n654 ) ;
 assign n765 = ( n766  &  n37 ) | ( n766  &  n179 ) ;
 assign n768 = ( i_10_ ) | ( n173 ) | ( (~ n383) ) | ( n652 ) ;
 assign n767 = ( n768  &  n26 ) | ( n768  &  n40 ) | ( n768  &  n125 ) ;
 assign n769 = ( n767  &  n654 ) | ( n767  &  n655 ) | ( n767  &  n32 ) ;
 assign n770 = ( n30  &  n34 ) | ( n30  &  (~ n53) ) | ( n34  &  (~ n101) ) | ( (~ n53)  &  (~ n101) ) ;
 assign n772 = ( (~ n101) ) | ( n125 ) | ( n178 ) | ( n668 ) ;
 assign n771 = ( i_4_  &  n772 ) | ( n42  &  n772 ) | ( (~ n716)  &  n772 ) ;
 assign n773 = ( (~ n51)  &  n116 ) | ( (~ n51)  &  n769  &  n770 ) ;
 assign n775 = ( i_10_  &  i_2_ ) | ( n402  &  i_2_ ) | ( i_10_  &  n428 ) | ( n402  &  n428 ) ;
 assign n777 = ( n42 ) | ( n697 ) | ( i_11_ ) | ( n317 ) ;
 assign n776 = ( n777  &  i_9_ ) | ( n777  &  n258 ) | ( n777  &  n73 ) ;
 assign n779 = ( (~ i_2_) ) | ( n61 ) | ( n429 ) ;
 assign n778 = ( n779  &  n241 ) | ( n779  &  n61 ) | ( n779  &  n197 ) ;
 assign n781 = ( i_10_ ) | ( (~ n296) ) | ( n398 ) ;
 assign n780 = ( (~ n185)  &  n781 ) | ( n253  &  n781 ) | ( n396  &  n781 ) ;
 assign n782 = ( (~ i_13_)  &  n780 ) | ( n470  &  n780 ) | ( n651  &  n780 ) ;
 assign n785 = ( n212 ) | ( (~ n268) ) | ( n665 ) ;
 assign n783 = ( (~ n102)  &  (~ n292)  &  n785 ) | ( n192  &  (~ n292)  &  n785 ) ;
 assign n788 = ( n187  &  n169 ) | ( n173  &  n169 ) | ( n187  &  n655 ) | ( n173  &  n655 ) ;
 assign n789 = ( n788  &  n163 ) | ( n788  &  n36 ) ;
 assign n790 = ( n156  &  n143 ) | ( n40  &  n143 ) | ( n156  &  n31 ) | ( n40  &  n31 ) ;
 assign n791 = ( n790  &  n789  &  n131 ) | ( n790  &  n789  &  n39 ) ;
 assign n792 = ( (~ n297)  &  n497 ) | ( (~ n297)  &  n753  &  n755 ) ;
 assign n794 = ( (~ i_7_)  &  n914 ) | ( n320  &  n914 ) ;
 assign n796 = ( (~ i_4_) ) | ( n73 ) | ( (~ n542) ) ;
 assign n795 = ( n796  &  i_8_ ) | ( n796  &  i_13_ ) | ( n796  &  n260 ) ;
 assign n797 = ( i_11_  &  (~ n406) ) | ( n178  &  (~ n406) ) | ( i_11_  &  (~ n670) ) | ( n178  &  (~ n670) ) ;
 assign n799 = ( (~ i_8_) ) | ( i_13_ ) | ( n260 ) ;
 assign n798 = ( (~ n421)  &  n799 ) | ( n667  &  (~ n670)  &  n799 ) ;
 assign n802 = ( (~ i_2_) ) | ( n312 ) | ( n376 ) ;
 assign n803 = ( i_7_  &  (~ n916) ) | ( n795  &  n797  &  (~ n916) ) ;
 assign n805 = ( (~ n448) ) | ( (~ n626) ) | ( (~ n702) ) ;
 assign n804 = ( n805  &  n437 ) | ( n805  &  n700 ) ;
 assign n806 = ( (~ n185)  &  n344 ) | ( (~ n185)  &  n428 ) | ( n344  &  n429 ) | ( n428  &  n429 ) ;
 assign n808 = ( i_3_ ) | ( i_6_ ) | ( (~ i_8_) ) | ( i_10_ ) | ( (~ n185) ) | ( n945 ) ;
 assign n807 = ( (~ n421)  &  n808 ) | ( n425  &  n808 ) ;
 assign n810 = ( n945 ) | ( n624 ) | ( i_10_ ) | ( i_13_ ) ;
 assign n809 = ( n810  &  n118 ) | ( n810  &  n701 ) ;
 assign n812 = ( i_10_ ) | ( i_8_ ) ;
 assign n813 = ( n205  &  n341 ) | ( n205  &  (~ n409) ) | ( n341  &  n812 ) | ( (~ n409)  &  n812 ) ;
 assign n814 = ( i_8_ ) | ( (~ n383) ) | ( n402 ) ;
 assign n816 = ( (~ i_6_) ) | ( (~ i_12_) ) | ( n453 ) | ( n685 ) ;
 assign n818 = ( (~ i_3_) ) | ( (~ i_9_) ) | ( (~ n479) ) | ( n652 ) ;
 assign n817 = ( n334  &  n818 ) | ( (~ n626)  &  n818 ) | ( n699  &  n818 ) ;
 assign n819 = ( n417  &  n434 ) | ( n365  &  n434 ) | ( n417  &  n99 ) | ( n365  &  n99 ) ;
 assign n821 = ( (~ i_6_)  &  n410 ) | ( i_6_  &  n422 ) | ( n410  &  n422 ) ;
 assign n822 = ( i_1_  &  n369 ) | ( (~ i_1_)  &  n392 ) | ( n369  &  n392 ) ;
 assign n820 = ( (~ i_12_)  &  n821  &  n822 ) | ( n430  &  n821  &  n822 ) ;
 assign n823 = ( n572  &  n470 ) | ( n568  &  n470 ) | ( n572  &  n573 ) | ( n568  &  n573 ) ;
 assign n824 = ( n46  &  n693 ) | ( (~ n280)  &  n693 ) | ( n46  &  n708 ) | ( (~ n280)  &  n708 ) ;
 assign n825 = ( n223  &  n483 ) | ( (~ n280)  &  n483 ) | ( n223  &  n693 ) | ( (~ n280)  &  n693 ) ;
 assign n826 = ( n223  &  n483 ) | ( (~ n271)  &  n483 ) | ( n223  &  n691 ) | ( (~ n271)  &  n691 ) ;
 assign n827 = ( n46  &  n691 ) | ( (~ n271)  &  n691 ) | ( n46  &  n708 ) | ( (~ n271)  &  n708 ) ;
 assign n828 = ( (~ n185)  &  n344 ) | ( n209  &  n344 ) | ( (~ n185)  &  n669 ) | ( n209  &  n669 ) ;
 assign n829 = ( (~ n104)  &  n118 ) | ( n114  &  n118 ) | ( (~ n104)  &  n565 ) | ( n114  &  n565 ) ;
 assign n830 = ( (~ i_7_)  &  i_10_ ) | ( i_3_  &  (~ i_8_)  &  i_10_ ) ;
 assign n832 = ( (~ i_8_) ) | ( n39 ) ;
 assign n834 = ( (~ i_2_)  &  n934 ) | ( n365  &  n934 ) | ( (~ n506)  &  n934 ) ;
 assign n833 = ( (~ i_3_)  &  (~ n280) ) | ( i_3_  &  n693 ) | ( (~ n280)  &  n693 ) ;
 assign n835 = ( i_0_  &  (~ i_7_) ) | ( (~ i_7_)  &  (~ n53) ) | ( i_0_  &  n483 ) | ( (~ n53)  &  n483 ) ;
 assign n838 = ( i_8_ ) | ( n36 ) | ( (~ n479) ) ;
 assign n837 = ( n838  &  n496 ) | ( n838  &  n454 ) ;
 assign n841 = ( (~ i_8_) ) | ( n114 ) | ( n173 ) ;
 assign n840 = ( (~ n421)  &  n841 ) | ( n495  &  n841 ) ;
 assign n844 = ( i_6_ ) | ( n494 ) | ( n417 ) ;
 assign n843 = ( n844  &  n486 ) | ( n844  &  n455 ) ;
 assign n845 = ( n173  &  (~ n276) ) | ( (~ n276)  &  n320 ) | ( n173  &  n659 ) | ( n320  &  n659 ) ;
 assign n846 = ( n39  &  n843  &  n845 ) | ( (~ n713)  &  n843  &  n845 ) ;
 assign n847 = ( i_0_  &  i_7_ ) | ( n491  &  i_7_ ) | ( i_0_  &  n482 ) | ( n491  &  n482 ) ;
 assign n848 = ( (~ i_1_)  &  (~ i_2_) ) | ( (~ i_2_)  &  n710 ) | ( (~ i_1_)  &  n711 ) | ( n710  &  n711 ) ;
 assign n849 = ( (~ i_1_)  &  (~ i_2_) ) | ( (~ i_2_)  &  (~ n584) ) | ( (~ i_1_)  &  n709 ) | ( (~ n584)  &  n709 ) ;
 assign n851 = ( n106  &  n455 ) | ( n671  &  n455 ) | ( n106  &  n551 ) | ( n671  &  n551 ) ;
 assign n852 = ( i_2_ ) | ( n107 ) | ( n344 ) ;
 assign n854 = ( n455  &  n568 ) | ( n570  &  n568 ) | ( n455  &  n323 ) | ( n570  &  n323 ) ;
 assign n857 = ( i_10_ ) | ( n106 ) | ( n234 ) ;
 assign n856 = ( (~ i_9_)  &  n857 ) | ( n670  &  n857 ) | ( n703  &  n857 ) ;
 assign n858 = ( (~ n453)  &  (~ n472)  &  n856 ) | ( n469  &  (~ n472)  &  n856 ) ;
 assign n863 = ( i_13_ ) | ( n348 ) | ( i_3_ ) ;
 assign n862 = ( (~ i_6_)  &  n922 ) | ( (~ i_12_)  &  n922 ) | ( n663  &  n922 ) ;
 assign n861 = ( (~ i_3_)  &  n336  &  n863 ) | ( n336  &  n863  &  n862 ) ;
 assign n867 = ( i_5_  &  n456 ) | ( (~ i_5_)  &  n466 ) | ( n456  &  n466 ) ;
 assign n865 = ( (~ i_1_)  &  n867  &  (~ n930) ) | ( n660  &  n867  &  (~ n930) ) ;
 assign n870 = ( i_8_ ) | ( (~ n575) ) | ( n703 ) ;
 assign n869 = ( n870  &  n232 ) | ( n870  &  n306 ) | ( n870  &  n403 ) ;
 assign n871 = ( (~ i_10_) ) | ( n116 ) | ( n497 ) ;
 assign n873 = ( n219 ) | ( n125 ) | ( n707 ) ;
 assign n872 = ( n873  &  n569 ) | ( n873  &  n110 ) ;
 assign n874 = ( n215 ) | ( n346 ) | ( (~ n383) ) ;
 assign n876 = ( n173  &  (~ n588) ) | ( (~ n588)  &  n828  &  n829 ) ;
 assign n878 = ( n239  &  n554 ) | ( n704  &  n554 ) | ( n239  &  n36 ) | ( n704  &  n36 ) ;
 assign n879 = ( n151  &  (~ n591)  &  (~ n592) ) | ( n550  &  (~ n591)  &  (~ n592) ) ;
 assign n882 = ( (~ n296)  &  (~ n421) ) | ( (~ n421)  &  n539 ) | ( (~ n296)  &  n540 ) | ( n539  &  n540 ) ;
 assign n884 = ( n705  &  n672 ) | ( n249  &  n672 ) | ( n705  &  n61 ) | ( n249  &  n61 ) ;
 assign n886 = ( n647 ) | ( n500 ) | ( n557 ) | ( i_5_ ) ;
 assign n885 = ( i_5_  &  n886  &  (~ n940) ) | ( n531  &  n886  &  (~ n940) ) ;
 assign n890 = ( n221  &  n736 ) | ( n196  &  n736 ) | ( n221  &  n346 ) | ( n196  &  n346 ) ;
 assign n891 = ( n46  &  (~ n609)  &  n890 ) | ( n428  &  (~ n609)  &  n890 ) ;
 assign n893 = ( n231  &  n204 ) | ( n428  &  n204 ) | ( n231  &  n402 ) | ( n428  &  n402 ) ;
 assign n895 = ( (~ i_5_) ) | ( i_9_ ) | ( (~ n241) ) ;
 assign n894 = ( n895  &  n893  &  i_0_ ) | ( n895  &  n893  &  i_5_ ) ;
 assign n896 = ( n44  &  n221 ) | ( n429  &  n221 ) | ( n44  &  n707 ) | ( n429  &  n707 ) ;
 assign n898 = ( i_10_ ) | ( n398 ) ;
 assign n899 = ( i_0_  &  i_2_ ) | ( n610  &  i_2_ ) | ( i_0_  &  n337 ) | ( n610  &  n337 ) ;
 assign n901 = ( i_6_ ) | ( n43 ) ;
 assign n900 = ( i_5_  &  (~ i_12_)  &  n901 ) | ( (~ i_12_)  &  n42  &  n901 ) ;
 assign n903 = ( (~ i_3_) ) | ( i_7_ ) | ( n251 ) ;
 assign n902 = ( n903  &  i_7_ ) | ( n903  &  n508 ) ;
 assign n904 = ( n683  &  n902 ) | ( (~ i_2_)  &  i_7_  &  n902 ) ;
 assign n905 = ( (~ i_2_)  &  (~ i_7_) ) | ( (~ i_7_)  &  n684 ) | ( (~ i_2_)  &  n733 ) | ( n684  &  n733 ) ;
 assign n906 = ( n246  &  (~ n625) ) | ( n494  &  n500  &  (~ n625) ) ;
 assign n908 = ( (~ i_0_) ) | ( n640 ) ;
 assign n909 = ( n623 ) | ( n497 ) ;
 assign n910 = ( (~ i_3_) ) | ( n323 ) | ( (~ n542) ) ;
 assign n911 = ( (~ i_8_) ) | ( (~ n421) ) | ( (~ n453) ) ;
 assign n912 = ( (~ i_5_) ) | ( n42 ) | ( (~ n647) ) | ( n685 ) ;
 assign n914 = ( i_7_ ) | ( n32 ) | ( (~ n276) ) ;
 assign n915 = ( i_7_  &  n713 ) | ( i_7_  &  n50 ) ;
 assign n916 = ( i_7_  &  (~ n798) ) | ( i_7_  &  (~ i_12_)  &  (~ n178) ) ;
 assign n920 = ( i_12_ ) | ( n648 ) ;
 assign n921 = ( i_8_ ) | ( (~ n186) ) | ( n699 ) ;
 assign n922 = ( i_6_ ) | ( (~ i_11_) ) | ( n661 ) ;
 assign n923 = ( (~ i_10_)  &  (~ n712) ) | ( (~ i_10_)  &  n63  &  n185 ) ;
 assign n927 = ( i_2_  &  i_12_  &  (~ n365) ) | ( i_2_  &  i_12_  &  (~ n494) ) ;
 assign n930 = ( (~ i_1_)  &  (~ n854) ) | ( (~ i_1_)  &  n185  &  (~ n671) ) ;
 assign n932 = ( (~ i_0_)  &  (~ i_4_)  &  n558 ) | ( (~ i_0_)  &  (~ i_4_)  &  n561 ) ;
 assign n933 = ( i_0_  &  (~ n858) ) | ( i_0_  &  (~ n861) ) | ( i_0_  &  (~ n865) ) ;
 assign n934 = ( n99 ) | ( n125 ) | ( i_2_ ) ;
 assign n935 = ( i_4_  &  (~ n840) ) | ( i_4_  &  (~ n56)  &  (~ n61) ) ;
 assign n937 = ( (~ i_4_)  &  (~ n837) ) | ( (~ i_4_)  &  (~ n508)  &  (~ n620) ) ;
 assign n941 = ( n498 ) | ( n646 ) | ( (~ n846) ) | ( (~ n847) ) | ( n935 ) | ( n937 ) ;
 assign n940 = ( i_5_  &  n941 ) ;
 assign n942 = ( (~ i_4_) ) | ( (~ i_5_) ) | ( n495 ) ;
 assign n943 = ( (~ i_6_)  &  (~ n186) ) | ( i_6_  &  n451 ) | ( (~ n186)  &  n451 ) ;
 assign n944 = ( i_6_  &  n454 ) | ( (~ i_6_)  &  n619 ) | ( n454  &  n619 ) ;
 assign n945 = ( i_2_  &  i_7_ ) ;
 assign n946 = ( n667  &  i_3_  &  n521 ) ;
 assign n951 = ( n714  &  n541  &  i_6_ ) ;


endmodule

