module frg2 (
	a, b, c, d, e, f, g, h, 
	i, j, k, l, m, n, o, p, q, r, 
	s, t, u, v, w, x, y, z, a0, b0, 
	c0, d0, e0, f0, g0, h0, i0, j0, k0, l0, 
	m0, n0, o0, p0, q0, s0, t0, u0, v0, w0, 
	x0, y0, z0, a1, b1, c1, d1, e1, f1, g1, 
	h1, i1, j1, k1, l1, m1, n1, o1, p1, q1, 
	r1, s1, t1, u1, v1, w1, x1, y1, z1, a2, 
	b2, c2, d2, e2, f2, g2, h2, i2, j2, k2, 
	l2, m2, n2, o2, p2, q2, r2, s2, t2, u2, 
	v2, w2, x2, y2, z2, a3, b3, c3, d3, e3, 
	f3, g3, h3, i3, j3, k3, l3, m3, n3, o3, 
	p3, q3, r3, s3, t3, u3, v3, w3, x3, y3, 
	z3, a4, b4, c4, d4, e4, f4, g4, h4, i4, 
	j4, k4, l4, m4, n4, o4, p4, q4, r4, s4, 
	t4, u4, v4, w4, x4, y4, z4, a5, b5, c5, 
	d5, e5, f5, g5, h5, i5, j5, k5, l5, m5, 
	n5, o5, p5, q5, r5, s5, t5, u5, v5, w5, 
	x5, y5, z5, a6, b6, c6, d6, e6, f6, g6, 
	h6, i6, j6, k6, l6, m6, n6, o6, p6, q6, 
	r6, s6, t6, u6, v6, w6, x6, y6, z6, a7, 
	b7, c7, d7, e7, f7, g7, h7, i7, j7, k7, 
	l7, m7, n7, o7, p7, q7, r7, s7, t7, u7, 
	v7, w7, x7, y7, z7, a8, b8, c8, d8, e8, 
	f8, g8, h8, i8, j8, k8, l8, m8, n8, o8, 
	p8, q8, r8, s8, t8, u8, v8, w8, x8, y8, 
	z8, a9, b9, c9, d9, e9, f9, g9, h9, i9, 
	j9, k9, l9, m9, n9, o9, p9, q9, r9, s9, 
	t9, u9, v9, w9);

input a, b, c, d, e, f, g, h, i, j, k, l, m, n, o, p, q, r, s, t, u, v, w, x, y, z, a0, b0, c0, d0, e0, f0, g0, h0, i0, j0, k0, l0, m0, n0, o0, p0, q0, s0, t0, u0, v0, w0, x0, y0, z0, a1, b1, c1, d1, e1, f1, g1, h1, i1, j1, k1, l1, m1, n1, o1, p1, q1, r1, s1, t1, u1, v1, w1, x1, y1, z1, a2, b2, c2, d2, e2, f2, g2, h2, i2, j2, k2, l2, m2, n2, o2, p2, q2, r2, s2, t2, u2, v2, w2, x2, y2, z2, a3, b3, c3, d3, e3, f3, g3, h3, i3, j3, k3, l3, m3, n3, o3, p3, q3, r3, s3, t3, u3, v3, w3, x3, y3, z3, a4, b4, c4, d4, e4, f4, g4, h4, i4, j4, k4, l4, m4, n4;

output o4, p4, q4, r4, s4, t4, u4, v4, w4, x4, y4, z4, a5, b5, c5, d5, e5, f5, g5, h5, i5, j5, k5, l5, m5, n5, o5, p5, q5, r5, s5, t5, u5, v5, w5, x5, y5, z5, a6, b6, c6, d6, e6, f6, g6, h6, i6, j6, k6, l6, m6, n6, o6, p6, q6, r6, s6, t6, u6, v6, w6, x6, y6, z6, a7, b7, c7, d7, e7, f7, g7, h7, i7, j7, k7, l7, m7, n7, o7, p7, q7, r7, s7, t7, u7, v7, w7, x7, y7, z7, a8, b8, c8, d8, e8, f8, g8, h8, i8, j8, k8, l8, m8, n8, o8, p8, q8, r8, s8, t8, u8, v8, w8, x8, y8, z8, a9, b9, c9, d9, e9, f9, g9, h9, i9, j9, k9, l9, m9, n9, o9, p9, q9, r9, s9, t9, u9, v9, w9;

wire g15, j15, k15, l15, m15, o15, t15, w15, x15, y15, z15, b16, c16, d16, f16, g16, h16, j16, l16, m16, p16, r16, s16, u16, v16, w16, x16, a17, b17, d17, e17, g17, i17, j17, l17, n17, o17, q17, s17, t17, v17, x17, y17, a18, c18, d18, f18, h18, i18, k18, m18, n18, p18, r18, s18, u18, w18, x18, z18, b19, c19, e19, g19, h19, j19, l19, m19, o19, q19, r19, t19, v19, w19, y19, a20, b20, d20, f20, g20, i20, k20, l20, n20, p20, q20, s20, u20, v20, x20, z20, a21, c21, e21, f21, h21, i21, j21, k21, l21, q21, r21, s21, t21, x21, y21, z21, a22, e22, f22, g22, h22, l22, m22, n22, o22, s22, t22, u22, v22, z22, a23, b23, c23, g23, h23, i23, j23, n23, o23, p23, q23, r23, s23, t23, u23, w23, y23, z23, a24, c24, d24, e24, g24, h24, i24, k24, l24, m24, o24, p24, q24, s24, t24, u24, w24, x24, y24, z24, a25, b25, c25, d25, e25, f25, g25, h25, i25, j25, k25, l25, m25, n25, o25, p25, q25, r25, s25, t25, w25, x25, z25, a26, c26, d26, f26, g26, i26, j26, l26, m26, o26, p26, r26, s26, u26, v26, x26, y26, a27, b27, d27, e27, g27, h27, j27, k27, m27, n27, p27, q27, s27, t27, v27, w27, y27, z27, b28, c28, e28, f28, h28, i28, j28, k28, l28, m28, n28, p28, q28, r28, s28, u28, v28, w28, x28, a29, b29, d29, e29, f29, g29, i29, j29, k29, l29, m29, n29, o29, p29, q29, r29, t29, u29, v29, w29, x29, y29, z29, a30, b30, c30, d30, e30, f30, g30, h30, j30, k30, l30, m30, n30, o30, p30, q30, r30, t30, u30, v30, w30, x30, b31, c31, d31, e31, f31, h31, i31, j31, k31, l31, m31, n31, o31, p31, q31, r31, s31, t31, u31, v31, w31, y31, z31, a32, b32, c32, d32, e32, f32, i32, j32, k32, l32, m32, n32, o32, p32, q32, r32, s32, t32, u32, w32, x32, y32, a33, b33, c33, d33, e33, h33, i33, j33, k33, l33, m33, n33, o33, p33, q33, r33, s33, t33, u33, v33, w33, x33, y33, z33, a34, b34, c34, d34, e34, f34, g34, h34, i34, k34, l34, m34, n34, o34, p34, q34, r34, s34, t34, v34, w34, x34, b35, d35, e35, f35, g35, h35, i35, j35, k35, l35, m35, n35, o35, p35, q35, r35;

assign o4 = ( (~ g1) ) ;
 assign p4 = ( (~ m0)  &  (~ j33) ) | ( (~ k0)  &  (~ h33)  &  (~ j33) ) | ( k0  &  (~ i33)  &  (~ j33) ) | ( (~ h33)  &  (~ i33)  &  (~ j33) ) ;
 assign q4 = ( (~ m0)  &  (~ m33) ) | ( (~ k0)  &  (~ k33)  &  (~ m33) ) | ( k0  &  (~ l33)  &  (~ m33) ) | ( (~ k33)  &  (~ l33)  &  (~ m33) ) ;
 assign r4 = ( (~ m0)  &  (~ p33) ) | ( (~ k0)  &  (~ n33)  &  (~ p33) ) | ( k0  &  (~ o33)  &  (~ p33) ) | ( (~ n33)  &  (~ o33)  &  (~ p33) ) ;
 assign s4 = ( (~ m0)  &  (~ s33) ) | ( (~ k0)  &  (~ q33)  &  (~ s33) ) | ( k0  &  (~ r33)  &  (~ s33) ) | ( (~ q33)  &  (~ r33)  &  (~ s33) ) ;
 assign v4 = ( m3  &  (~ t33) ) | ( k0  &  l0  &  (~ t33) ) | ( (~ k0)  &  (~ l0)  &  (~ t33) ) ;
 assign w4 = ( n3  &  (~ u33) ) | ( k0  &  l0  &  (~ u33) ) | ( (~ k0)  &  (~ l0)  &  (~ u33) ) ;
 assign x4 = ( o3  &  (~ v33) ) | ( k0  &  l0  &  (~ v33) ) | ( (~ k0)  &  (~ l0)  &  (~ v33) ) ;
 assign y4 = ( p3  &  (~ w33) ) | ( k0  &  l0  &  (~ w33) ) | ( (~ k0)  &  (~ l0)  &  (~ w33) ) ;
 assign z4 = ( q3  &  (~ x33) ) | ( k0  &  l0  &  (~ x33) ) | ( (~ k0)  &  (~ l0)  &  (~ x33) ) ;
 assign a5 = ( r3  &  (~ y33) ) | ( k0  &  l0  &  (~ y33) ) | ( (~ k0)  &  (~ l0)  &  (~ y33) ) ;
 assign b5 = ( s3  &  (~ z33) ) | ( k0  &  l0  &  (~ z33) ) | ( (~ k0)  &  (~ l0)  &  (~ z33) ) ;
 assign c5 = ( t3  &  (~ a34) ) | ( k0  &  l0  &  (~ a34) ) | ( (~ k0)  &  (~ l0)  &  (~ a34) ) ;
 assign d5 = ( m3  &  m0 ) ;
 assign e5 = ( n3  &  m0 ) ;
 assign f5 = ( o3  &  m0 ) ;
 assign g5 = ( p3  &  m0 ) ;
 assign h5 = ( q3  &  m0 ) ;
 assign i5 = ( r3  &  m0 ) ;
 assign j5 = ( s3  &  m0 ) ;
 assign k5 = ( t3  &  m0 ) ;
 assign l5 = ( (~ j4)  &  g1 ) ;
 assign n5 = ( (~ b34) ) ;
 assign o5 = ( (~ c34) ) ;
 assign p5 = ( (~ d34) ) ;
 assign q5 = ( (~ e34) ) ;
 assign r5 = ( (~ f34) ) ;
 assign s5 = ( (~ g30)  &  n1 ) | ( (~ g34)  &  n1 ) | ( (~ h34)  &  n1 ) | ( (~ g30)  &  (~ i34) ) | ( (~ g34)  &  (~ i34) ) | ( (~ h34)  &  (~ i34) ) ;
 assign t5 = ( (~ g30)  &  n1 ) | ( (~ g34)  &  n1 ) | ( (~ h34)  &  n1 ) | ( (~ g30)  &  (~ i34) ) | ( (~ g34)  &  (~ i34) ) | ( (~ h34)  &  (~ i34) ) ;
 assign u5 = ( (~ g30)  &  n1 ) | ( (~ g34)  &  n1 ) | ( (~ h34)  &  n1 ) | ( (~ g30)  &  (~ i34) ) | ( (~ g34)  &  (~ i34) ) | ( (~ h34)  &  (~ i34) ) ;
 assign v5 = ( (~ g30)  &  n1 ) | ( (~ g34)  &  n1 ) | ( (~ h34)  &  n1 ) | ( (~ g30)  &  (~ i34) ) | ( (~ g34)  &  (~ i34) ) | ( (~ h34)  &  (~ i34) ) ;
 assign w5 = ( (~ g30)  &  n1 ) | ( (~ g34)  &  n1 ) | ( (~ h34)  &  n1 ) | ( (~ g30)  &  (~ i34) ) | ( (~ g34)  &  (~ i34) ) | ( (~ h34)  &  (~ i34) ) ;
 assign x5 = ( (~ k34) ) ;
 assign y5 = ( (~ l34) ) ;
 assign z5 = ( (~ m34) ) ;
 assign a6 = ( (~ n34) ) ;
 assign b6 = ( (~ o34) ) ;
 assign c6 = ( (~ p34) ) ;
 assign d6 = ( (~ q34) ) ;
 assign e6 = ( (~ r34) ) ;
 assign f6 = ( (~ s34) ) ;
 assign g6 = ( (~ t34) ) ;
 assign h6 = ( (~ h1) ) ;
 assign i6 = ( (~ i1) ) ;
 assign j6 = ( (~ j1) ) ;
 assign k6 = ( (~ k1) ) ;
 assign l6 = ( (~ l1) ) ;
 assign n6 = ( f1  &  i4 ) | ( (~ f1)  &  (~ i4) ) ;
 assign o6 = ( (~ c4)  &  (~ b4)  &  (~ v34) ) ;
 assign p6 = ( (~ g15)  &  (~ q0)  &  o0 ) ;
 assign q6 = ( (~ n0)  &  (~ j15)  &  (~ k15) ) | ( o0  &  (~ l15)  &  (~ m15) ) ;
 assign r6 = ( (~ t15)  &  (~ g1)  &  (~ y15) ) | ( n0  &  (~ g1)  &  (~ y15) ) | ( (~ w15)  &  (~ g1)  &  (~ y15) ) | ( (~ t15)  &  (~ x15)  &  (~ y15) ) | ( n0  &  (~ x15)  &  (~ y15) ) | ( (~ w15)  &  (~ x15)  &  (~ y15) ) ;
 assign s6 = ( (~ t15)  &  (~ g1)  &  (~ c16) ) | ( n0  &  (~ g1)  &  (~ c16) ) | ( (~ b16)  &  (~ g1)  &  (~ c16) ) | ( (~ t15)  &  (~ x15)  &  (~ c16) ) | ( n0  &  (~ x15)  &  (~ c16) ) | ( (~ b16)  &  (~ x15)  &  (~ c16) ) ;
 assign t6 = ( (~ t15)  &  (~ g1)  &  (~ g16) ) | ( n0  &  (~ g1)  &  (~ g16) ) | ( (~ f16)  &  (~ g1)  &  (~ g16) ) | ( (~ t15)  &  (~ x15)  &  (~ g16) ) | ( n0  &  (~ x15)  &  (~ g16) ) | ( (~ f16)  &  (~ x15)  &  (~ g16) ) ;
 assign u6 = ( (~ j16)  &  (~ l16) ) | ( (~ g1)  &  l1  &  (~ l16) ) ;
 assign v6 = ( m1  &  (~ p16) ) | ( (~ n0)  &  p0  &  (~ p16) ) ;
 assign w6 = ( a17  &  n1  &  (~ v16) ) | ( (~ r16)  &  n1  &  (~ v16) ) | ( (~ s16)  &  n1  &  (~ v16) ) | ( a17  &  (~ n0)  &  (~ v16) ) | ( (~ r16)  &  (~ n0)  &  (~ v16) ) | ( (~ s16)  &  (~ n0)  &  (~ v16) ) | ( a17  &  (~ u16)  &  (~ v16) ) | ( (~ r16)  &  (~ u16)  &  (~ v16) ) | ( (~ s16)  &  (~ u16)  &  (~ v16) ) ;
 assign x6 = ( a17  &  o1  &  (~ d17) ) | ( (~ b17)  &  o1  &  (~ d17) ) | ( (~ s16)  &  o1  &  (~ d17) ) | ( a17  &  (~ n0)  &  (~ d17) ) | ( (~ b17)  &  (~ n0)  &  (~ d17) ) | ( (~ s16)  &  (~ n0)  &  (~ d17) ) | ( a17  &  (~ u16)  &  (~ d17) ) | ( (~ b17)  &  (~ u16)  &  (~ d17) ) | ( (~ s16)  &  (~ u16)  &  (~ d17) ) ;
 assign y6 = ( a17  &  p1  &  (~ i17) ) | ( (~ g17)  &  p1  &  (~ i17) ) | ( (~ s16)  &  p1  &  (~ i17) ) | ( a17  &  (~ n0)  &  (~ i17) ) | ( (~ g17)  &  (~ n0)  &  (~ i17) ) | ( (~ s16)  &  (~ n0)  &  (~ i17) ) | ( a17  &  (~ u16)  &  (~ i17) ) | ( (~ g17)  &  (~ u16)  &  (~ i17) ) | ( (~ s16)  &  (~ u16)  &  (~ i17) ) ;
 assign z6 = ( a17  &  q1  &  (~ n17) ) | ( (~ l17)  &  q1  &  (~ n17) ) | ( (~ s16)  &  q1  &  (~ n17) ) | ( a17  &  (~ n0)  &  (~ n17) ) | ( (~ l17)  &  (~ n0)  &  (~ n17) ) | ( (~ s16)  &  (~ n0)  &  (~ n17) ) | ( a17  &  (~ u16)  &  (~ n17) ) | ( (~ l17)  &  (~ u16)  &  (~ n17) ) | ( (~ s16)  &  (~ u16)  &  (~ n17) ) ;
 assign a7 = ( a17  &  r1  &  (~ s17) ) | ( (~ q17)  &  r1  &  (~ s17) ) | ( (~ s16)  &  r1  &  (~ s17) ) | ( a17  &  (~ n0)  &  (~ s17) ) | ( (~ q17)  &  (~ n0)  &  (~ s17) ) | ( (~ s16)  &  (~ n0)  &  (~ s17) ) | ( a17  &  (~ u16)  &  (~ s17) ) | ( (~ q17)  &  (~ u16)  &  (~ s17) ) | ( (~ s16)  &  (~ u16)  &  (~ s17) ) ;
 assign b7 = ( a17  &  s1  &  (~ x17) ) | ( (~ v17)  &  s1  &  (~ x17) ) | ( (~ s16)  &  s1  &  (~ x17) ) | ( a17  &  (~ n0)  &  (~ x17) ) | ( (~ v17)  &  (~ n0)  &  (~ x17) ) | ( (~ s16)  &  (~ n0)  &  (~ x17) ) | ( a17  &  (~ u16)  &  (~ x17) ) | ( (~ v17)  &  (~ u16)  &  (~ x17) ) | ( (~ s16)  &  (~ u16)  &  (~ x17) ) ;
 assign c7 = ( a17  &  t1  &  (~ c18) ) | ( (~ a18)  &  t1  &  (~ c18) ) | ( (~ s16)  &  t1  &  (~ c18) ) | ( a17  &  (~ n0)  &  (~ c18) ) | ( (~ a18)  &  (~ n0)  &  (~ c18) ) | ( (~ s16)  &  (~ n0)  &  (~ c18) ) | ( a17  &  (~ u16)  &  (~ c18) ) | ( (~ a18)  &  (~ u16)  &  (~ c18) ) | ( (~ s16)  &  (~ u16)  &  (~ c18) ) ;
 assign d7 = ( a17  &  u1  &  (~ h18) ) | ( (~ f18)  &  u1  &  (~ h18) ) | ( (~ s16)  &  u1  &  (~ h18) ) | ( a17  &  (~ n0)  &  (~ h18) ) | ( (~ f18)  &  (~ n0)  &  (~ h18) ) | ( (~ s16)  &  (~ n0)  &  (~ h18) ) | ( a17  &  (~ u16)  &  (~ h18) ) | ( (~ f18)  &  (~ u16)  &  (~ h18) ) | ( (~ s16)  &  (~ u16)  &  (~ h18) ) ;
 assign e7 = ( a17  &  v1  &  (~ m18) ) | ( (~ k18)  &  v1  &  (~ m18) ) | ( (~ s16)  &  v1  &  (~ m18) ) | ( a17  &  (~ n0)  &  (~ m18) ) | ( (~ k18)  &  (~ n0)  &  (~ m18) ) | ( (~ s16)  &  (~ n0)  &  (~ m18) ) | ( a17  &  (~ u16)  &  (~ m18) ) | ( (~ k18)  &  (~ u16)  &  (~ m18) ) | ( (~ s16)  &  (~ u16)  &  (~ m18) ) ;
 assign f7 = ( a17  &  w1  &  (~ r18) ) | ( (~ p18)  &  w1  &  (~ r18) ) | ( (~ s16)  &  w1  &  (~ r18) ) | ( a17  &  (~ n0)  &  (~ r18) ) | ( (~ p18)  &  (~ n0)  &  (~ r18) ) | ( (~ s16)  &  (~ n0)  &  (~ r18) ) | ( a17  &  (~ u16)  &  (~ r18) ) | ( (~ p18)  &  (~ u16)  &  (~ r18) ) | ( (~ s16)  &  (~ u16)  &  (~ r18) ) ;
 assign g7 = ( a17  &  x1  &  (~ w18) ) | ( (~ u18)  &  x1  &  (~ w18) ) | ( (~ s16)  &  x1  &  (~ w18) ) | ( a17  &  (~ n0)  &  (~ w18) ) | ( (~ u18)  &  (~ n0)  &  (~ w18) ) | ( (~ s16)  &  (~ n0)  &  (~ w18) ) | ( a17  &  (~ u16)  &  (~ w18) ) | ( (~ u18)  &  (~ u16)  &  (~ w18) ) | ( (~ s16)  &  (~ u16)  &  (~ w18) ) ;
 assign h7 = ( a17  &  y1  &  (~ b19) ) | ( (~ z18)  &  y1  &  (~ b19) ) | ( (~ s16)  &  y1  &  (~ b19) ) | ( a17  &  (~ n0)  &  (~ b19) ) | ( (~ z18)  &  (~ n0)  &  (~ b19) ) | ( (~ s16)  &  (~ n0)  &  (~ b19) ) | ( a17  &  (~ u16)  &  (~ b19) ) | ( (~ z18)  &  (~ u16)  &  (~ b19) ) | ( (~ s16)  &  (~ u16)  &  (~ b19) ) ;
 assign i7 = ( a17  &  z1  &  (~ g19) ) | ( (~ e19)  &  z1  &  (~ g19) ) | ( (~ s16)  &  z1  &  (~ g19) ) | ( a17  &  (~ n0)  &  (~ g19) ) | ( (~ e19)  &  (~ n0)  &  (~ g19) ) | ( (~ s16)  &  (~ n0)  &  (~ g19) ) | ( a17  &  (~ u16)  &  (~ g19) ) | ( (~ e19)  &  (~ u16)  &  (~ g19) ) | ( (~ s16)  &  (~ u16)  &  (~ g19) ) ;
 assign j7 = ( a17  &  a2  &  (~ l19) ) | ( (~ j19)  &  a2  &  (~ l19) ) | ( (~ s16)  &  a2  &  (~ l19) ) | ( a17  &  (~ n0)  &  (~ l19) ) | ( (~ j19)  &  (~ n0)  &  (~ l19) ) | ( (~ s16)  &  (~ n0)  &  (~ l19) ) | ( a17  &  (~ u16)  &  (~ l19) ) | ( (~ j19)  &  (~ u16)  &  (~ l19) ) | ( (~ s16)  &  (~ u16)  &  (~ l19) ) ;
 assign k7 = ( a17  &  b2  &  (~ q19) ) | ( (~ o19)  &  b2  &  (~ q19) ) | ( (~ s16)  &  b2  &  (~ q19) ) | ( a17  &  (~ n0)  &  (~ q19) ) | ( (~ o19)  &  (~ n0)  &  (~ q19) ) | ( (~ s16)  &  (~ n0)  &  (~ q19) ) | ( a17  &  (~ u16)  &  (~ q19) ) | ( (~ o19)  &  (~ u16)  &  (~ q19) ) | ( (~ s16)  &  (~ u16)  &  (~ q19) ) ;
 assign l7 = ( a17  &  c2  &  (~ v19) ) | ( (~ t19)  &  c2  &  (~ v19) ) | ( (~ s16)  &  c2  &  (~ v19) ) | ( a17  &  (~ n0)  &  (~ v19) ) | ( (~ t19)  &  (~ n0)  &  (~ v19) ) | ( (~ s16)  &  (~ n0)  &  (~ v19) ) | ( a17  &  (~ u16)  &  (~ v19) ) | ( (~ t19)  &  (~ u16)  &  (~ v19) ) | ( (~ s16)  &  (~ u16)  &  (~ v19) ) ;
 assign m7 = ( a17  &  d2  &  (~ a20) ) | ( (~ y19)  &  d2  &  (~ a20) ) | ( (~ s16)  &  d2  &  (~ a20) ) | ( a17  &  (~ n0)  &  (~ a20) ) | ( (~ y19)  &  (~ n0)  &  (~ a20) ) | ( (~ s16)  &  (~ n0)  &  (~ a20) ) | ( a17  &  (~ u16)  &  (~ a20) ) | ( (~ y19)  &  (~ u16)  &  (~ a20) ) | ( (~ s16)  &  (~ u16)  &  (~ a20) ) ;
 assign n7 = ( a17  &  e2  &  (~ f20) ) | ( (~ d20)  &  e2  &  (~ f20) ) | ( (~ s16)  &  e2  &  (~ f20) ) | ( a17  &  (~ n0)  &  (~ f20) ) | ( (~ d20)  &  (~ n0)  &  (~ f20) ) | ( (~ s16)  &  (~ n0)  &  (~ f20) ) | ( a17  &  (~ u16)  &  (~ f20) ) | ( (~ d20)  &  (~ u16)  &  (~ f20) ) | ( (~ s16)  &  (~ u16)  &  (~ f20) ) ;
 assign o7 = ( a17  &  f2  &  (~ k20) ) | ( (~ i20)  &  f2  &  (~ k20) ) | ( (~ s16)  &  f2  &  (~ k20) ) | ( a17  &  (~ n0)  &  (~ k20) ) | ( (~ i20)  &  (~ n0)  &  (~ k20) ) | ( (~ s16)  &  (~ n0)  &  (~ k20) ) | ( a17  &  (~ u16)  &  (~ k20) ) | ( (~ i20)  &  (~ u16)  &  (~ k20) ) | ( (~ s16)  &  (~ u16)  &  (~ k20) ) ;
 assign p7 = ( a17  &  g2  &  (~ p20) ) | ( (~ n20)  &  g2  &  (~ p20) ) | ( (~ s16)  &  g2  &  (~ p20) ) | ( a17  &  (~ n0)  &  (~ p20) ) | ( (~ n20)  &  (~ n0)  &  (~ p20) ) | ( (~ s16)  &  (~ n0)  &  (~ p20) ) | ( a17  &  (~ u16)  &  (~ p20) ) | ( (~ n20)  &  (~ u16)  &  (~ p20) ) | ( (~ s16)  &  (~ u16)  &  (~ p20) ) ;
 assign q7 = ( a17  &  h2  &  (~ u20) ) | ( (~ s20)  &  h2  &  (~ u20) ) | ( (~ s16)  &  h2  &  (~ u20) ) | ( a17  &  (~ n0)  &  (~ u20) ) | ( (~ s20)  &  (~ n0)  &  (~ u20) ) | ( (~ s16)  &  (~ n0)  &  (~ u20) ) | ( a17  &  (~ u16)  &  (~ u20) ) | ( (~ s20)  &  (~ u16)  &  (~ u20) ) | ( (~ s16)  &  (~ u16)  &  (~ u20) ) ;
 assign r7 = ( a17  &  i2  &  (~ z20) ) | ( (~ x20)  &  i2  &  (~ z20) ) | ( (~ s16)  &  i2  &  (~ z20) ) | ( a17  &  (~ n0)  &  (~ z20) ) | ( (~ x20)  &  (~ n0)  &  (~ z20) ) | ( (~ s16)  &  (~ n0)  &  (~ z20) ) | ( a17  &  (~ u16)  &  (~ z20) ) | ( (~ x20)  &  (~ u16)  &  (~ z20) ) | ( (~ s16)  &  (~ u16)  &  (~ z20) ) ;
 assign s7 = ( a17  &  j2  &  (~ e21) ) | ( (~ c21)  &  j2  &  (~ e21) ) | ( (~ s16)  &  j2  &  (~ e21) ) | ( a17  &  (~ n0)  &  (~ e21) ) | ( (~ c21)  &  (~ n0)  &  (~ e21) ) | ( (~ s16)  &  (~ n0)  &  (~ e21) ) | ( a17  &  (~ u16)  &  (~ e21) ) | ( (~ c21)  &  (~ u16)  &  (~ e21) ) | ( (~ s16)  &  (~ u16)  &  (~ e21) ) ;
 assign t7 = ( (~ q0)  &  o0  &  (~ h21) ) ;
 assign u7 = ( (~ q0)  &  o0  &  (~ q21) ) ;
 assign v7 = ( (~ q0)  &  o0  &  (~ x21) ) ;
 assign w7 = ( (~ q0)  &  o0  &  (~ e22) ) ;
 assign x7 = ( (~ q0)  &  o0  &  (~ l22) ) ;
 assign y7 = ( (~ q0)  &  o0  &  (~ s22) ) ;
 assign z7 = ( (~ q0)  &  o0  &  (~ z22) ) ;
 assign a8 = ( (~ q0)  &  o0  &  (~ g23) ) ;
 assign b8 = ( (~ q0)  &  o0  &  (~ n23) ) ;
 assign c8 = ( (~ q0)  &  o0  &  (~ y23) ) ;
 assign d8 = ( (~ q0)  &  o0  &  (~ c24) ) ;
 assign e8 = ( (~ q0)  &  o0  &  (~ g24) ) ;
 assign f8 = ( (~ q0)  &  o0  &  (~ k24) ) ;
 assign g8 = ( (~ q0)  &  o0  &  (~ o24) ) ;
 assign h8 = ( (~ q0)  &  o0  &  (~ s24) ) ;
 assign i8 = ( (~ w24)  &  (~ x24)  &  (~ s23) ) | ( o0  &  (~ y24)  &  (~ z24) ) ;
 assign j8 = ( (~ a25)  &  (~ b25)  &  (~ c25) ) | ( o0  &  (~ d25)  &  (~ e25) ) ;
 assign k8 = ( (~ a25)  &  (~ w25)  &  (~ c25) ) | ( o0  &  (~ x25)  &  (~ e25) ) ;
 assign l8 = ( (~ a25)  &  (~ z25)  &  (~ c25) ) | ( o0  &  (~ a26)  &  (~ e25) ) ;
 assign m8 = ( (~ a25)  &  (~ c26)  &  (~ c25) ) | ( o0  &  (~ d26)  &  (~ e25) ) ;
 assign n8 = ( (~ a25)  &  (~ f26)  &  (~ c25) ) | ( o0  &  (~ g26)  &  (~ e25) ) ;
 assign o8 = ( (~ a25)  &  (~ i26)  &  (~ c25) ) | ( o0  &  (~ j26)  &  (~ e25) ) ;
 assign p8 = ( (~ a25)  &  (~ l26)  &  (~ c25) ) | ( o0  &  (~ m26)  &  (~ e25) ) ;
 assign q8 = ( (~ a25)  &  (~ o26)  &  (~ c25) ) | ( o0  &  (~ p26)  &  (~ e25) ) ;
 assign r8 = ( (~ a25)  &  (~ r26)  &  (~ c25) ) | ( o0  &  (~ s26)  &  (~ e25) ) ;
 assign s8 = ( (~ a25)  &  (~ u26)  &  (~ c25) ) | ( o0  &  (~ v26)  &  (~ e25) ) ;
 assign t8 = ( (~ a25)  &  (~ x26)  &  (~ c25) ) | ( o0  &  (~ y26)  &  (~ e25) ) ;
 assign u8 = ( (~ a25)  &  (~ a27)  &  (~ c25) ) | ( o0  &  (~ b27)  &  (~ e25) ) ;
 assign v8 = ( (~ a25)  &  (~ d27)  &  (~ c25) ) | ( o0  &  (~ e27)  &  (~ e25) ) ;
 assign w8 = ( (~ a25)  &  (~ g27)  &  (~ c25) ) | ( o0  &  (~ h27)  &  (~ e25) ) ;
 assign x8 = ( (~ a25)  &  (~ j27)  &  (~ c25) ) | ( o0  &  (~ k27)  &  (~ e25) ) ;
 assign y8 = ( (~ a25)  &  (~ m27)  &  (~ c25) ) | ( o0  &  (~ n27)  &  (~ e25) ) ;
 assign z8 = ( (~ a25)  &  (~ p27)  &  (~ c25) ) | ( o0  &  (~ q27)  &  (~ e25) ) ;
 assign a9 = ( (~ a25)  &  (~ s27)  &  (~ c25) ) | ( o0  &  (~ t27)  &  (~ e25) ) ;
 assign b9 = ( (~ a25)  &  (~ v27)  &  (~ c25) ) | ( o0  &  (~ w27)  &  (~ e25) ) ;
 assign c9 = ( (~ a25)  &  (~ y27)  &  (~ c25) ) | ( o0  &  (~ z27)  &  (~ e25) ) ;
 assign d9 = ( (~ a25)  &  (~ b28)  &  (~ c25) ) | ( o0  &  (~ c28)  &  (~ e25) ) ;
 assign e9 = ( (~ a25)  &  (~ e28)  &  (~ c25) ) | ( o0  &  (~ f28)  &  (~ e25) ) ;
 assign f9 = ( (~ h28)  &  (~ i28)  &  (~ j28) ) | ( o0  &  (~ k28)  &  (~ l28) ) ;
 assign g9 = ( x3  &  (~ a29) ) | ( l4  &  (~ a17)  &  (~ a29) ) ;
 assign h9 = ( (~ o0) ) | ( (~ e29) ) | ( y3  &  (~ d29) ) ;
 assign i9 = ( (~ o0) ) | ( (~ j29) ) | ( z3  &  (~ i29) ) ;
 assign j9 = ( (~ q0)  &  o0  &  (~ n29) ) ;
 assign k9 = ( (~ c30) ) | ( (~ x29)  &  (~ y29)  &  (~ z29) ) | ( o0  &  (~ a30)  &  (~ b30) ) ;
 assign l9 = ( (~ m30) ) | ( (~ j30)  &  (~ y29)  &  (~ z29) ) | ( o0  &  (~ k30)  &  (~ l30) ) ;
 assign m9 = ( o0  &  (~ t30)  &  (~ u30) ) | ( (~ n0)  &  o0  &  (~ v30) ) ;
 assign n9 = ( (~ o0) ) | ( (~ c31) ) | ( e4  &  (~ b31) ) ;
 assign o9 = ( (~ o0) ) | ( (~ i31) ) | ( f4  &  (~ h31) ) ;
 assign p9 = ( (~ r31) ) | ( (~ n31)  &  (~ o31)  &  (~ z29) ) | ( o0  &  (~ p31)  &  (~ q31) ) ;
 assign q9 = ( (~ c30) ) | ( (~ y31)  &  (~ a25)  &  (~ z29) ) | ( o0  &  (~ z31)  &  (~ a32) ) ;
 assign r9 = ( i4  &  l4  &  (~ i32) ) | ( n1  &  l4  &  (~ i32) ) ;
 assign s9 = ( (~ k32)  &  (~ l32)  &  (~ j28) ) | ( o0  &  (~ m32)  &  (~ n32) ) ;
 assign t9 = ( (~ c4)  &  (~ b4)  &  (~ a33) ) ;
 assign u9 = ( m1  &  (~ c33) ) ;
 assign v9 = ( (~ g15)  &  (~ e33) ) | ( (~ d33)  &  (~ e33) ) ;
 assign w9 = ( k4  &  (~ a25) ) ;
 assign g15 = ( (~ h35) ) | ( (~ x0)  &  h1  &  (~ g35) ) | ( (~ y0)  &  i1  &  (~ g35) ) ;
 assign j15 = ( c1 ) | ( q0 ) | ( (~ o0) ) ;
 assign k15 = ( (~ t15) ) | ( e1 ) | ( d1 ) ;
 assign l15 = ( (~ h1) ) | ( g1 ) | ( q0 ) ;
 assign m15 = ( t15  &  (~ n0)  &  (~ o15) ) ;
 assign o15 = ( d1  &  e1 ) | ( e1  &  c1 ) ;
 assign t15 = ( (~ l1)  &  (~ k1)  &  (~ p35) ) ;
 assign w15 = ( (~ c1)  &  (~ d1) ) | ( (~ c1)  &  (~ e1) ) | ( d1  &  (~ e1) ) ;
 assign x15 = ( (~ t15) ) | ( e1 ) | ( n0 ) ;
 assign y15 = ( q0 ) | ( (~ o0) ) | ( (~ z15) ) ;
 assign z15 = ( i1 ) | ( (~ n0)  &  (~ e1)  &  t15 ) ;
 assign b16 = ( (~ c1)  &  (~ d1) ) | ( c1  &  (~ e1) ) | ( (~ d1)  &  (~ e1) ) ;
 assign c16 = ( q0 ) | ( (~ o0) ) | ( (~ d16) ) ;
 assign d16 = ( j1 ) | ( (~ n0)  &  (~ e1)  &  t15 ) ;
 assign f16 = ( (~ c1)  &  (~ d1) ) | ( (~ c1)  &  (~ e1) ) | ( (~ d1)  &  (~ e1) ) ;
 assign g16 = ( q0 ) | ( (~ o0) ) | ( (~ h16) ) ;
 assign h16 = ( k1 ) | ( (~ n0)  &  (~ e1)  &  t15 ) ;
 assign j16 = ( c1 ) | ( n0 ) | ( (~ m16) ) ;
 assign l16 = ( q0 ) | ( (~ o0) ) | ( (~ n0)  &  (~ e1)  &  t15 ) ;
 assign m16 = ( t15  &  (~ d1) ) ;
 assign p16 = ( q0 ) | ( (~ o0) ) | ( (~ g15)  &  m1 ) ;
 assign r16 = ( l4  &  (~ o1) ) ;
 assign s16 = ( (~ t15) ) | ( n0 ) ;
 assign u16 = ( (~ l4) ) | ( a17 ) ;
 assign v16 = ( (~ x16) ) | ( (~ n1)  &  (~ t15)  &  (~ w16) ) ;
 assign w16 = ( l4  &  (~ a17) ) ;
 assign x16 = ( j0  &  o0  &  (~ q0) ) | ( n0  &  o0  &  (~ q0) ) | ( (~ t15)  &  o0  &  (~ q0) ) ;
 assign a17 = ( (~ c4)  &  (~ b4)  &  (~ q35) ) ;
 assign b17 = ( l4  &  (~ p1) ) ;
 assign d17 = ( (~ e17) ) | ( (~ o1)  &  (~ t15)  &  (~ w16) ) ;
 assign e17 = ( i0  &  o0  &  (~ q0) ) | ( n0  &  o0  &  (~ q0) ) | ( (~ t15)  &  o0  &  (~ q0) ) ;
 assign g17 = ( l4  &  (~ q1) ) ;
 assign i17 = ( (~ j17) ) | ( (~ p1)  &  (~ t15)  &  (~ w16) ) ;
 assign j17 = ( h0  &  o0  &  (~ q0) ) | ( n0  &  o0  &  (~ q0) ) | ( (~ t15)  &  o0  &  (~ q0) ) ;
 assign l17 = ( l4  &  (~ r1) ) ;
 assign n17 = ( (~ o17) ) | ( (~ q1)  &  (~ t15)  &  (~ w16) ) ;
 assign o17 = ( g0  &  o0  &  (~ q0) ) | ( n0  &  o0  &  (~ q0) ) | ( (~ t15)  &  o0  &  (~ q0) ) ;
 assign q17 = ( l4  &  (~ s1) ) ;
 assign s17 = ( (~ t17) ) | ( (~ r1)  &  (~ t15)  &  (~ w16) ) ;
 assign t17 = ( f0  &  o0  &  (~ q0) ) | ( n0  &  o0  &  (~ q0) ) | ( (~ t15)  &  o0  &  (~ q0) ) ;
 assign v17 = ( l4  &  (~ t1) ) ;
 assign x17 = ( (~ y17) ) | ( (~ s1)  &  (~ t15)  &  (~ w16) ) ;
 assign y17 = ( e0  &  o0  &  (~ q0) ) | ( n0  &  o0  &  (~ q0) ) | ( (~ t15)  &  o0  &  (~ q0) ) ;
 assign a18 = ( l4  &  (~ u1) ) ;
 assign c18 = ( (~ d18) ) | ( (~ t1)  &  (~ t15)  &  (~ w16) ) ;
 assign d18 = ( d0  &  o0  &  (~ q0) ) | ( n0  &  o0  &  (~ q0) ) | ( (~ t15)  &  o0  &  (~ q0) ) ;
 assign f18 = ( l4  &  (~ v1) ) ;
 assign h18 = ( (~ i18) ) | ( (~ u1)  &  (~ t15)  &  (~ w16) ) ;
 assign i18 = ( m0  &  o0  &  (~ q0) ) | ( n0  &  o0  &  (~ q0) ) | ( (~ t15)  &  o0  &  (~ q0) ) ;
 assign k18 = ( l4  &  (~ w1) ) ;
 assign m18 = ( (~ n18) ) | ( (~ v1)  &  (~ t15)  &  (~ w16) ) ;
 assign n18 = ( k0  &  o0  &  (~ q0) ) | ( n0  &  o0  &  (~ q0) ) | ( (~ t15)  &  o0  &  (~ q0) ) ;
 assign p18 = ( l4  &  (~ x1) ) ;
 assign r18 = ( (~ s18) ) | ( (~ w1)  &  (~ t15)  &  (~ w16) ) ;
 assign s18 = ( l0  &  o0  &  (~ q0) ) | ( n0  &  o0  &  (~ q0) ) | ( (~ t15)  &  o0  &  (~ q0) ) ;
 assign u18 = ( l4  &  (~ y1) ) ;
 assign w18 = ( (~ x18) ) | ( (~ x1)  &  (~ t15)  &  (~ w16) ) ;
 assign x18 = ( q  &  o0  &  (~ q0) ) | ( n0  &  o0  &  (~ q0) ) | ( (~ t15)  &  o0  &  (~ q0) ) ;
 assign z18 = ( l4  &  (~ z1) ) ;
 assign b19 = ( (~ c19) ) | ( (~ y1)  &  (~ t15)  &  (~ w16) ) ;
 assign c19 = ( r  &  o0  &  (~ q0) ) | ( n0  &  o0  &  (~ q0) ) | ( (~ t15)  &  o0  &  (~ q0) ) ;
 assign e19 = ( l4  &  (~ a2) ) ;
 assign g19 = ( (~ h19) ) | ( (~ z1)  &  (~ t15)  &  (~ w16) ) ;
 assign h19 = ( s  &  o0  &  (~ q0) ) | ( n0  &  o0  &  (~ q0) ) | ( (~ t15)  &  o0  &  (~ q0) ) ;
 assign j19 = ( l4  &  (~ b2) ) ;
 assign l19 = ( (~ m19) ) | ( (~ a2)  &  (~ t15)  &  (~ w16) ) ;
 assign m19 = ( t  &  o0  &  (~ q0) ) | ( n0  &  o0  &  (~ q0) ) | ( (~ t15)  &  o0  &  (~ q0) ) ;
 assign o19 = ( l4  &  (~ c2) ) ;
 assign q19 = ( (~ r19) ) | ( (~ b2)  &  (~ t15)  &  (~ w16) ) ;
 assign r19 = ( u  &  o0  &  (~ q0) ) | ( n0  &  o0  &  (~ q0) ) | ( (~ t15)  &  o0  &  (~ q0) ) ;
 assign t19 = ( l4  &  (~ d2) ) ;
 assign v19 = ( (~ w19) ) | ( (~ c2)  &  (~ t15)  &  (~ w16) ) ;
 assign w19 = ( v  &  o0  &  (~ q0) ) | ( n0  &  o0  &  (~ q0) ) | ( (~ t15)  &  o0  &  (~ q0) ) ;
 assign y19 = ( l4  &  (~ e2) ) ;
 assign a20 = ( (~ b20) ) | ( (~ d2)  &  (~ t15)  &  (~ w16) ) ;
 assign b20 = ( w  &  o0  &  (~ q0) ) | ( n0  &  o0  &  (~ q0) ) | ( (~ t15)  &  o0  &  (~ q0) ) ;
 assign d20 = ( l4  &  (~ f2) ) ;
 assign f20 = ( (~ g20) ) | ( (~ e2)  &  (~ t15)  &  (~ w16) ) ;
 assign g20 = ( x  &  o0  &  (~ q0) ) | ( n0  &  o0  &  (~ q0) ) | ( (~ t15)  &  o0  &  (~ q0) ) ;
 assign i20 = ( l4  &  (~ g2) ) ;
 assign k20 = ( (~ l20) ) | ( (~ f2)  &  (~ t15)  &  (~ w16) ) ;
 assign l20 = ( y  &  o0  &  (~ q0) ) | ( n0  &  o0  &  (~ q0) ) | ( (~ t15)  &  o0  &  (~ q0) ) ;
 assign n20 = ( l4  &  (~ h2) ) ;
 assign p20 = ( (~ q20) ) | ( (~ g2)  &  (~ t15)  &  (~ w16) ) ;
 assign q20 = ( z  &  o0  &  (~ q0) ) | ( n0  &  o0  &  (~ q0) ) | ( (~ t15)  &  o0  &  (~ q0) ) ;
 assign s20 = ( l4  &  (~ i2) ) ;
 assign u20 = ( (~ v20) ) | ( (~ h2)  &  (~ t15)  &  (~ w16) ) ;
 assign v20 = ( a0  &  o0  &  (~ q0) ) | ( n0  &  o0  &  (~ q0) ) | ( (~ t15)  &  o0  &  (~ q0) ) ;
 assign x20 = ( l4  &  (~ j2) ) ;
 assign z20 = ( (~ a21) ) | ( (~ i2)  &  (~ t15)  &  (~ w16) ) ;
 assign a21 = ( b0  &  o0  &  (~ q0) ) | ( n0  &  o0  &  (~ q0) ) | ( (~ t15)  &  o0  &  (~ q0) ) ;
 assign c21 = ( l4  &  (~ k2) ) ;
 assign e21 = ( (~ f21) ) | ( (~ j2)  &  (~ t15)  &  (~ w16) ) ;
 assign f21 = ( c0  &  o0  &  (~ q0) ) | ( n0  &  o0  &  (~ q0) ) | ( (~ t15)  &  o0  &  (~ q0) ) ;
 assign h21 = ( (~ l21) ) | ( (~ m0)  &  (~ s16)  &  (~ i21) ) | ( (~ a17)  &  (~ j21)  &  (~ k21) ) ;
 assign i21 = ( (~ k0)  &  a ) | ( l0  &  a ) | ( k0  &  (~ l0)  &  i ) ;
 assign j21 = ( (~ l4) ) | ( l2 ) ;
 assign k21 = ( t15  &  (~ n0)  &  (~ m0) ) ;
 assign l21 = ( k2 ) | ( (~ a17)  &  l4 ) | ( (~ m0)  &  (~ n0)  &  t15 ) ;
 assign q21 = ( (~ t21) ) | ( (~ m0)  &  (~ s16)  &  (~ r21) ) | ( (~ a17)  &  (~ s21)  &  (~ k21) ) ;
 assign r21 = ( (~ k0)  &  b ) | ( l0  &  b ) | ( k0  &  (~ l0)  &  j ) ;
 assign s21 = ( (~ l4) ) | ( m2 ) ;
 assign t21 = ( l2 ) | ( (~ a17)  &  l4 ) | ( (~ m0)  &  (~ n0)  &  t15 ) ;
 assign x21 = ( (~ a22) ) | ( (~ m0)  &  (~ s16)  &  (~ y21) ) | ( (~ a17)  &  (~ z21)  &  (~ k21) ) ;
 assign y21 = ( (~ k0)  &  c ) | ( l0  &  c ) | ( k0  &  (~ l0)  &  k ) ;
 assign z21 = ( (~ l4) ) | ( n2 ) ;
 assign a22 = ( m2 ) | ( (~ a17)  &  l4 ) | ( (~ m0)  &  (~ n0)  &  t15 ) ;
 assign e22 = ( (~ h22) ) | ( (~ m0)  &  (~ s16)  &  (~ f22) ) | ( (~ a17)  &  (~ g22)  &  (~ k21) ) ;
 assign f22 = ( (~ k0)  &  d ) | ( l0  &  d ) | ( k0  &  (~ l0)  &  l ) ;
 assign g22 = ( (~ l4) ) | ( o2 ) ;
 assign h22 = ( n2 ) | ( (~ a17)  &  l4 ) | ( (~ m0)  &  (~ n0)  &  t15 ) ;
 assign l22 = ( (~ o22) ) | ( (~ m0)  &  (~ s16)  &  (~ m22) ) | ( (~ a17)  &  (~ n22)  &  (~ k21) ) ;
 assign m22 = ( (~ k0)  &  e ) | ( l0  &  e ) | ( k0  &  (~ l0)  &  m ) ;
 assign n22 = ( (~ l4) ) | ( p2 ) ;
 assign o22 = ( o2 ) | ( (~ a17)  &  l4 ) | ( (~ m0)  &  (~ n0)  &  t15 ) ;
 assign s22 = ( (~ v22) ) | ( (~ m0)  &  (~ s16)  &  (~ t22) ) | ( (~ a17)  &  (~ u22)  &  (~ k21) ) ;
 assign t22 = ( (~ k0)  &  f ) | ( l0  &  f ) | ( k0  &  (~ l0)  &  n ) ;
 assign u22 = ( (~ l4) ) | ( q2 ) ;
 assign v22 = ( p2 ) | ( (~ a17)  &  l4 ) | ( (~ m0)  &  (~ n0)  &  t15 ) ;
 assign z22 = ( (~ c23) ) | ( (~ m0)  &  (~ s16)  &  (~ a23) ) | ( (~ a17)  &  (~ b23)  &  (~ k21) ) ;
 assign a23 = ( (~ k0)  &  g ) | ( l0  &  g ) | ( k0  &  (~ l0)  &  o ) ;
 assign b23 = ( (~ l4) ) | ( r2 ) ;
 assign c23 = ( q2 ) | ( (~ a17)  &  l4 ) | ( (~ m0)  &  (~ n0)  &  t15 ) ;
 assign g23 = ( (~ j23) ) | ( (~ m0)  &  (~ s16)  &  (~ h23) ) | ( (~ a17)  &  (~ i23)  &  (~ k21) ) ;
 assign h23 = ( (~ k0)  &  h ) | ( l0  &  h ) | ( k0  &  (~ l0)  &  p ) ;
 assign i23 = ( (~ l4) ) | ( s2 ) ;
 assign j23 = ( r2 ) | ( (~ a17)  &  l4 ) | ( (~ m0)  &  (~ n0)  &  t15 ) ;
 assign n23 = ( (~ p23)  &  (~ q23) ) | ( (~ s2)  &  a17  &  (~ q23) ) | ( (~ s2)  &  (~ o23)  &  (~ q23) ) | ( (~ a17)  &  (~ o23)  &  (~ q23) ) ;
 assign o23 = ( l4  &  t2 ) ;
 assign p23 = ( n0 ) | ( m0 ) | ( (~ w23) ) ;
 assign q23 = ( i  &  (~ r23)  &  (~ s23) ) | ( (~ l4)  &  s2  &  (~ t23) ) ;
 assign r23 = ( (~ t15) ) | ( n0 ) | ( m0 ) ;
 assign s23 = ( (~ k0)  &  l0 ) | ( k0  &  (~ l0) ) ;
 assign t23 = ( (~ n0)  &  (~ m0)  &  (~ u23) ) ;
 assign u23 = ( (~ t15) ) | ( (~ k0)  &  l0 ) | ( k0  &  (~ l0) ) ;
 assign w23 = ( k0  &  l0  &  t15 ) | ( (~ k0)  &  (~ l0)  &  t15 ) ;
 assign y23 = ( (~ p23)  &  (~ a24) ) | ( (~ t2)  &  a17  &  (~ a24) ) | ( (~ t2)  &  (~ z23)  &  (~ a24) ) | ( (~ a17)  &  (~ z23)  &  (~ a24) ) ;
 assign z23 = ( l4  &  u2 ) ;
 assign a24 = ( j  &  (~ r23)  &  (~ s23) ) | ( (~ l4)  &  t2  &  (~ t23) ) ;
 assign c24 = ( (~ p23)  &  (~ e24) ) | ( (~ u2)  &  a17  &  (~ e24) ) | ( (~ u2)  &  (~ d24)  &  (~ e24) ) | ( (~ a17)  &  (~ d24)  &  (~ e24) ) ;
 assign d24 = ( l4  &  v2 ) ;
 assign e24 = ( k  &  (~ r23)  &  (~ s23) ) | ( (~ l4)  &  u2  &  (~ t23) ) ;
 assign g24 = ( (~ p23)  &  (~ i24) ) | ( (~ v2)  &  a17  &  (~ i24) ) | ( (~ v2)  &  (~ h24)  &  (~ i24) ) | ( (~ a17)  &  (~ h24)  &  (~ i24) ) ;
 assign h24 = ( l4  &  w2 ) ;
 assign i24 = ( l  &  (~ r23)  &  (~ s23) ) | ( (~ l4)  &  v2  &  (~ t23) ) ;
 assign k24 = ( (~ p23)  &  (~ m24) ) | ( (~ w2)  &  a17  &  (~ m24) ) | ( (~ w2)  &  (~ l24)  &  (~ m24) ) | ( (~ a17)  &  (~ l24)  &  (~ m24) ) ;
 assign l24 = ( l4  &  x2 ) ;
 assign m24 = ( m  &  (~ r23)  &  (~ s23) ) | ( (~ l4)  &  w2  &  (~ t23) ) ;
 assign o24 = ( (~ p23)  &  (~ q24) ) | ( (~ x2)  &  a17  &  (~ q24) ) | ( (~ x2)  &  (~ p24)  &  (~ q24) ) | ( (~ a17)  &  (~ p24)  &  (~ q24) ) ;
 assign p24 = ( l4  &  y2 ) ;
 assign q24 = ( n  &  (~ r23)  &  (~ s23) ) | ( (~ l4)  &  x2  &  (~ t23) ) ;
 assign s24 = ( (~ p23)  &  (~ u24) ) | ( (~ y2)  &  a17  &  (~ u24) ) | ( (~ y2)  &  (~ t24)  &  (~ u24) ) | ( (~ a17)  &  (~ t24)  &  (~ u24) ) ;
 assign t24 = ( l4  &  z2 ) ;
 assign u24 = ( o  &  (~ r23)  &  (~ s23) ) | ( (~ l4)  &  y2  &  (~ t23) ) ;
 assign w24 = ( n0 ) | ( m0 ) | ( (~ p) ) ;
 assign x24 = ( (~ t15) ) | ( q0 ) | ( (~ o0) ) ;
 assign y24 = ( (~ z2) ) | ( q0 ) ;
 assign z24 = ( l4  &  (~ a17) ) | ( (~ m0)  &  (~ s16)  &  (~ s23) ) ;
 assign a25 = ( (~ l25) ) | ( q0 ) | ( (~ o0) ) ;
 assign b25 = ( (~ k4) ) | ( (~ b3) ) | ( j25 ) ;
 assign c25 = ( (~ r25) ) | ( h1  &  (~ p25) ) | ( i1  &  (~ q25) ) ;
 assign d25 = ( (~ a3) ) | ( q0 ) ;
 assign e25 = ( (~ h1)  &  (~ i1)  &  (~ h25) ) | ( (~ f25)  &  (~ i1)  &  (~ h25) ) | ( (~ h1)  &  (~ g25)  &  (~ h25) ) | ( (~ f25)  &  (~ g25)  &  (~ h25) ) ;
 assign f25 = ( j1 ) | ( i1 ) | ( (~ o25) ) ;
 assign g25 = ( l1 ) | ( k1 ) | ( j1 ) ;
 assign h25 = ( (~ k4) ) | ( (~ i25) ) | ( l1  &  k1 ) ;
 assign i25 = ( (~ l1)  &  (~ j25)  &  (~ k25) ) | ( (~ j1)  &  (~ j25)  &  (~ k25) ) ;
 assign j25 = ( (~ h4)  &  (~ r35) ) ;
 assign k25 = ( (~ l25) ) | ( (~ m25) ) | ( k1  &  j1 ) ;
 assign l25 = ( (~ x34) ) | ( h1  &  (~ x0) ) | ( i1  &  (~ y0) ) ;
 assign m25 = ( l1 ) | ( k1 ) | ( (~ n25) ) ;
 assign n25 = ( (~ j1)  &  (~ i1)  &  (~ h1) ) ;
 assign o25 = ( (~ l1)  &  (~ k1) ) ;
 assign p25 = ( (~ j1)  &  (~ i1)  &  (~ t25) ) ;
 assign q25 = ( (~ l1)  &  (~ k1)  &  (~ j1) ) ;
 assign r25 = ( i1  &  (~ s25) ) | ( h1  &  (~ s25) ) | ( (~ q25)  &  (~ s25) ) ;
 assign s25 = ( j1  &  k1 ) | ( j1  &  l1 ) | ( k1  &  l1 ) ;
 assign t25 = ( l1 ) | ( k1 ) ;
 assign w25 = ( (~ k4) ) | ( (~ c3) ) | ( j25 ) ;
 assign x25 = ( (~ b3) ) | ( q0 ) ;
 assign z25 = ( (~ k4) ) | ( (~ d3) ) | ( j25 ) ;
 assign a26 = ( (~ c3) ) | ( q0 ) ;
 assign c26 = ( (~ k4) ) | ( (~ e3) ) | ( j25 ) ;
 assign d26 = ( (~ d3) ) | ( q0 ) ;
 assign f26 = ( (~ k4) ) | ( (~ f3) ) | ( j25 ) ;
 assign g26 = ( (~ e3) ) | ( q0 ) ;
 assign i26 = ( (~ k4) ) | ( (~ g3) ) | ( j25 ) ;
 assign j26 = ( (~ f3) ) | ( q0 ) ;
 assign l26 = ( (~ k4) ) | ( (~ h3) ) | ( j25 ) ;
 assign m26 = ( (~ g3) ) | ( q0 ) ;
 assign o26 = ( (~ k4) ) | ( (~ i3) ) | ( j25 ) ;
 assign p26 = ( (~ h3) ) | ( q0 ) ;
 assign r26 = ( (~ k4) ) | ( (~ j3) ) | ( j25 ) ;
 assign s26 = ( (~ i3) ) | ( q0 ) ;
 assign u26 = ( (~ k4) ) | ( (~ k3) ) | ( j25 ) ;
 assign v26 = ( (~ j3) ) | ( q0 ) ;
 assign x26 = ( (~ k4) ) | ( (~ l3) ) | ( j25 ) ;
 assign y26 = ( (~ k3) ) | ( q0 ) ;
 assign a27 = ( (~ k4) ) | ( (~ m3) ) | ( j25 ) ;
 assign b27 = ( (~ l3) ) | ( q0 ) ;
 assign d27 = ( (~ k4) ) | ( (~ n3) ) | ( j25 ) ;
 assign e27 = ( (~ m3) ) | ( q0 ) ;
 assign g27 = ( (~ k4) ) | ( (~ o3) ) | ( j25 ) ;
 assign h27 = ( (~ n3) ) | ( q0 ) ;
 assign j27 = ( (~ k4) ) | ( (~ p3) ) | ( j25 ) ;
 assign k27 = ( (~ o3) ) | ( q0 ) ;
 assign m27 = ( (~ k4) ) | ( (~ q3) ) | ( j25 ) ;
 assign n27 = ( (~ p3) ) | ( q0 ) ;
 assign p27 = ( (~ k4) ) | ( (~ r3) ) | ( j25 ) ;
 assign q27 = ( (~ q3) ) | ( q0 ) ;
 assign s27 = ( (~ k4) ) | ( (~ s3) ) | ( j25 ) ;
 assign t27 = ( (~ r3) ) | ( q0 ) ;
 assign v27 = ( (~ k4) ) | ( (~ t3) ) | ( j25 ) ;
 assign w27 = ( (~ s3) ) | ( q0 ) ;
 assign y27 = ( (~ k4) ) | ( (~ u3) ) | ( j25 ) ;
 assign z27 = ( (~ t3) ) | ( q0 ) ;
 assign b28 = ( (~ k4) ) | ( (~ v3) ) | ( j25 ) ;
 assign c28 = ( (~ u3) ) | ( q0 ) ;
 assign e28 = ( (~ k4) ) | ( (~ w3) ) | ( j25 ) ;
 assign f28 = ( (~ v3) ) | ( q0 ) ;
 assign h28 = ( q0 ) | ( (~ o0) ) ;
 assign i28 = ( (~ k4) ) | ( j25 ) | ( (~ l25) ) ;
 assign j28 = ( (~ s0)  &  h1 ) | ( (~ r28)  &  h1 ) | ( (~ q25)  &  h1 ) | ( (~ s0)  &  (~ s28) ) | ( (~ r28)  &  (~ s28) ) | ( (~ q25)  &  (~ s28) ) ;
 assign k28 = ( (~ w3) ) | ( q0 ) ;
 assign l28 = ( (~ h1)  &  (~ i1)  &  (~ m28) ) | ( (~ f25)  &  (~ i1)  &  (~ m28) ) | ( (~ h1)  &  (~ g25)  &  (~ m28) ) | ( (~ f25)  &  (~ g25)  &  (~ m28) ) ;
 assign m28 = ( (~ k4) ) | ( j25 ) | ( (~ n28) ) ;
 assign n28 = ( (~ l1)  &  l25  &  (~ p28) ) | ( (~ k1)  &  l25  &  (~ p28) ) ;
 assign p28 = ( (~ q28) ) | ( (~ i1)  &  (~ h1)  &  (~ g25) ) ;
 assign q28 = ( (~ j1) ) | ( (~ k1)  &  (~ l1) ) ;
 assign r28 = ( (~ i1)  &  h1 ) ;
 assign s28 = ( (~ i1)  &  (~ u28) ) | ( i1  &  (~ g25)  &  t0 ) ;
 assign u28 = ( (~ u0)  &  (~ w0)  &  (~ w28) ) | ( (~ u0)  &  j1  &  (~ w28) ) | ( (~ w0)  &  (~ j1)  &  (~ w28) ) | ( (~ w0)  &  (~ o25)  &  (~ w28) ) | ( j1  &  (~ o25)  &  (~ w28) ) | ( (~ u0)  &  (~ v28)  &  (~ w28) ) | ( (~ j1)  &  (~ v28)  &  (~ w28) ) | ( (~ o25)  &  (~ v28)  &  (~ w28) ) ;
 assign v28 = ( l1  &  (~ k1) ) ;
 assign w28 = ( (~ l1)  &  (~ x28) ) ;
 assign x28 = ( (~ k1) ) | ( j1 ) | ( (~ v0) ) ;
 assign a29 = ( (~ b29) ) | ( l4  &  x3  &  (~ a17) ) ;
 assign b29 = ( n0  &  o0  &  (~ q0) ) | ( (~ t15)  &  o0  &  (~ q0) ) ;
 assign d29 = ( l4  &  (~ x3)  &  (~ a17) ) ;
 assign e29 = ( (~ t15)  &  (~ q0)  &  (~ f29) ) | ( n0  &  (~ q0)  &  (~ f29) ) ;
 assign f29 = ( l4  &  (~ g29) ) ;
 assign g29 = ( y3 ) | ( x3 ) | ( a17 ) ;
 assign i29 = ( (~ x3)  &  (~ a17)  &  (~ m29) ) ;
 assign j29 = ( (~ t15)  &  (~ q0)  &  (~ k29) ) | ( n0  &  (~ q0)  &  (~ k29) ) ;
 assign k29 = ( l4  &  (~ z3)  &  (~ l29) ) ;
 assign l29 = ( (~ y3) ) | ( x3 ) | ( a17 ) ;
 assign m29 = ( (~ l4) ) | ( (~ y3) ) ;
 assign n29 = ( (~ o29)  &  (~ a4)  &  (~ r29) ) | ( (~ p29)  &  (~ a4)  &  (~ r29) ) | ( (~ s16)  &  (~ a4)  &  (~ r29) ) | ( (~ o29)  &  (~ n0)  &  (~ r29) ) | ( (~ p29)  &  (~ n0)  &  (~ r29) ) | ( (~ s16)  &  (~ n0)  &  (~ r29) ) | ( (~ o29)  &  (~ q29)  &  (~ r29) ) | ( (~ p29)  &  (~ q29)  &  (~ r29) ) | ( (~ s16)  &  (~ q29)  &  (~ r29) ) ;
 assign o29 = ( y3  &  (~ x3)  &  (~ a17) ) ;
 assign p29 = ( l4  &  (~ a4)  &  z3 ) ;
 assign q29 = ( x3 ) | ( a17 ) | ( (~ w29) ) ;
 assign r29 = ( m0  &  a4  &  (~ t29) ) | ( m0  &  t15  &  (~ t29) ) | ( a4  &  (~ t15)  &  (~ t29) ) | ( a4  &  (~ s23)  &  (~ t29) ) | ( t15  &  (~ s23)  &  (~ t29) ) ;
 assign t29 = ( t15  &  n0 ) | ( (~ t15)  &  (~ u29)  &  (~ v29) ) ;
 assign u29 = ( x3 ) | ( a17 ) ;
 assign v29 = ( (~ l4) ) | ( (~ z3) ) | ( (~ y3) ) ;
 assign w29 = ( l4  &  z3  &  y3 ) ;
 assign x29 = ( (~ o0) ) | ( (~ g30) ) | ( (~ h30) ) ;
 assign y29 = ( x3 ) | ( a17 ) | ( q0 ) ;
 assign z29 = ( t15  &  (~ n0) ) ;
 assign a30 = ( (~ b4) ) | ( q0 ) ;
 assign b30 = ( t15  &  (~ n0) ) | ( (~ a17)  &  (~ e30)  &  (~ f30) ) ;
 assign c30 = ( (~ t15) ) | ( q0 ) | ( (~ d30) ) ;
 assign d30 = ( o0  &  (~ n0)  &  m0 ) ;
 assign e30 = ( (~ y3) ) | ( x3 ) ;
 assign f30 = ( (~ l4) ) | ( a4 ) | ( (~ z3) ) ;
 assign g30 = ( z3  &  y3 ) ;
 assign h30 = ( l4  &  (~ b4)  &  (~ a4) ) ;
 assign j30 = ( (~ o0) ) | ( (~ q30) ) | ( (~ r30) ) ;
 assign k30 = ( (~ c4) ) | ( q0 ) ;
 assign l30 = ( t15  &  (~ n0) ) | ( (~ a17)  &  (~ o30)  &  (~ p30) ) ;
 assign m30 = ( (~ t15) ) | ( q0 ) | ( (~ n30) ) ;
 assign n30 = ( o0  &  (~ n0)  &  (~ m0) ) ;
 assign o30 = ( (~ z3) ) | ( (~ y3) ) | ( x3 ) ;
 assign p30 = ( (~ l4) ) | ( b4 ) | ( a4 ) ;
 assign q30 = ( (~ a4)  &  z3  &  y3 ) ;
 assign r30 = ( l4  &  (~ c4)  &  (~ b4) ) ;
 assign t30 = ( g1 ) | ( q0 ) ;
 assign u30 = ( (~ d4)  &  (~ x30) ) | ( (~ j25)  &  l25  &  (~ w30) ) ;
 assign v30 = ( (~ t15) ) | ( q0 ) ;
 assign w30 = ( (~ k4) ) | ( (~ d4) ) ;
 assign x30 = ( k4  &  (~ j25)  &  l25 ) ;
 assign b31 = ( (~ j25)  &  l25  &  (~ f31) ) ;
 assign c31 = ( (~ q0)  &  (~ g1)  &  (~ d31) ) ;
 assign d31 = ( t15  &  (~ n0) ) | ( (~ j25)  &  l25  &  (~ e31) ) ;
 assign e31 = ( (~ k4) ) | ( e4 ) | ( d4 ) ;
 assign f31 = ( (~ k4) ) | ( d4 ) ;
 assign h31 = ( (~ j25)  &  l25  &  (~ m31) ) ;
 assign i31 = ( (~ q0)  &  (~ g1)  &  (~ j31) ) ;
 assign j31 = ( t15  &  (~ n0) ) | ( l25  &  (~ k31)  &  (~ l31) ) ;
 assign k31 = ( d4 ) | ( j25 ) ;
 assign l31 = ( (~ k4) ) | ( f4 ) | ( (~ e4) ) ;
 assign m31 = ( (~ k4) ) | ( (~ e4) ) | ( d4 ) ;
 assign n31 = ( (~ o0) ) | ( (~ v31) ) | ( (~ w31) ) ;
 assign o31 = ( j25 ) | ( (~ l25) ) | ( q0 ) ;
 assign p31 = ( (~ g4) ) | ( g1 ) | ( q0 ) ;
 assign q31 = ( t15  &  (~ n0) ) | ( l25  &  (~ k31)  &  (~ u31) ) ;
 assign r31 = ( (~ t15) ) | ( q0 ) | ( (~ s31) ) ;
 assign s31 = ( o0  &  (~ t31) ) ;
 assign t31 = ( n0 ) | ( (~ k0)  &  l0  &  m0 ) | ( k0  &  (~ l0)  &  m0 ) ;
 assign u31 = ( (~ k4) ) | ( (~ f4) ) | ( (~ e4) ) ;
 assign v31 = ( e4  &  (~ d4)  &  (~ g1) ) ;
 assign w31 = ( k4  &  (~ g4)  &  f4 ) ;
 assign y31 = ( (~ d32) ) | ( (~ e32) ) | ( (~ f32) ) ;
 assign z31 = ( (~ h4) ) | ( g1 ) | ( q0 ) ;
 assign a32 = ( t15  &  (~ n0) ) | ( l25  &  (~ b32)  &  (~ c32) ) ;
 assign b32 = ( (~ e4) ) | ( d4 ) | ( j25 ) ;
 assign c32 = ( (~ k4) ) | ( g4 ) | ( (~ f4) ) ;
 assign d32 = ( (~ g1)  &  (~ j25) ) ;
 assign e32 = ( f4  &  e4  &  (~ d4) ) ;
 assign f32 = ( k4  &  (~ h4)  &  (~ g4) ) ;
 assign i32 = ( (~ j32) ) | ( i4  &  n1 ) ;
 assign j32 = ( (~ a17)  &  (~ q0)  &  o0 ) ;
 assign k32 = ( q0 ) | ( (~ o0) ) | ( (~ y32) ) ;
 assign l32 = ( g1 ) | ( j25 ) | ( (~ l25) ) ;
 assign m32 = ( (~ j4) ) | ( g1 ) | ( q0 ) ;
 assign n32 = ( (~ h1)  &  (~ o32)  &  (~ r32) ) | ( (~ h1)  &  (~ p32)  &  (~ r32) ) | ( h1  &  (~ q32)  &  (~ r32) ) | ( (~ o32)  &  (~ q32)  &  (~ r32) ) | ( (~ p32)  &  (~ q32)  &  (~ r32) ) ;
 assign o32 = ( (~ j1)  &  (~ i1) ) ;
 assign p32 = ( (~ w0)  &  (~ k1) ) | ( (~ v0)  &  (~ l1) ) | ( (~ k1)  &  (~ l1) ) ;
 assign q32 = ( i1 ) | ( (~ s0) ) | ( (~ q25) ) ;
 assign r32 = ( (~ u32) ) | ( i1  &  (~ t32) ) | ( (~ h1)  &  (~ u0)  &  (~ s32) ) ;
 assign s32 = ( l1 ) | ( k1 ) | ( i1 ) ;
 assign t32 = ( (~ j1)  &  t0  &  (~ t25) ) ;
 assign u32 = ( n4  &  k4  &  (~ w32) ) ;
 assign w32 = ( (~ l25) ) | ( (~ x32) ) | ( l1  &  k1 ) ;
 assign x32 = ( (~ j1)  &  (~ j25) ) | ( (~ k1)  &  (~ l1)  &  (~ j25) ) ;
 assign y32 = ( n4  &  k4  &  (~ j4) ) ;
 assign a33 = ( (~ o0) ) | ( (~ b33) ) | ( (~ q30) ) ;
 assign b33 = ( m1  &  (~ q0) ) ;
 assign c33 = ( a17 ) | ( q0 ) | ( (~ o0) ) ;
 assign d33 = ( (~ n4) ) | ( (~ b35) ) | ( h1  &  (~ x0) ) ;
 assign e33 = ( q0 ) | ( (~ o0) ) | ( (~ l25)  &  d33 ) ;
 assign h33 = ( (~ l0)  &  (~ d3) ) | ( l0  &  (~ l3) ) | ( (~ d3)  &  (~ l3) ) ;
 assign i33 = ( l0  &  (~ d3) ) | ( (~ l0)  &  (~ l3) ) | ( (~ d3)  &  (~ l3) ) ;
 assign j33 = ( (~ t3)  &  (~ m0) ) ;
 assign k33 = ( (~ l0)  &  (~ c3) ) | ( l0  &  (~ k3) ) | ( (~ c3)  &  (~ k3) ) ;
 assign l33 = ( l0  &  (~ c3) ) | ( (~ l0)  &  (~ k3) ) | ( (~ c3)  &  (~ k3) ) ;
 assign m33 = ( (~ s3)  &  (~ m0) ) ;
 assign n33 = ( (~ l0)  &  (~ b3) ) | ( l0  &  (~ j3) ) | ( (~ b3)  &  (~ j3) ) ;
 assign o33 = ( l0  &  (~ b3) ) | ( (~ l0)  &  (~ j3) ) | ( (~ b3)  &  (~ j3) ) ;
 assign p33 = ( (~ r3)  &  (~ m0) ) ;
 assign q33 = ( (~ l0)  &  (~ a3) ) | ( l0  &  (~ i3) ) | ( (~ a3)  &  (~ i3) ) ;
 assign r33 = ( l0  &  (~ a3) ) | ( (~ l0)  &  (~ i3) ) | ( (~ a3)  &  (~ i3) ) ;
 assign s33 = ( (~ q3)  &  (~ m0) ) ;
 assign t33 = ( (~ m0) ) | ( k0  &  l0  &  (~ e3) ) | ( (~ k0)  &  (~ l0)  &  (~ e3) ) ;
 assign u33 = ( (~ m0) ) | ( k0  &  l0  &  (~ f3) ) | ( (~ k0)  &  (~ l0)  &  (~ f3) ) ;
 assign v33 = ( (~ m0) ) | ( k0  &  l0  &  (~ g3) ) | ( (~ k0)  &  (~ l0)  &  (~ g3) ) ;
 assign w33 = ( (~ m0) ) | ( k0  &  l0  &  (~ h3) ) | ( (~ k0)  &  (~ l0)  &  (~ h3) ) ;
 assign x33 = ( (~ m0) ) | ( k0  &  l0  &  (~ i3) ) | ( (~ k0)  &  (~ l0)  &  (~ i3) ) ;
 assign y33 = ( (~ m0) ) | ( k0  &  l0  &  (~ j3) ) | ( (~ k0)  &  (~ l0)  &  (~ j3) ) ;
 assign z33 = ( (~ m0) ) | ( k0  &  l0  &  (~ k3) ) | ( (~ k0)  &  (~ l0)  &  (~ k3) ) ;
 assign a34 = ( (~ m0) ) | ( k0  &  l0  &  (~ l3) ) | ( (~ k0)  &  (~ l0)  &  (~ l3) ) ;
 assign b34 = ( (~ k4)  &  h1  &  (~ n0) ) ;
 assign c34 = ( (~ k4)  &  i1  &  (~ n0) ) ;
 assign d34 = ( (~ k4)  &  j1  &  (~ n0) ) ;
 assign e34 = ( (~ k4)  &  k1  &  (~ n0) ) ;
 assign f34 = ( (~ k4)  &  l1  &  (~ n0) ) ;
 assign g34 = ( (~ c4)  &  (~ b4)  &  (~ a4) ) ;
 assign h34 = ( (~ f1)  &  i4 ) | ( f1  &  (~ i4) ) ;
 assign i34 = ( (~ z3) ) | ( (~ y3) ) | ( (~ g34) ) ;
 assign k34 = ( (~ k4)  &  m1  &  h1 ) ;
 assign l34 = ( (~ k4)  &  m1  &  i1 ) ;
 assign m34 = ( (~ k4)  &  m1  &  j1 ) ;
 assign n34 = ( (~ k4)  &  m1  &  k1 ) ;
 assign o34 = ( (~ k4)  &  m1  &  l1 ) ;
 assign p34 = ( l4  &  h1 ) ;
 assign q34 = ( l4  &  i1 ) ;
 assign r34 = ( l4  &  j1 ) ;
 assign s34 = ( l4  &  k1 ) ;
 assign t34 = ( l4  &  l1 ) ;
 assign v34 = ( (~ y3) ) | ( (~ x3) ) | ( (~ w34) ) ;
 assign w34 = ( (~ a4)  &  z3 ) ;
 assign x34 = ( z0  &  a1  &  b1 ) | ( (~ j1)  &  a1  &  b1 ) | ( z0  &  (~ k1)  &  b1 ) | ( (~ j1)  &  (~ k1)  &  b1 ) | ( z0  &  a1  &  (~ l1) ) | ( (~ j1)  &  a1  &  (~ l1) ) | ( z0  &  (~ k1)  &  (~ l1) ) | ( (~ j1)  &  (~ k1)  &  (~ l1) ) ;
 assign b35 = ( (~ i1)  &  (~ j1)  &  (~ d35) ) | ( y0  &  (~ j1)  &  (~ d35) ) | ( (~ i1)  &  z0  &  (~ d35) ) | ( y0  &  z0  &  (~ d35) ) ;
 assign d35 = ( (~ e35) ) | ( k1  &  (~ a1) ) | ( l1  &  (~ b1) ) ;
 assign e35 = ( h4 ) | ( (~ f35) ) ;
 assign f35 = ( (~ g4)  &  f4  &  e4 ) ;
 assign g35 = ( f4  &  e4  &  (~ o35) ) ;
 assign h35 = ( (~ i35)  &  (~ j35) ) | ( (~ j1)  &  (~ k1)  &  (~ j35) ) | ( (~ k1)  &  z0  &  (~ j35) ) | ( (~ j1)  &  a1  &  (~ j35) ) | ( z0  &  a1  &  (~ j35) ) ;
 assign i35 = ( (~ f4) ) | ( (~ e4) ) | ( (~ n35) ) ;
 assign j35 = ( (~ n4)  &  (~ k35) ) | ( (~ i35)  &  (~ k35) ) | ( (~ b1)  &  l1  &  (~ k35) ) ;
 assign k35 = ( (~ h4)  &  (~ g4)  &  (~ l35) ) ;
 assign l35 = ( (~ d4) ) | ( g1 ) | ( (~ m35) ) ;
 assign m35 = ( f4  &  e4 ) ;
 assign n35 = ( (~ h4)  &  (~ g4) ) ;
 assign o35 = ( h4 ) | ( g4 ) ;
 assign p35 = ( j1 ) | ( i1 ) | ( h1 ) ;
 assign q35 = ( (~ y3) ) | ( x3 ) | ( (~ w34) ) ;
 assign r35 = ( g4 ) | ( (~ f4) ) | ( (~ e4) ) ;
 assign t4 = ( u3 ) ;
 assign u4 = ( v3 ) ;
 assign m5 = ( m4 ) ;
 assign m6 = ( k4 ) ;


endmodule

