module k2_2 (
	a, b, c, d, e, f, g, h, 
	i, j, k, l, m, n, o, p, q, r, 
	s, t, u, v, w, x, y, z, a0, b0, 
	c0, d0, e0, f0, g0, h0, i0, j0, k0, l0, 
	m0, n0, o0, p0, q0, r0, s0, t0, u0, v0, 
	w0, x0, y0, z0, a1, b1, c1, d1, e1, f1, 
	g1, h1, i1, j1, k1, l1, m1, n1, o1, p1, 
	q1, r1, s1, t1, u1, v1, w1, x1, y1, z1, 
	a2, b2, c2, d2, e2, f2, g2, h2, i2, j2, 
	k2, l2);

input a, b, c, d, e, f, g, h, i, j, k, l, m, n, o, p, q, r, s, t, u, v, w, x, y, z, a0, b0, c0, d0, e0, f0, g0, h0, i0, j0, k0, l0, m0, n0, o0, p0, q0, r0, s0;

output t0, u0, v0, w0, x0, y0, z0, a1, b1, c1, d1, e1, f1, g1, h1, i1, j1, k1, l1, m1, n1, o1, p1, q1, r1, s1, t1, u1, v1, w1, x1, y1, z1, a2, b2, c2, d2, e2, f2, g2, h2, i2, j2, k2, l2;

wire d5, x5, y5, z5, a6, b6, c6, d6, e6, f6, g6, h6, i6, j6, k6, l6, m6, n6, o6, p6, q6, r6, s6, t6, u6, v6, w6, x6, y6, z6, a7, b7, c7, d7, e7, f7, g7, h7, i7, j7, k7, l7, m7, n7, o7, p7, q7, r7, s7, t7, u7, v7, w7, x7, y7, z7, a8, b8, c8, d8, e8, f8, g8, h8, i8, j8, k8, l8, m8, n8, o8, p8, q8, r8, s8, t8, u8, v8, w8, x8, y8, z8, a9, b9, c9, d9, e9, f9, g9, h9, i9, j9, k9, l9, m9, n9, o9, p9, q9, r9, s9, t9, u9, v9, w9, x9, y9, z9, a10, b10, c10, d10, e10, f10, g10, h10, i10, j10, k10, l10, m10, n10, o10, p10, q10, r10, s10, t10, u10, v10, w10, x10, y10, z10, a11, b11, c11, d11, e11, f11, g11, h11, i11, j11, k11, l11, m11, n11, o11, p11, q11, r11, s11, t11, u11, v11, w11, x11, y11, z11, a12, b12, c12, d12, e12, f12, g12, h12, i12, j12, k12, l12, m12, n12, o12, p12, q12, r12, s12, t12, u12, v12;

assign v0 =((~ a) & a);
 assign j2 =((~ a) & a);
 assign t0 = ( g9 ) | ( l6 ) | ( m9 ) | ( n9 ) | ( e10 ) | ( l11 ) ;
 assign u0 = ( g9 ) | ( l11 ) ;
 assign w0 = ( m9 ) | ( n9 ) ;
 assign x0 = ( l6 ) | ( n9 ) | ( l11 ) ;
 assign y0 = ( h9 ) | ( m6 ) | ( f10 ) | ( t10 ) ;
 assign z0 = ( w8 ) | ( a9 ) | ( b9 ) | ( c9 ) | ( d9 ) | ( i2 ) | ( k10 ) | ( w10 ) | ( z10 ) | ( c11 ) | ( f11 ) | ( t11 ) | ( x11 ) | ( d12 ) | ( k12 ) | ( v12 ) | ( s11 ) | ( u6 ) | ( q12 ) | ( q6 ) | ( s6 ) | ( k6 ) | ( p6 ) | ( e6 ) | ( b6 ) | ( a6 ) | ( z5 ) | ( n8 ) | ( j8 ) | ( g8 ) ;
 assign a1 = ( a9 ) | ( b9 ) | ( w10 ) | ( z10 ) | ( p6 ) | ( e6 ) ;
 assign b1 = ( w8 ) | ( a9 ) | ( c9 ) | ( i2 ) | ( k10 ) | ( w10 ) | ( c11 ) | ( t11 ) | ( k12 ) | ( s11 ) | ( s6 ) | ( k6 ) | ( e6 ) | ( z5 ) | ( j8 ) ;
 assign c1 = ( x11 ) | ( d12 ) | ( g8 ) ;
 assign d1 = ( x8 ) | ( e9 ) | ( f9 ) | ( i9 ) | ( o9 ) | ( p9 ) | ( o6 ) | ( y9 ) | ( g10 ) | ( l10 ) | ( x10 ) | ( a11 ) | ( d11 ) | ( e11 ) | ( g11 ) | ( h11 ) | ( x9 ) | ( u11 ) | ( y11 ) | ( d7 ) | ( l12 ) | ( n12 ) | ( i12 ) | ( u12 ) | ( r11 ) | ( g12 ) | ( n1 ) | ( o1 ) | ( j6 ) | ( g6 ) | ( f6 ) | ( y5 ) | ( m8 ) | ( i8 ) | ( f8 ) | ( d8 ) | ( z7 ) | ( y7 ) | ( x7 ) | ( w7 ) | ( v7 ) | ( u7 ) | ( t7 ) | ( q7 ) ;
 assign e1 = ( x8 ) | ( y8 ) | ( e9 ) | ( f9 ) | ( i9 ) | ( j9 ) | ( o9 ) | ( p9 ) | ( r9 ) | ( s9 ) | ( o6 ) | ( t6 ) | ( y9 ) | ( z9 ) | ( g10 ) | ( h10 ) | ( l10 ) | ( m10 ) | ( x10 ) | ( y10 ) | ( b11 ) | ( d11 ) | ( e11 ) | ( g11 ) | ( h11 ) | ( x9 ) | ( u11 ) | ( y11 ) | ( d7 ) | ( l12 ) | ( u12 ) | ( g12 ) | ( r6 ) | ( f6 ) | ( d6 ) | ( m8 ) | ( h8 ) | ( f8 ) | ( o7 ) ;
 assign f1 = ( x8 ) | ( y8 ) | ( e9 ) | ( f9 ) | ( i9 ) | ( j9 ) | ( r9 ) | ( s9 ) | ( o6 ) | ( t6 ) | ( y9 ) | ( z9 ) | ( g10 ) | ( h10 ) | ( l10 ) | ( m10 ) | ( x10 ) | ( y10 ) | ( a11 ) | ( b11 ) | ( d11 ) | ( e11 ) | ( g11 ) | ( h11 ) | ( l9 ) | ( t9 ) | ( x9 ) | ( b10 ) | ( u11 ) | ( y11 ) | ( d7 ) | ( l12 ) | ( n12 ) | ( i12 ) | ( u12 ) | ( r11 ) | ( g12 ) | ( r6 ) | ( n1 ) | ( o1 ) | ( j6 ) | ( g6 ) | ( f6 ) | ( d6 ) | ( y5 ) | ( m8 ) | ( i8 ) | ( h8 ) | ( f8 ) | ( d8 ) | ( q7 ) | ( p7 ) ;
 assign g1 = ( r8 ) | ( u8 ) | ( o9 ) | ( p9 ) | ( a11 ) | ( l9 ) | ( t9 ) | ( b10 ) | ( p11 ) | ( c12 ) | ( m12 ) | ( n12 ) | ( v10 ) | ( i12 ) | ( j12 ) | ( p12 ) | ( s12 ) | ( o12 ) | ( r11 ) | ( o11 ) | ( y6 ) | ( x6 ) | ( w6 ) | ( v6 ) | ( r6 ) | ( n1 ) | ( o1 ) | ( n6 ) | ( j6 ) | ( h6 ) | ( g6 ) | ( c6 ) | ( d6 ) | ( y5 ) | ( e12 ) | ( i8 ) | ( h8 ) | ( z7 ) | ( w7 ) | ( v7 ) | ( u7 ) | ( t7 ) | ( q7 ) ;
 assign h1 = ( f9 ) | ( p9 ) | ( t6 ) | ( z9 ) | ( a11 ) | ( e11 ) | ( h11 ) | ( t9 ) | ( n12 ) | ( i12 ) | ( o12 ) | ( r11 ) | ( o11 ) | ( r6 ) | ( n1 ) | ( o1 ) | ( j6 ) | ( g6 ) | ( d6 ) | ( y5 ) | ( i8 ) | ( h8 ) | ( c8 ) | ( z7 ) | ( x7 ) | ( v7 ) | ( t7 ) | ( r7 ) ;
 assign i1 = ( r8 ) | ( u8 ) | ( x8 ) | ( e9 ) | ( i9 ) | ( o9 ) | ( p9 ) | ( o6 ) | ( y9 ) | ( f10 ) | ( g10 ) | ( i10 ) | ( l10 ) | ( x10 ) | ( a11 ) | ( d11 ) | ( g11 ) | ( x9 ) | ( c10 ) | ( d10 ) | ( u11 ) | ( x11 ) | ( y11 ) | ( z11 ) | ( d7 ) | ( q11 ) | ( f12 ) | ( k12 ) | ( l12 ) | ( m12 ) | ( n12 ) | ( i12 ) | ( t12 ) | ( u12 ) | ( r11 ) | ( u9 ) | ( w6 ) | ( g12 ) | ( n1 ) | ( o1 ) | ( j6 ) | ( g6 ) | ( c6 ) | ( f6 ) | ( y5 ) | ( o8 ) | ( m8 ) | ( k8 ) | ( i8 ) | ( g8 ) | ( f8 ) | ( e8 ) | ( s7 ) | ( o7 ) | ( n7 ) | ( m7 ) | ( l7 ) | ( j7 ) | ( i7 ) | ( g7 ) ;
 assign j1 = ( r8 ) | ( u8 ) | ( e9 ) | ( a11 ) | ( d11 ) | ( g11 ) | ( c10 ) | ( d10 ) | ( x11 ) | ( d5 ) | ( a12 ) | ( q11 ) | ( f12 ) | ( k12 ) | ( n12 ) | ( i12 ) | ( p12 ) | ( s12 ) | ( t12 ) | ( o12 ) | ( r11 ) | ( o11 ) | ( u9 ) | ( y6 ) | ( w6 ) | ( v6 ) | ( r6 ) | ( n1 ) | ( o1 ) | ( n6 ) | ( j6 ) | ( h6 ) | ( g6 ) | ( c6 ) | ( d6 ) | ( y5 ) | ( e12 ) | ( q8 ) | ( o8 ) | ( m8 ) | ( k8 ) | ( i8 ) | ( h8 ) | ( g8 ) | ( e8 ) | ( d8 ) | ( z7 ) | ( y7 ) | ( x7 ) | ( w7 ) | ( v7 ) | ( u7 ) | ( t7 ) | ( q7 ) ;
 assign k1 = ( r8 ) | ( u8 ) | ( x8 ) | ( y8 ) | ( e9 ) | ( f9 ) | ( i9 ) | ( j9 ) | ( o9 ) | ( p9 ) | ( r9 ) | ( s9 ) | ( o6 ) | ( t6 ) | ( y9 ) | ( z9 ) | ( g10 ) | ( h10 ) | ( j10 ) | ( l10 ) | ( m10 ) | ( x10 ) | ( y10 ) | ( a11 ) | ( b11 ) | ( e11 ) | ( h11 ) | ( i11 ) | ( l9 ) | ( t9 ) | ( x9 ) | ( b10 ) | ( u11 ) | ( y11 ) | ( z11 ) | ( d7 ) | ( l12 ) | ( m12 ) | ( p12 ) | ( u12 ) | ( o12 ) | ( r11 ) | ( o11 ) | ( y6 ) | ( x6 ) | ( w6 ) | ( g12 ) | ( r6 ) | ( n1 ) | ( o1 ) | ( j6 ) | ( g6 ) | ( c6 ) | ( f6 ) | ( d6 ) | ( y5 ) | ( q8 ) | ( i8 ) | ( f8 ) | ( e8 ) | ( c8 ) | ( s7 ) | ( r7 ) | ( p7 ) | ( o7 ) | ( n7 ) | ( h7 ) | ( g7 ) ;
 assign l1 = ( r8 ) | ( u8 ) | ( x8 ) | ( i9 ) | ( o9 ) | ( p9 ) | ( o6 ) | ( y9 ) | ( f10 ) | ( g10 ) | ( j10 ) | ( l10 ) | ( x10 ) | ( x9 ) | ( p11 ) | ( u11 ) | ( y11 ) | ( z11 ) | ( c12 ) | ( d7 ) | ( l12 ) | ( m12 ) | ( n12 ) | ( v10 ) | ( i12 ) | ( j12 ) | ( p12 ) | ( s12 ) | ( u12 ) | ( b7 ) | ( y6 ) | ( v6 ) | ( g12 ) | ( n6 ) | ( h6 ) | ( f6 ) | ( e12 ) | ( h8 ) | ( f8 ) | ( e8 ) | ( j7 ) | ( i7 ) | ( h7 ) | ( g7 ) ;
 assign m1 = ( x8 ) | ( e9 ) | ( i9 ) | ( o9 ) | ( p9 ) | ( o6 ) | ( y9 ) | ( f10 ) | ( g10 ) | ( l10 ) | ( x10 ) | ( d11 ) | ( g11 ) | ( x9 ) | ( p11 ) | ( u11 ) | ( y11 ) | ( d5 ) | ( a12 ) | ( c12 ) | ( d7 ) | ( l12 ) | ( m12 ) | ( v10 ) | ( i12 ) | ( j12 ) | ( p12 ) | ( u12 ) | ( o12 ) | ( o11 ) | ( x6 ) | ( w6 ) | ( v6 ) | ( g12 ) | ( r6 ) | ( n6 ) | ( h6 ) | ( c6 ) | ( f6 ) | ( d6 ) | ( e12 ) | ( m8 ) | ( h8 ) | ( f8 ) | ( e8 ) | ( s7 ) | ( o7 ) | ( l7 ) | ( k7 ) | ( i7 ) ;
 assign n1 = ( (~ r)  &  s  &  (~ t)  &  u  &  (~ v)  &  a0  &  (~ c0)  &  d0  &  e0 ) ;
 assign o1 = ( s  &  (~ t)  &  u  &  (~ v)  &  a0  &  c0  &  d0  &  (~ e0) ) ;
 assign p1 = ( r8 ) | ( x8 ) | ( y8 ) | ( z8 ) | ( e9 ) | ( f9 ) | ( i9 ) | ( j9 ) | ( o9 ) | ( p9 ) | ( q9 ) | ( r9 ) | ( s9 ) | ( o6 ) | ( t6 ) | ( y9 ) | ( z9 ) | ( f10 ) | ( g10 ) | ( h10 ) | ( i10 ) | ( j10 ) | ( l10 ) | ( m10 ) | ( r10 ) | ( s10 ) | ( x10 ) | ( y10 ) | ( a11 ) | ( b11 ) | ( d11 ) | ( e11 ) | ( g11 ) | ( h11 ) | ( i11 ) | ( l9 ) | ( t9 ) | ( k11 ) | ( x9 ) | ( b10 ) | ( p11 ) | ( c10 ) | ( d10 ) | ( u11 ) | ( x11 ) | ( d5 ) | ( z11 ) | ( a12 ) | ( c12 ) | ( d7 ) | ( q11 ) | ( f12 ) | ( k12 ) | ( m12 ) | ( n12 ) | ( v10 ) | ( i12 ) | ( j12 ) | ( p12 ) | ( s12 ) | ( t12 ) | ( u12 ) | ( o12 ) | ( r11 ) | ( o11 ) | ( u9 ) | ( b7 ) | ( z6 ) | ( y6 ) | ( x6 ) | ( w6 ) | ( v6 ) | ( g12 ) | ( r6 ) | ( n1 ) | ( o1 ) | ( n6 ) | ( j6 ) | ( i6 ) | ( h6 ) | ( g6 ) | ( c6 ) | ( f6 ) | ( d6 ) | ( y5 ) | ( e12 ) | ( q8 ) | ( o8 ) | ( m8 ) | ( k8 ) | ( i8 ) | ( h8 ) | ( g8 ) | ( f8 ) | ( e8 ) | ( d8 ) | ( c8 ) | ( z7 ) | ( y7 ) | ( x7 ) | ( w7 ) | ( v7 ) | ( u7 ) | ( t7 ) | ( s7 ) | ( r7 ) | ( q7 ) | ( p7 ) | ( o7 ) | ( n7 ) | ( m7 ) | ( l7 ) | ( k7 ) | ( j7 ) | ( i7 ) | ( h7 ) | ( g7 ) ;
 assign q1 = ( e9 ) | ( d11 ) | ( g11 ) ;
 assign d5 = ( (~ s)  &  (~ t)  &  u  &  (~ v)  &  w  &  (~ d0)  &  e0 ) ;
 assign s1 = ( u8 ) | ( z8 ) | ( q9 ) | ( r10 ) | ( s10 ) | ( k11 ) | ( m11 ) | ( p11 ) | ( d5 ) | ( z11 ) | ( b12 ) | ( c12 ) | ( m12 ) | ( v10 ) | ( j12 ) | ( p12 ) | ( s12 ) | ( q10 ) | ( b7 ) | ( z6 ) | ( y6 ) | ( x6 ) | ( w6 ) | ( v6 ) | ( n6 ) | ( i6 ) | ( h6 ) | ( c6 ) | ( e12 ) | ( n7 ) ;
 assign t1 = ( p11 ) | ( c12 ) | ( j12 ) | ( e12 ) ;
 assign u1 = ( c10 ) | ( d10 ) | ( x11 ) | ( q11 ) | ( f12 ) | ( k12 ) | ( t12 ) | ( u9 ) | ( o8 ) | ( k8 ) | ( g8 ) ;
 assign v1 = ( y8 ) | ( z8 ) | ( f9 ) | ( j9 ) | ( q9 ) | ( r9 ) | ( s9 ) | ( t6 ) | ( v9 ) | ( a7 ) | ( k9 ) | ( j10 ) | ( p10 ) | ( x5 ) | ( r10 ) | ( s10 ) | ( e7 ) | ( u10 ) | ( b11 ) | ( h11 ) | ( i11 ) | ( l9 ) | ( t9 ) | ( k11 ) | ( m11 ) | ( b10 ) | ( d5 ) | ( a12 ) | ( b12 ) | ( q10 ) | ( b7 ) | ( z6 ) | ( s7 ) | ( p7 ) | ( m7 ) | ( l7 ) | ( k7 ) | ( j7 ) | ( i7 ) | ( h7 ) | ( g7 ) | ( f7 ) ;
 assign w1 = ( w8 ) | ( a9 ) | ( b9 ) | ( c9 ) | ( d9 ) | ( h9 ) | ( m6 ) | ( i2 ) | ( f10 ) | ( k10 ) | ( w10 ) | ( z10 ) | ( c11 ) | ( f11 ) | ( t10 ) | ( t11 ) | ( x11 ) | ( d12 ) | ( k12 ) | ( v12 ) | ( u6 ) | ( b6 ) | ( n8 ) | ( g8 ) ;
 assign x1 = ( s11 ) | ( q12 ) | ( k6 ) | ( p6 ) | ( e6 ) | ( j8 ) ;
 assign y1 = ( s11 ) | ( q6 ) | ( s6 ) | ( a6 ) | ( z5 ) | ( j8 ) ;
 assign z1 = ( (~ m)  &  (~ n)  &  (~ o)  &  v  &  (~ b0)  &  (~ c0)  &  (~ d0)  &  (~ e0) ) ;
 assign a2 = ( o8 ) | ( k8 ) | ( i8 ) | ( g8 ) | ( f8 ) ;
 assign b2 = ( l6 ) | ( m9 ) | ( n9 ) | ( m6 ) | ( o6 ) | ( z9 ) | ( h10 ) | ( i10 ) | ( m10 ) | ( y10 ) | ( e11 ) | ( u11 ) | ( v11 ) | ( x11 ) | ( d7 ) | ( j11 ) | ( k12 ) | ( u12 ) | ( r12 ) | ( o12 ) | ( s11 ) | ( o11 ) | ( g12 ) | ( r6 ) | ( q6 ) | ( s6 ) | ( f6 ) | ( d6 ) | ( a6 ) | ( z5 ) | ( n8 ) | ( m8 ) | ( l8 ) | ( j8 ) | ( c8 ) | ( b8 ) | ( a8 ) | ( z7 ) | ( y7 ) | ( x7 ) | ( w7 ) | ( v7 ) | ( t7 ) | ( r7 ) | ( q7 ) | ( o7 ) ;
 assign c2 = ( w8 ) | ( x8 ) | ( a9 ) | ( b9 ) | ( c9 ) | ( d9 ) | ( e9 ) | ( h9 ) | ( i9 ) | ( o9 ) | ( p9 ) | ( m6 ) | ( o6 ) | ( i2 ) | ( y9 ) | ( f10 ) | ( g10 ) | ( k10 ) | ( l10 ) | ( w10 ) | ( x10 ) | ( z10 ) | ( a11 ) | ( c11 ) | ( d11 ) | ( f11 ) | ( g11 ) | ( t10 ) | ( x9 ) | ( p11 ) | ( t11 ) | ( w11 ) | ( x11 ) | ( z11 ) | ( c12 ) | ( d12 ) | ( h12 ) | ( n11 ) | ( k12 ) | ( m12 ) | ( v10 ) | ( j12 ) | ( v12 ) | ( o12 ) | ( s11 ) | ( r11 ) | ( o11 ) | ( w6 ) | ( v6 ) | ( u6 ) | ( q12 ) | ( q6 ) | ( s6 ) | ( n6 ) | ( k6 ) | ( h6 ) | ( p6 ) | ( e6 ) | ( c6 ) | ( b6 ) | ( a6 ) | ( z5 ) | ( e12 ) | ( q8 ) | ( o8 ) | ( l8 ) | ( k8 ) | ( j8 ) | ( h8 ) | ( f8 ) | ( d8 ) | ( u7 ) | ( n7 ) ;
 assign d2 = ( s8 ) | ( t8 ) | ( v8 ) | ( z1 ) | ( x8 ) | ( e9 ) | ( i9 ) | ( l6 ) | ( m9 ) | ( n9 ) | ( o6 ) | ( w9 ) | ( y9 ) | ( a10 ) | ( c7 ) | ( g10 ) | ( i10 ) | ( l10 ) | ( n10 ) | ( o10 ) | ( p8 ) | ( x10 ) | ( y10 ) | ( a11 ) | ( d11 ) | ( g11 ) | ( x9 ) | ( t11 ) | ( v11 ) | ( d12 ) | ( j11 ) | ( v12 ) | ( r12 ) | ( s11 ) | ( u6 ) | ( q12 ) | ( r6 ) | ( k6 ) | ( p6 ) | ( e6 ) | ( b6 ) | ( d6 ) | ( q8 ) | ( m8 ) | ( j8 ) | ( h8 ) | ( g8 ) | ( c8 ) | ( u7 ) | ( r7 ) ;
 assign e2 = ( r8 ) | ( s8 ) | ( t8 ) | ( v8 ) | ( z1 ) | ( w8 ) | ( x8 ) | ( y8 ) | ( z8 ) | ( a9 ) | ( b9 ) | ( c9 ) | ( d9 ) | ( e9 ) | ( f9 ) | ( h9 ) | ( i9 ) | ( j9 ) | ( l6 ) | ( m9 ) | ( n9 ) | ( o9 ) | ( p9 ) | ( q9 ) | ( r9 ) | ( s9 ) | ( m6 ) | ( o6 ) | ( t6 ) | ( v9 ) | ( w9 ) | ( i2 ) | ( y9 ) | ( z9 ) | ( a10 ) | ( a7 ) | ( c7 ) | ( k9 ) | ( f10 ) | ( g10 ) | ( h10 ) | ( i10 ) | ( j10 ) | ( k10 ) | ( l10 ) | ( m10 ) | ( n10 ) | ( o10 ) | ( p10 ) | ( x5 ) | ( r10 ) | ( s10 ) | ( e7 ) | ( u10 ) | ( p8 ) | ( w10 ) | ( x10 ) | ( y10 ) | ( z10 ) | ( a11 ) | ( b11 ) | ( c11 ) | ( d11 ) | ( e11 ) | ( f11 ) | ( g11 ) | ( h11 ) | ( i11 ) | ( l9 ) | ( t9 ) | ( k11 ) | ( m11 ) | ( t10 ) | ( x9 ) | ( b10 ) | ( p11 ) | ( c10 ) | ( d10 ) | ( t11 ) | ( u11 ) | ( v11 ) | ( w11 ) | ( x11 ) | ( y11 ) | ( d5 ) | ( z11 ) | ( a12 ) | ( b12 ) | ( c12 ) | ( d12 ) | ( d7 ) | ( j11 ) | ( h12 ) | ( n11 ) | ( q11 ) | ( f12 ) | ( k12 ) | ( l12 ) | ( m12 ) | ( n12 ) | ( v10 ) | ( i12 ) | ( j12 ) | ( p12 ) | ( s12 ) | ( t12 ) | ( v12 ) | ( u12 ) | ( r12 ) | ( o12 ) | ( s11 ) | ( r11 ) | ( o11 ) | ( u9 ) | ( q10 ) | ( b7 ) | ( z6 ) | ( y6 ) | ( x6 ) | ( w6 ) | ( v6 ) | ( u6 ) | ( g12 ) | ( q12 ) | ( r6 ) | ( n1 ) | ( q6 ) | ( s6 ) | ( o1 ) | ( n6 ) | ( k6 ) | ( j6 ) | ( i6 ) | ( h6 ) | ( p6 ) | ( e6 ) | ( g6 ) | ( c6 ) | ( b6 ) | ( f6 ) | ( d6 ) | ( a6 ) | ( z5 ) | ( y5 ) | ( e12 ) | ( q8 ) | ( o8 ) | ( n8 ) | ( m8 ) | ( l8 ) | ( k8 ) | ( j8 ) | ( i8 ) | ( h8 ) | ( g8 ) | ( f8 ) | ( e8 ) | ( d8 ) | ( c8 ) | ( b8 ) | ( a8 ) | ( z7 ) | ( y7 ) | ( x7 ) | ( w7 ) | ( v7 ) | ( u7 ) | ( t7 ) | ( s7 ) | ( r7 ) | ( q7 ) | ( p7 ) | ( o7 ) | ( n7 ) | ( m7 ) | ( l7 ) | ( k7 ) | ( j7 ) | ( i7 ) | ( h7 ) | ( g7 ) | ( f7 ) | ( s  &  t  &  u  &  v  &  a0  &  e0 ) ;
 assign f2 = ( g9 ) | ( e10 ) | ( l11 ) | ( (~ s)  &  t  &  v  &  c0  &  (~ d0)  &  e0  &  (~ a) ) | ( (~ b)  &  (~ s)  &  t  &  (~ u)  &  (~ v)  &  w  &  d0  &  (~ e0) ) | ( (~ s)  &  (~ t)  &  u  &  v  &  w  &  (~ d0)  &  e0  &  (~ a) ) | ( s  &  t  &  (~ u)  &  (~ v)  &  w  &  d0  &  (~ e0)  &  (~ a) ) | ( (~ s)  &  (~ t)  &  u  &  v  &  (~ d0)  &  e0  &  (~ a)  &  a0 ) | ( (~ s)  &  (~ t)  &  u  &  v  &  (~ d0)  &  e0  &  (~ a)  &  z ) | ( s  &  t  &  (~ u)  &  (~ v)  &  d0  &  (~ e0)  &  (~ a)  &  z ) | ( s  &  t  &  u  &  (~ v)  &  (~ d0)  &  (~ a)  &  d  &  b0 ) | ( (~ b)  &  (~ s)  &  t  &  (~ u)  &  (~ v)  &  d0  &  (~ e0)  &  x ) | ( (~ b)  &  (~ s)  &  t  &  (~ u)  &  v  &  w  &  (~ c0)  &  (~ d0)  &  e0 ) | ( (~ s)  &  t  &  u  &  (~ v)  &  w  &  c0  &  d0  &  (~ e0)  &  (~ a) ) | ( s  &  t  &  (~ u)  &  (~ v)  &  c0  &  (~ d0)  &  e0  &  (~ a)  &  a0 ) | ( s  &  t  &  (~ u)  &  (~ v)  &  (~ c0)  &  d0  &  (~ e0)  &  (~ a)  &  a0 ) | ( (~ b)  &  (~ s)  &  t  &  (~ u)  &  v  &  (~ c0)  &  (~ d0)  &  e0  &  x ) | ( (~ s)  &  (~ t)  &  u  &  (~ v)  &  (~ c0)  &  d0  &  (~ e0)  &  (~ a)  &  x ) | ( s  &  (~ t)  &  u  &  (~ v)  &  c0  &  (~ d0)  &  e0  &  (~ a)  &  a0  &  l ) | ( s  &  (~ t)  &  u  &  (~ v)  &  (~ c0)  &  d0  &  (~ e0)  &  (~ a)  &  a0  &  r ) | ( s  &  (~ t)  &  u  &  (~ v)  &  (~ c0)  &  d0  &  (~ e0)  &  (~ a)  &  a0  &  (~ r) ) | ( s  &  t  &  u  &  (~ v)  &  c0  &  d0  &  (~ e0)  &  (~ a)  &  (~ b0)  &  (~ e) ) | ( (~ s)  &  t  &  u  &  (~ v)  &  w  &  (~ c0)  &  d0  &  (~ e0)  &  (~ a)  &  (~ f) ) | ( (~ s)  &  (~ t)  &  (~ u)  &  (~ v)  &  (~ c0)  &  d0  &  (~ e0)  &  (~ a)  &  (~ d)  &  (~ f) ) | ( s  &  t  &  u  &  (~ v)  &  (~ c0)  &  d0  &  e0  &  (~ a)  &  (~ b0)  &  (~ f) ) | ( s  &  (~ t)  &  u  &  v  &  (~ c0)  &  (~ d0)  &  e0  &  (~ a)  &  (~ f)  &  (~ p) ) | ( (~ s)  &  (~ t)  &  u  &  (~ v)  &  c0  &  (~ d0)  &  e0  &  (~ a)  &  (~ d)  &  c ) | ( (~ s)  &  (~ t)  &  (~ u)  &  (~ v)  &  c0  &  (~ d0)  &  e0  &  (~ a)  &  (~ d)  &  (~ c) ) | ( (~ s)  &  t  &  u  &  v  &  w  &  (~ c0)  &  (~ d0)  &  e0  &  (~ a)  &  (~ f)  &  (~ p) ) ;
 assign g2 = ( x8 ) | ( e9 ) | ( i9 ) | ( o9 ) | ( p9 ) | ( o6 ) | ( y9 ) | ( g10 ) | ( l10 ) | ( x10 ) | ( a11 ) | ( d11 ) | ( g11 ) | ( x9 ) | ( y11 ) | ( d7 ) | ( l12 ) | ( n12 ) | ( i12 ) | ( t12 ) | ( u9 ) | ( n1 ) | ( o1 ) | ( j6 ) | ( g6 ) | ( y5 ) | ( k8 ) | ( f8 ) ;
 assign h2 = ( v9 ) | ( p10 ) | ( x5 ) | ( c10 ) | ( d10 ) | ( t12 ) | ( o8 ) ;
 assign i2 = ( a  &  (~ f)  &  (~ p)  &  (~ s)  &  t  &  u  &  v  &  w  &  (~ c0)  &  (~ d0)  &  e0 ) ;
 assign k2 = ( d5 ) | ( z11 ) ;
 assign x5 = ( f  &  k  &  s  &  (~ t)  &  u  &  v  &  z  &  (~ c0)  &  (~ d0)  &  e0 ) ;
 assign y5 = ( s  &  t  &  (~ u)  &  (~ v)  &  a0  &  c0  &  d0  &  (~ e0) ) ;
 assign z5 = ( a  &  (~ l)  &  s  &  t  &  (~ u)  &  (~ v)  &  a0  &  c0  &  (~ d0)  &  e0 ) ;
 assign a6 = ( a  &  l  &  s  &  t  &  (~ u)  &  (~ v)  &  a0  &  c0  &  (~ d0)  &  e0 ) ;
 assign b6 = ( a  &  s  &  t  &  (~ u)  &  (~ v)  &  a0  &  (~ c0)  &  d0  &  (~ e0) ) ;
 assign c6 = ( s  &  t  &  (~ u)  &  (~ v)  &  a0  &  (~ c0)  &  (~ d0)  &  e0 ) ;
 assign d6 = ( s  &  t  &  (~ u)  &  (~ v)  &  a0  &  c0  &  (~ d0)  &  (~ e0) ) ;
 assign e6 = ( a  &  k  &  (~ l)  &  s  &  t  &  (~ u)  &  (~ v)  &  z  &  d0  &  (~ e0) ) ;
 assign f6 = ( s  &  t  &  (~ u)  &  (~ v)  &  a0  &  (~ c0)  &  d0  &  e0 ) ;
 assign g6 = ( s  &  t  &  (~ u)  &  (~ v)  &  z  &  d0  &  e0 ) ;
 assign h6 = ( k  &  s  &  t  &  (~ u)  &  (~ v)  &  z  &  (~ d0)  &  e0 ) ;
 assign i6 = ( (~ k)  &  s  &  t  &  (~ u)  &  (~ v)  &  z  &  (~ d0)  &  e0 ) ;
 assign j6 = ( s  &  t  &  (~ u)  &  (~ v)  &  w  &  d0  &  e0 ) ;
 assign k6 = ( a  &  s  &  t  &  (~ u)  &  (~ v)  &  w  &  d0  &  (~ e0) ) ;
 assign l6 = ( (~ s)  &  t  &  v  &  y  &  (~ c0)  &  (~ d0)  &  e0 ) ;
 assign m6 = ( a  &  (~ s)  &  t  &  v  &  c0  &  (~ d0)  &  e0 ) ;
 assign n6 = ( s  &  t  &  (~ u)  &  (~ v)  &  w  &  (~ d0)  &  e0 ) ;
 assign o6 = ( (~ s)  &  t  &  v  &  c0  &  d0  &  (~ e0) ) ;
 assign p6 = ( a  &  k  &  l  &  s  &  t  &  (~ u)  &  (~ v)  &  z  &  d0  &  (~ e0) ) ;
 assign q6 = ( a  &  (~ l)  &  s  &  (~ t)  &  u  &  (~ v)  &  a0  &  c0  &  (~ d0)  &  e0 ) ;
 assign r6 = ( r  &  s  &  (~ t)  &  u  &  (~ v)  &  a0  &  c0  &  (~ d0)  &  (~ e0) ) ;
 assign s6 = ( a  &  l  &  s  &  (~ t)  &  u  &  (~ v)  &  a0  &  c0  &  (~ d0)  &  e0 ) ;
 assign t6 = ( (~ s)  &  t  &  v  &  c0  &  d0  &  e0 ) ;
 assign u6 = ( a  &  r  &  s  &  (~ t)  &  u  &  (~ v)  &  a0  &  (~ c0)  &  d0  &  (~ e0) ) ;
 assign v6 = ( (~ r)  &  s  &  (~ t)  &  u  &  (~ v)  &  a0  &  (~ c0)  &  (~ d0)  &  e0 ) ;
 assign w6 = ( r  &  s  &  (~ t)  &  u  &  (~ v)  &  a0  &  (~ c0)  &  (~ d0)  &  e0 ) ;
 assign x6 = ( s  &  (~ t)  &  u  &  (~ v)  &  x  &  e0 ) ;
 assign y6 = ( s  &  (~ t)  &  u  &  (~ v)  &  w  &  e0 ) ;
 assign z6 = ( (~ k)  &  s  &  (~ t)  &  (~ u)  &  (~ v)  &  z  &  e0 ) ;
 assign a7 = ( i  &  q  &  (~ s)  &  t  &  u  &  v  &  w  &  c0  &  (~ d0)  &  (~ e0) ) ;
 assign b7 = ( k  &  s  &  (~ t)  &  (~ u)  &  (~ v)  &  z  &  e0 ) ;
 assign c7 = ( (~ h)  &  (~ q)  &  (~ s)  &  t  &  u  &  v  &  w  &  c0  &  (~ d0)  &  (~ e0) ) ;
 assign d7 = ( (~ s)  &  (~ t)  &  u  &  (~ v)  &  (~ c0)  &  d0  &  e0 ) ;
 assign e7 = ( i  &  q  &  s  &  (~ t)  &  u  &  v  &  c0 ) ;
 assign f7 = ( (~ s)  &  (~ t)  &  (~ u)  &  v  &  x  &  d0  &  (~ e0)  &  (~ f0)  &  (~ g0)  &  (~ h0)  &  (~ i0)  &  (~ j0)  &  (~ k0)  &  (~ l0) ) ;
 assign g7 = ( (~ s)  &  (~ t)  &  (~ u)  &  v  &  x  &  d0  &  (~ e0)  &  (~ f0)  &  (~ g0)  &  (~ h0)  &  (~ i0)  &  (~ j0)  &  (~ k0)  &  l0 ) ;
 assign h7 = ( (~ s)  &  (~ t)  &  (~ u)  &  v  &  x  &  d0  &  (~ e0)  &  (~ f0)  &  (~ g0)  &  (~ h0)  &  (~ i0)  &  (~ j0)  &  k0 ) ;
 assign i7 = ( (~ s)  &  (~ t)  &  (~ u)  &  v  &  x  &  d0  &  (~ e0)  &  (~ f0)  &  (~ g0)  &  (~ h0)  &  (~ i0)  &  j0 ) ;
 assign j7 = ( (~ s)  &  (~ t)  &  (~ u)  &  v  &  x  &  d0  &  (~ e0)  &  (~ f0)  &  (~ g0)  &  (~ h0)  &  i0 ) ;
 assign k7 = ( (~ s)  &  (~ t)  &  (~ u)  &  v  &  x  &  d0  &  (~ e0)  &  (~ f0)  &  (~ g0)  &  h0 ) ;
 assign l7 = ( (~ s)  &  (~ t)  &  (~ u)  &  v  &  x  &  d0  &  (~ e0)  &  (~ f0)  &  g0 ) ;
 assign m7 = ( (~ s)  &  (~ t)  &  (~ u)  &  v  &  x  &  d0  &  (~ e0)  &  f0 ) ;
 assign n7 = ( (~ s)  &  (~ t)  &  (~ u)  &  v  &  x  &  (~ d0)  &  e0 ) ;
 assign o7 = ( (~ j)  &  (~ s)  &  (~ t)  &  (~ u)  &  v  &  w  &  (~ c0)  &  d0  &  (~ e0)  &  (~ m0)  &  (~ n0)  &  (~ o0)  &  (~ p0)  &  (~ q0)  &  r0  &  (~ s0) ) ;
 assign p7 = ( (~ j)  &  (~ s)  &  (~ t)  &  (~ u)  &  v  &  w  &  (~ c0)  &  d0  &  (~ e0)  &  (~ m0)  &  (~ n0)  &  (~ o0)  &  (~ p0)  &  (~ q0)  &  (~ r0)  &  (~ s0) ) ;
 assign q7 = ( (~ j)  &  (~ s)  &  (~ t)  &  (~ u)  &  v  &  w  &  (~ c0)  &  d0  &  (~ e0)  &  (~ m0)  &  (~ n0)  &  (~ o0)  &  (~ p0)  &  (~ q0)  &  (~ r0)  &  s0 ) ;
 assign r7 = ( (~ j)  &  (~ s)  &  (~ t)  &  (~ u)  &  v  &  w  &  (~ c0)  &  d0  &  (~ e0)  &  (~ m0)  &  (~ n0)  &  o0  &  (~ p0)  &  (~ q0) ) ;
 assign s7 = ( (~ s)  &  (~ t)  &  (~ u)  &  v  &  w  &  c0  &  e0 ) ;
 assign t7 = ( (~ s)  &  (~ t)  &  (~ u)  &  v  &  w  &  (~ c0)  &  d0  &  e0 ) ;
 assign u7 = ( (~ j)  &  (~ s)  &  (~ t)  &  (~ u)  &  v  &  w  &  (~ c0)  &  d0  &  (~ e0)  &  (~ m0)  &  n0  &  (~ p0)  &  q0 ) ;
 assign v7 = ( (~ j)  &  (~ s)  &  (~ t)  &  (~ u)  &  v  &  w  &  (~ c0)  &  d0  &  (~ e0)  &  (~ m0)  &  n0  &  (~ p0)  &  (~ q0) ) ;
 assign w7 = ( (~ j)  &  (~ s)  &  (~ t)  &  (~ u)  &  v  &  w  &  (~ c0)  &  d0  &  (~ e0)  &  (~ m0)  &  (~ n0)  &  (~ p0)  &  q0 ) ;
 assign x7 = ( (~ j)  &  (~ s)  &  (~ t)  &  (~ u)  &  v  &  w  &  (~ c0)  &  d0  &  (~ e0)  &  (~ m0)  &  p0 ) ;
 assign y7 = ( (~ j)  &  (~ s)  &  (~ t)  &  (~ u)  &  v  &  w  &  (~ c0)  &  d0  &  (~ e0)  &  m0 ) ;
 assign z7 = ( j  &  (~ s)  &  (~ t)  &  (~ u)  &  v  &  w  &  (~ c0)  &  (~ d0)  &  e0  &  (~ f0)  &  (~ h0)  &  n0 ) ;
 assign a8 = ( j  &  (~ s)  &  (~ t)  &  (~ u)  &  v  &  w  &  (~ c0)  &  (~ d0)  &  e0  &  (~ f0)  &  (~ h0)  &  (~ n0) ) ;
 assign b8 = ( j  &  (~ s)  &  (~ t)  &  (~ u)  &  v  &  w  &  (~ c0)  &  (~ d0)  &  e0  &  f0 ) ;
 assign c8 = ( j  &  (~ s)  &  (~ t)  &  (~ u)  &  v  &  w  &  (~ c0)  &  (~ d0)  &  e0  &  h0 ) ;
 assign d8 = ( (~ j)  &  (~ s)  &  (~ t)  &  (~ u)  &  v  &  w  &  (~ c0)  &  (~ d0)  &  e0 ) ;
 assign e8 = ( s  &  t  &  u  &  (~ v)  &  b0  &  (~ c0)  &  d0  &  (~ e0) ) ;
 assign f8 = ( s  &  t  &  u  &  (~ v)  &  b0  &  (~ d0)  &  e0 ) ;
 assign g8 = ( a  &  d  &  s  &  t  &  u  &  (~ v)  &  b0  &  (~ d0)  &  (~ e0) ) ;
 assign h8 = ( (~ d)  &  s  &  t  &  u  &  (~ v)  &  b0  &  (~ d0)  &  (~ e0) ) ;
 assign i8 = ( s  &  t  &  u  &  (~ v)  &  (~ b0)  &  c0  &  d0  &  e0 ) ;
 assign j8 = ( (~ a)  &  (~ e)  &  s  &  t  &  u  &  (~ v)  &  (~ b0)  &  c0  &  d0  &  (~ e0) ) ;
 assign k8 = ( e  &  s  &  t  &  u  &  (~ v)  &  (~ b0)  &  c0  &  d0  &  (~ e0) ) ;
 assign l8 = ( s  &  t  &  u  &  (~ v)  &  (~ b0)  &  c0  &  (~ d0)  &  e0 ) ;
 assign m8 = ( s  &  t  &  u  &  (~ v)  &  (~ b0)  &  c0  &  (~ d0)  &  (~ e0) ) ;
 assign n8 = ( a  &  (~ f)  &  s  &  t  &  u  &  (~ v)  &  (~ b0)  &  (~ c0)  &  d0  &  e0 ) ;
 assign o8 = ( f  &  s  &  t  &  u  &  (~ v)  &  (~ b0)  &  (~ c0)  &  d0  &  e0 ) ;
 assign p8 = ( (~ i)  &  q  &  s  &  (~ t)  &  u  &  v  &  c0 ) ;
 assign q8 = ( s  &  t  &  u  &  (~ v)  &  (~ b0)  &  (~ c0)  &  d0  &  (~ e0) ) ;
 assign r8 = ( o  &  (~ b0)  &  (~ c0)  &  (~ d0)  &  (~ e0) ) ;
 assign s8 = ( (~ o)  &  (~ s)  &  (~ t)  &  u  &  (~ v)  &  (~ x)  &  (~ b0)  &  (~ c0)  &  (~ d0)  &  (~ e0) ) ;
 assign t8 = ( (~ o)  &  s  &  (~ t)  &  (~ u)  &  (~ v)  &  (~ b0)  &  (~ c0)  &  (~ d0)  &  (~ e0) ) ;
 assign u8 = ( n  &  (~ o)  &  v  &  (~ b0)  &  (~ c0)  &  (~ d0)  &  (~ e0) ) ;
 assign v8 = ( n  &  (~ o)  &  (~ v)  &  (~ b0)  &  (~ c0)  &  (~ d0)  &  (~ e0) ) ;
 assign w8 = ( a  &  (~ s)  &  (~ t)  &  u  &  v  &  w  &  (~ d0)  &  e0 ) ;
 assign x8 = ( (~ s)  &  (~ t)  &  u  &  v  &  (~ a0)  &  d0  &  (~ e0) ) ;
 assign y8 = ( (~ s)  &  (~ t)  &  u  &  v  &  (~ a0)  &  d0  &  e0 ) ;
 assign z8 = ( (~ k)  &  (~ s)  &  (~ t)  &  u  &  v  &  z ) ;
 assign a9 = ( a  &  k  &  (~ l)  &  (~ s)  &  (~ t)  &  u  &  v  &  z  &  (~ d0)  &  e0 ) ;
 assign b9 = ( a  &  k  &  l  &  (~ s)  &  (~ t)  &  u  &  v  &  z  &  (~ d0)  &  e0 ) ;
 assign c9 = ( a  &  (~ l)  &  (~ s)  &  (~ t)  &  u  &  v  &  a0  &  (~ d0)  &  e0 ) ;
 assign d9 = ( a  &  l  &  (~ s)  &  (~ t)  &  u  &  v  &  a0  &  (~ d0)  &  e0 ) ;
 assign e9 = ( (~ s)  &  (~ t)  &  u  &  v  &  a0  &  d0  &  (~ e0) ) ;
 assign f9 = ( (~ s)  &  (~ t)  &  u  &  v  &  a0  &  d0  &  e0 ) ;
 assign g9 = ( (~ a)  &  (~ s)  &  (~ t)  &  u  &  v  &  y  &  (~ d0)  &  e0 ) ;
 assign h9 = ( a  &  (~ s)  &  (~ t)  &  u  &  v  &  y  &  (~ d0)  &  e0 ) ;
 assign i9 = ( (~ s)  &  (~ t)  &  u  &  v  &  y  &  d0  &  (~ e0) ) ;
 assign j9 = ( (~ s)  &  (~ t)  &  u  &  v  &  y  &  d0  &  e0 ) ;
 assign k9 = ( h  &  (~ q)  &  (~ s)  &  t  &  u  &  v  &  w  &  c0  &  (~ d0)  &  (~ e0) ) ;
 assign l9 = ( k  &  s  &  t  &  (~ u)  &  v  &  z  &  e0 ) ;
 assign m9 = ( k  &  (~ s)  &  t  &  v  &  z  &  (~ c0)  &  (~ d0)  &  e0 ) ;
 assign n9 = ( (~ s)  &  t  &  v  &  a0  &  (~ c0)  &  (~ d0)  &  e0 ) ;
 assign o9 = ( b  &  (~ s)  &  t  &  (~ u)  &  v  &  w  &  (~ c0)  &  (~ d0)  &  e0 ) ;
 assign p9 = ( b  &  (~ s)  &  t  &  (~ u)  &  v  &  x  &  (~ c0)  &  (~ d0)  &  e0 ) ;
 assign q9 = ( (~ k)  &  (~ s)  &  t  &  v  &  z  &  (~ c0)  &  (~ d0)  &  e0 ) ;
 assign r9 = ( (~ s)  &  t  &  (~ u)  &  v  &  w  &  (~ c0)  &  d0  &  (~ e0) ) ;
 assign s9 = ( (~ s)  &  t  &  (~ u)  &  v  &  x  &  (~ c0)  &  d0  &  (~ e0) ) ;
 assign t9 = ( s  &  t  &  (~ u)  &  v  &  a0  &  e0 ) ;
 assign u9 = ( c  &  (~ d)  &  (~ s)  &  t  &  u  &  (~ v)  &  w  &  c0  &  (~ d0)  &  e0 ) ;
 assign v9 = ( f  &  (~ s)  &  t  &  u  &  v  &  w  &  (~ c0)  &  (~ d0)  &  e0 ) ;
 assign w9 = ( (~ f)  &  p  &  (~ s)  &  t  &  u  &  v  &  w  &  (~ c0)  &  (~ d0)  &  e0 ) ;
 assign x9 = ( s  &  t  &  u  &  v  &  d0  &  (~ e0) ) ;
 assign y9 = ( (~ s)  &  t  &  u  &  v  &  w  &  (~ c0)  &  d0  &  (~ e0) ) ;
 assign z9 = ( (~ s)  &  t  &  u  &  v  &  w  &  (~ c0)  &  d0  &  e0 ) ;
 assign a10 = ( (~ i)  &  q  &  (~ s)  &  t  &  u  &  v  &  w  &  c0  &  (~ d0)  &  (~ e0) ) ;
 assign b10 = ( s  &  t  &  u  &  v  &  d0  &  e0 ) ;
 assign c10 = ( d  &  (~ s)  &  (~ t)  &  (~ u)  &  (~ v)  &  (~ c0)  &  d0  &  (~ e0) ) ;
 assign d10 = ( (~ d)  &  f  &  (~ s)  &  (~ t)  &  (~ u)  &  (~ v)  &  (~ c0)  &  d0  &  (~ e0) ) ;
 assign e10 = ( (~ a)  &  s  &  (~ t)  &  (~ u)  &  v  &  (~ c0)  &  (~ d0)  &  e0 ) ;
 assign f10 = ( a  &  s  &  (~ t)  &  (~ u)  &  v  &  (~ c0)  &  (~ d0)  &  e0 ) ;
 assign g10 = ( s  &  (~ t)  &  (~ u)  &  v  &  (~ c0)  &  d0  &  (~ e0) ) ;
 assign h10 = ( s  &  (~ t)  &  (~ u)  &  v  &  (~ c0)  &  d0  &  e0 ) ;
 assign i10 = ( s  &  (~ t)  &  (~ u)  &  v  &  c0  &  (~ d0)  &  (~ e0) ) ;
 assign j10 = ( s  &  (~ t)  &  (~ u)  &  v  &  c0  &  (~ d0)  &  e0 ) ;
 assign k10 = ( a  &  (~ f)  &  (~ p)  &  s  &  (~ t)  &  u  &  v  &  w  &  (~ c0)  &  (~ d0)  &  e0 ) ;
 assign l10 = ( s  &  (~ t)  &  u  &  v  &  w  &  (~ c0)  &  d0  &  (~ e0) ) ;
 assign m10 = ( s  &  (~ t)  &  u  &  v  &  w  &  (~ c0)  &  d0  &  e0 ) ;
 assign n10 = ( (~ f)  &  p  &  s  &  (~ t)  &  u  &  v  &  (~ c0)  &  (~ d0)  &  e0 ) ;
 assign o10 = ( (~ h)  &  (~ q)  &  s  &  (~ t)  &  u  &  v  &  c0 ) ;
 assign p10 = ( f  &  s  &  (~ t)  &  u  &  v  &  (~ z)  &  (~ c0)  &  (~ d0)  &  e0 ) ;
 assign q10 = ( s  &  (~ t)  &  (~ u)  &  (~ v)  &  w  &  e0 ) ;
 assign r10 = ( f  &  (~ k)  &  s  &  (~ t)  &  u  &  v  &  z  &  (~ c0)  &  (~ d0)  &  e0 ) ;
 assign s10 = ( a  &  (~ f)  &  (~ k)  &  (~ p)  &  s  &  (~ t)  &  u  &  v  &  z  &  (~ c0)  &  (~ d0)  &  e0 ) ;
 assign t10 = ( a  &  s  &  t  &  u  &  v  &  (~ d0)  &  e0 ) ;
 assign u10 = ( h  &  (~ q)  &  s  &  (~ t)  &  u  &  v  &  c0 ) ;
 assign v10 = ( (~ s)  &  t  &  (~ u)  &  (~ v)  &  x  &  (~ d0)  &  e0 ) ;
 assign w10 = ( a  &  (~ f)  &  k  &  (~ l)  &  (~ p)  &  s  &  (~ t)  &  u  &  v  &  z  &  (~ c0)  &  (~ d0)  &  e0 ) ;
 assign x10 = ( (~ l)  &  s  &  (~ t)  &  u  &  v  &  z  &  (~ c0)  &  d0  &  (~ e0) ) ;
 assign y10 = ( (~ l)  &  s  &  (~ t)  &  u  &  v  &  z  &  (~ c0)  &  d0  &  e0 ) ;
 assign z10 = ( a  &  (~ f)  &  k  &  l  &  (~ p)  &  s  &  (~ t)  &  u  &  v  &  z  &  (~ c0)  &  (~ d0)  &  e0 ) ;
 assign a11 = ( l  &  s  &  (~ t)  &  u  &  v  &  z  &  (~ c0)  &  d0  &  (~ e0) ) ;
 assign b11 = ( l  &  s  &  (~ t)  &  u  &  v  &  z  &  (~ c0)  &  d0  &  e0 ) ;
 assign c11 = ( a  &  (~ f)  &  (~ l)  &  (~ p)  &  s  &  (~ t)  &  u  &  v  &  a0  &  (~ c0)  &  (~ d0)  &  e0 ) ;
 assign d11 = ( (~ l)  &  s  &  (~ t)  &  u  &  v  &  a0  &  (~ c0)  &  d0  &  (~ e0) ) ;
 assign e11 = ( (~ l)  &  s  &  (~ t)  &  u  &  v  &  a0  &  (~ c0)  &  d0  &  e0 ) ;
 assign f11 = ( a  &  (~ f)  &  l  &  (~ p)  &  s  &  (~ t)  &  u  &  v  &  a0  &  (~ c0)  &  (~ d0)  &  e0 ) ;
 assign g11 = ( l  &  s  &  (~ t)  &  u  &  v  &  a0  &  (~ c0)  &  d0  &  (~ e0) ) ;
 assign h11 = ( l  &  s  &  (~ t)  &  u  &  v  &  a0  &  (~ c0)  &  d0  &  e0 ) ;
 assign i11 = ( s  &  t  &  (~ u)  &  v  &  w  &  e0 ) ;
 assign j11 = ( (~ s)  &  (~ t)  &  u  &  (~ v)  &  c0  &  (~ d0)  &  (~ e0) ) ;
 assign k11 = ( (~ k)  &  s  &  t  &  (~ u)  &  v  &  z  &  e0 ) ;
 assign l11 = ( (~ a)  &  s  &  t  &  u  &  v  &  y  &  (~ d0)  &  e0 ) ;
 assign m11 = ( s  &  t  &  u  &  v  &  w  &  e0 ) ;
 assign n11 = ( (~ c)  &  (~ d)  &  (~ g)  &  (~ s)  &  (~ t)  &  u  &  (~ v)  &  c0  &  (~ d0)  &  e0 ) ;
 assign o11 = ( (~ c)  &  (~ d)  &  (~ s)  &  t  &  u  &  (~ v)  &  w  &  c0  &  (~ d0)  &  e0 ) ;
 assign p11 = ( (~ s)  &  (~ t)  &  (~ u)  &  (~ v)  &  (~ c0)  &  (~ d0)  &  e0 ) ;
 assign q11 = ( d  &  g  &  (~ s)  &  (~ t)  &  u  &  (~ v)  &  c0  &  (~ d0)  &  e0 ) ;
 assign r11 = ( (~ s)  &  t  &  u  &  (~ v)  &  w  &  c0  &  d0  &  e0 ) ;
 assign s11 = ( a  &  (~ s)  &  t  &  u  &  (~ v)  &  w  &  c0  &  d0  &  (~ e0) ) ;
 assign t11 = ( a  &  (~ d)  &  (~ f)  &  (~ s)  &  (~ t)  &  (~ u)  &  (~ v)  &  (~ c0)  &  d0  &  (~ e0) ) ;
 assign u11 = ( (~ s)  &  (~ t)  &  (~ u)  &  (~ v)  &  (~ c0)  &  d0  &  e0 ) ;
 assign v11 = ( (~ s)  &  (~ t)  &  (~ u)  &  (~ v)  &  c0  &  (~ d0)  &  (~ e0) ) ;
 assign w11 = ( (~ c)  &  (~ d)  &  (~ s)  &  (~ t)  &  (~ u)  &  (~ v)  &  c0  &  (~ d0)  &  e0 ) ;
 assign x11 = ( a  &  c  &  (~ d)  &  (~ s)  &  (~ t)  &  (~ u)  &  (~ v)  &  c0  &  (~ d0)  &  e0 ) ;
 assign y11 = ( (~ s)  &  (~ t)  &  (~ u)  &  (~ v)  &  c0  &  d0  &  (~ e0) ) ;
 assign z11 = ( (~ s)  &  (~ t)  &  u  &  (~ v)  &  y  &  (~ d0)  &  e0 ) ;
 assign a12 = ( (~ s)  &  (~ t)  &  u  &  (~ v)  &  y  &  d0  &  (~ e0) ) ;
 assign b12 = ( (~ s)  &  (~ t)  &  u  &  (~ v)  &  a0  &  (~ d0)  &  e0 ) ;
 assign c12 = ( (~ s)  &  (~ t)  &  u  &  (~ v)  &  x  &  (~ c0)  &  (~ d0)  &  e0 ) ;
 assign d12 = ( a  &  (~ s)  &  (~ t)  &  u  &  (~ v)  &  x  &  (~ c0)  &  d0  &  (~ e0) ) ;
 assign e12 = ( s  &  t  &  u  &  (~ v)  &  (~ b0)  &  (~ c0)  &  (~ d0)  &  e0 ) ;
 assign f12 = ( (~ c)  &  (~ d)  &  g  &  (~ s)  &  (~ t)  &  u  &  (~ v)  &  c0  &  (~ d0)  &  e0 ) ;
 assign g12 = ( r  &  s  &  (~ t)  &  u  &  (~ v)  &  a0  &  (~ c0)  &  d0  &  (~ e0) ) ;
 assign h12 = ( d  &  (~ g)  &  (~ s)  &  (~ t)  &  u  &  (~ v)  &  c0  &  (~ d0)  &  e0 ) ;
 assign i12 = ( b  &  (~ s)  &  t  &  (~ u)  &  (~ v)  &  x  &  d0  &  (~ e0) ) ;
 assign j12 = ( (~ s)  &  t  &  u  &  (~ v)  &  w  &  (~ c0)  &  (~ d0)  &  e0 ) ;
 assign k12 = ( a  &  (~ c)  &  (~ d)  &  (~ s)  &  (~ t)  &  u  &  (~ v)  &  c0  &  (~ d0)  &  e0 ) ;
 assign l12 = ( (~ s)  &  (~ t)  &  u  &  (~ v)  &  c0  &  d0  &  (~ e0) ) ;
 assign m12 = ( (~ s)  &  t  &  (~ u)  &  (~ v)  &  w  &  (~ d0)  &  e0 ) ;
 assign n12 = ( b  &  (~ s)  &  t  &  (~ u)  &  (~ v)  &  w  &  d0  &  (~ e0) ) ;
 assign o12 = ( d  &  (~ s)  &  t  &  u  &  (~ v)  &  w  &  c0  &  (~ d0)  &  e0 ) ;
 assign p12 = ( (~ s)  &  t  &  u  &  (~ v)  &  x  &  (~ c0)  &  (~ d0)  &  e0 ) ;
 assign q12 = ( a  &  (~ r)  &  s  &  (~ t)  &  u  &  (~ v)  &  a0  &  (~ c0)  &  d0  &  (~ e0) ) ;
 assign r12 = ( (~ s)  &  t  &  u  &  (~ v)  &  w  &  c0  &  (~ d0)  &  (~ e0) ) ;
 assign s12 = ( (~ s)  &  t  &  u  &  (~ v)  &  a0  &  (~ c0)  &  (~ d0)  &  e0 ) ;
 assign t12 = ( f  &  (~ s)  &  t  &  u  &  (~ v)  &  w  &  (~ c0)  &  d0  &  (~ e0) ) ;
 assign u12 = ( (~ s)  &  t  &  u  &  (~ v)  &  w  &  (~ c0)  &  d0  &  e0 ) ;
 assign v12 = ( a  &  (~ f)  &  (~ s)  &  t  &  u  &  (~ v)  &  w  &  (~ c0)  &  d0  &  (~ e0) ) ;
 assign r1 = ( d5 ) ;
 assign l2 = ( d5 ) ;


endmodule

