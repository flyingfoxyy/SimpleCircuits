module ex1010_mapped (
	i_9_, i_7_, i_8_, i_5_, i_6_, i_3_, i_4_, i_1_, 
	i_2_, i_0_, o_1_, o_2_, o_0_, o_9_, o_7_, o_8_, o_5_, o_6_, 
	o_3_, o_4_);

input i_9_, i_7_, i_8_, i_5_, i_6_, i_3_, i_4_, i_1_, i_2_, i_0_;

output o_1_, o_2_, o_0_, o_9_, o_7_, o_8_, o_5_, o_6_, o_3_, o_4_;

wire n_n1005, n_n1004, wire12040, wire12041, wire12585, wire12586, wire12588, wire12589, n_n621, n_n620, wire13136, wire13147, n_n3986, wire13572, wire13573, n_n3253, wire14216, wire14222, n_n3622, wire14777, wire14778, wire14779, n_n2525, n_n2523, wire15299, wire15300, n_n2898, wire15816, wire15817, n_n1784, wire16323, wire16324, wire16830, wire16831, n_n1038, wire11502, n_n1014, n_n942, n_n941, n_n937, wire11745, n_n4309, n_n1012, wire11832, n_n1007, n_n1009, wire12036, wire12037, n_n1456, n_n1455, wire12197, wire12200, n_n1396, n_n1415, wire12223, wire12224, wire12247, n_n1397, n_n1418, wire12432, n_n1398, wire25, n_n473, n_n65, n_n5305, wire15, n_n482, n_n5293, wire19, n_n526, n_n5296, n_n522, n_n491, n_n5284, n_n559, wire12601, n_n543, n_n4379, n_n4399, wire12699, wire12700, n_n562, n_n4458, n_n4488, wire12706, wire12707, n_n561, n_n4350, n_n4331, wire12713, wire12714, n_n563, wire22, n_n5297, n_n4378, n_n4408, wire13622, wire13623, n_n3936, n_n3931, n_n3929, wire13643, wire13644, n_n3920, n_n4362, n_n4312, wire13674, wire13679, n_n3194, wire13714, wire13728, wire13729, n_n3187, n_n3202, wire13760, n_n3192, n_n3201, wire13767, wire13768, wire13782, n_n3191, n_n3629, wire14513, wire14514, wire14540, n_n3635, wire14614, n_n3624, n_n3639, wire14655, wire14684, n_n3641, wire14750, wire14751, wire14772, n_n3626, n_n524, n_n464, wire148, n_n2548, wire14935, n_n2530, n_n2551, wire15006, n_n2531, n_n2533, wire15150, wire15151, wire15169, n_n2528, wire15206, n_n4436, n_n4417, wire15307, wire15308, n_n2845, n_n4355, n_n4335, wire15321, wire15322, n_n2846, n_n2841, wire15328, n_n2827, n_n2837, n_n2824, n_n2835, wire15400, n_n2821, n_n2839, wire15412, wire15413, wire15418, n_n2826, n_n2929, wire15437, wire15438, wire15463, n_n2907, wire15501, wire15502, wire15504, n_n2906, n_n2934, wire15543, wire15544, wire15549, n_n2908, n_n2905, wire15743, wire16025, wire16028, n_n1793, n_n1813, n_n1812, wire16072, n_n1792, n_n1818, wire16086, wire16087, wire16114, n_n1794, n_n1789, n_n1790, wire16240, wire16241, n_n1797, wire16263, n_n1787, wire16316, wire16318, n_n1786, n_n4404, n_n4413, wire16475, wire16476, n_n2104, wire16492, wire16493, wire16494, wire16497, n_n2087, n_n2099, wire16503, wire16504, wire16516, n_n2086, n_n2190, wire16545, n_n2166, n_n4367, n_n4374, wire16651, wire16745, wire16763, wire16, n_n518, n_n4338, wire21, n_n536, n_n4339, n_n4337, n_n4401, n_n4403, n_n4400, wire13, n_n4464, n_n455, n_n4467, wire11, n_n4463, wire10, n_n532, n_n4666, wire24, n_n390, n_n4667, n_n534, n_n4664, n_n509, n_n325, n_n4737, wire14, n_n4738, n_n4735, n_n528, n_n4782, n_n4784, n_n4779, wire17, n_n535, n_n4830, n_n260, n_n4831, n_n4900, n_n520, n_n4902, n_n4898, wire18, n_n4976, n_n195, n_n4977, n_n4975, n_n5038, n_n5040, n_n5034, wire12, n_n5092, wire20, n_n130, n_n5093, n_n5091, n_n4440, n_n4434, n_n4432, wire98, wire233, wire236, n_n4720, n_n4718, n_n4717, n_n4857, n_n4862, n_n4856, wire40, wire102, wire245, n_n4991, n_n4996, n_n4992, n_n4995, n_n4990, n_n4998, wire23, n_n4999, n_n500, wire103, n_n4617, n_n4637, n_n4613, n_n4927, n_n4958, n_n4920, n_n4325, n_n4327, n_n4324, n_n4382, n_n4383, n_n530, n_n4380, n_n4923, n_n4924, n_n4921, n_n4982, n_n4983, n_n4981, n_n5035, n_n5032, n_n5111, n_n5112, n_n5109, n_n5171, n_n5174, n_n5167, n_n4597, n_n4598, n_n4602, n_n4593, n_n4601, wire108, n_n4744, n_n4754, n_n4757, n_n4749, n_n4756, wire109, n_n4887, n_n4888, n_n4885, n_n3450, n_n4882, n_n4884, n_n4883, n_n5026, n_n5027, n_n5025, wire114, n_n5181, n_n5184, n_n5183, wire112, n_n5318, n_n5314, n_n5320, wire459, n_n4615, n_n4616, n_n4607, wire396, wire14071, wire14072, n_n3346, n_n4641, n_n4634, n_n4648, n_n4618, n_n4628, wire26, wire118, wire309, wire14078, n_n3281, n_n5050, n_n5060, n_n5055, n_n5054, n_n5059, n_n5048, n_n5028, n_n5036, wire50, n_n5039, wire97, wire13983, wire231, wire356, n_n4571, n_n4578, n_n4570, n_n4849, n_n4853, n_n4847, n_n5096, n_n5099, n_n5085, n_n4314, n_n4389, n_n4369, n_n4381, n_n4340, wire280, n_n5101, n_n5110, n_n5142, n_n5107, n_n5130, n_n5123, n_n5129, n_n5156, n_n4317, n_n4318, n_n4388, n_n4459, n_n4461, n_n4455, n_n4513, n_n4515, n_n4512, n_n4790, n_n4791, n_n4787, n_n4859, n_n4860, n_n4858, n_n4926, n_n4928, n_n4925, n_n4988, n_n4987, n_n5041, n_n5042, n_n5100, n_n4724, n_n4727, n_n4739, wire95, wire244, n_n4864, n_n4868, n_n5018, n_n5022, n_n5017, wire135, wire296, n_n4993, n_n4994, n_n1576, wire134, wire252, n_n5005, n_n5004, n_n5000, wire136, wire393, n_n4907, n_n4913, n_n4922, n_n4934, wire14801, wire14802, wire14803, wire14807, n_n2451, n_n4951, n_n5010, wire14810, wire14814, n_n2462, n_n4886, n_n4865, wire14819, n_n2464, wire31, n_n4453, n_n4420, n_n4407, n_n2470, wire14833, wire14834, wire14848, n_n2455, n_n2467, wire14861, wire14862, wire14870, n_n2454, n_n4391, wire14875, wire14876, n_n2472, n_n4316, n_n4313, wire14881, wire14882, n_n2473, wire234, n_n4372, n_n4373, n_n4371, n_n4431, n_n4433, n_n4430, n_n4494, n_n4491, n_n4834, n_n4835, n_n4832, n_n4909, n_n4911, n_n4903, n_n4979, n_n5049, n_n5179, n_n5239, n_n5240, n_n5238, n_n4514, wire791, n_n4247, n_n4646, n_n4644, n_n4651, n_n4649, wire311, n_n4952, n_n4950, n_n3803, n_n4942, wire59, n_n4945, n_n4946, n_n4949, wire12166, wire16327, n_n2222, n_n5244, n_n5245, wire318, wire16686, n_n4450, n_n4445, n_n4444, n_n4442, n_n4441, wire368, n_n4470, n_n4460, n_n4473, n_n4466, n_n4895, n_n4890, wire260, wire16331, n_n4850, wire277, wire295, wire16334, n_n2228, n_n4881, n_n4878, n_n4880, n_n4869, n_n4877, wire174, wire16342, n_n2178, n_n5321, n_n5323, n_n5324, n_n5322, n_n2274, n_n5307, n_n5326, n_n5325, n_n5332, n_n5329, wire115, wire16291, wire117, wire269, n_n2230, n_n2229, wire16362, wire16363, n_n2179, n_n4776, n_n4774, n_n4786, wire131, wire313, wire16374, wire16375, n_n2162, n_n4755, n_n4759, n_n4760, n_n4758, n_n2238, wire16394, wire16395, wire16399, n_n2182, n_n2242, wire16410, wire16411, wire16415, n_n2183, wire16423, wire16424, n_n2163, n_n4963, n_n4959, n_n4960, n_n4964, n_n2223, wire16449, wire16450, wire16456, n_n2177, wire250, n_n4817, n_n4827, n_n4816, n_n5097, n_n5019, n_n4416, n_n4523, n_n4547, n_n4539, n_n4521, n_n4544, n_n4557, n_n4560, n_n4553, n_n4800, n_n4777, n_n4778, n_n4780, n_n2130, n_n4803, n_n4783, n_n4812, n_n4811, n_n4781, n_n4674, n_n4661, wire16508, wire16509, n_n4361, n_n4363, n_n4359, n_n4438, n_n4439, n_n4437, n_n4825, n_n4828, n_n4824, n_n4879, n_n4937, n_n4938, n_n4936, n_n5037, n_n1570, n_n5043, n_n5045, n_n5302, n_n5294, n_n4894, n_n4916, n_n4930, n_n4947, wire96, n_n5131, n_n5137, n_n5136, n_n5200, n_n5206, n_n5146, n_n5204, n_n5191, n_n5113, n_n5081, n_n5089, n_n5124, wire335, n_n5258, n_n5274, n_n5232, n_n5255, n_n5267, n_n5222, n_n5212, n_n4344, n_n4345, n_n4343, n_n4392, n_n4393, n_n4612, n_n4611, n_n4669, n_n4673, n_n4668, n_n4734, n_n4733, n_n4792, n_n4854, n_n4855, n_n4912, n_n4908, n_n4966, n_n4968, n_n5014, n_n5015, n_n5012, n_n5067, n_n5069, n_n5066, n_n5241, n_n5243, n_n5300, n_n5299, n_n4364, n_n3533, n_n4366, n_n4365, wire11607, n_n1308, n_n4770, n_n4769, n_n4767, n_n4764, n_n4905, wire352, n_n5046, n_n5056, n_n5057, wire166, wire292, n_n4843, n_n4845, n_n4846, n_n4848, n_n4839, n_n4840, n_n4838, n_n3820, n_n4384, n_n4390, n_n4638, n_n4633, n_n5155, n_n5161, n_n4425, n_n4482, n_n4489, n_n4504, n_n4511, n_n4526, n_n4533, n_n4554, n_n4561, n_n4568, n_n4575, n_n4590, n_n4640, n_n4647, n_n4662, n_n4690, n_n4704, n_n4711, n_n4748, n_n4821, n_n4901, n_n4974, n_n5003, n_n5047, n_n5098, n_n5105, n_n5120, n_n5127, n_n5186, n_n5193, n_n5251, n_n5266, n_n5273, n_n4347, n_n4397, n_n4398, n_n4396, n_n4524, n_n4522, wire170, n_n4246, n_n4670, n_n4732, n_n4789, n_n4906, n_n4967, n_n5086, n_n5087, n_n4589, n_n4587, n_n881, n_n4594, n_n4083, n_n4639, n_n4904, n_n4319, n_n4320, n_n4451, n_n4918, n_n4919, n_n4917, n_n4985, n_n4984, n_n5031, n_n5114, n_n5116, n_n5162, n_n4582, n_n4584, n_n4586, wire365, wire14091, wire14092, n_n3348, n_n4876, n_n4870, n_n4871, n_n4872, wire461, wire13850, n_n3326, n_n5327, n_n2643, n_n4577, n_n4576, n_n4569, n_n4574, n_n4581, n_n4572, n_n4573, n_n4579, wire14087, wire14088, wire14101, n_n3282, n_n4538, n_n4525, n_n4531, n_n4551, n_n4552, n_n3871, wire212, n_n4550, n_n4543, wire14107, wire202, wire14115, wire14116, n_n3260, n_n4629, n_n4583, n_n4842, n_n4844, n_n5303, n_n5182, n_n5173, n_n5165, n_n5230, n_n5166, n_n5163, n_n5214, n_n5002, n_n5053, n_n5033, n_n5051, n_n5006, n_n4454, n_n4518, n_n4517, wire664, n_n3152, n_n4725, n_n4726, n_n4861, n_n5103, n_n5104, n_n5102, n_n4395, n_n4357, wire15032, wire15033, n_n2638, wire425, wire15028, wire15029, n_n2560, n_n4426, n_n4409, wire15048, wire15049, n_n2635, wire37, wire15044, n_n2559, n_n4315, n_n4360, n_n4487, n_n4483, n_n4837, n_n4899, n_n4986, n_n5044, n_n5115, n_n5175, n_n5177, n_n5311, n_n4798, n_n4804, n_n4794, n_n4795, n_n4793, n_n4796, n_n4797, n_n4801, n_n4933, n_n4935, wire249, wire289, n_n4497, wire65, wire66, n_n4478, n_n4477, n_n4475, n_n4476, wire70, wire184, wire16576, wire693, wire388, wire16351, wire16352, wire176, wire16355, wire16356, n_n4822, n_n4823, n_n4806, n_n4820, n_n4818, n_n4810, wire186, n_n4415, wire16520, wire16521, n_n2263, wire16527, n_n4326, n_n2446, n_n4336, wire14473, n_n2443, n_n4328, n_n4330, n_n2445, wire171, wire198, wire283, n_n2435, n_n4386, wire12447, wire14460, wire54, n_n4370, n_n4368, wire282, wire423, n_n4503, n_n4502, n_n4500, n_n4546, n_n4555, wire213, n_n4656, n_n4659, n_n5106, n_n4341, n_n5117, n_n5223, n_n5328, n_n5254, n_n5249, n_n5233, n_n5236, n_n5262, n_n5278, wire449, wire16774, wire16775, wire16776, wire16777, n_n2083, n_n4375, n_n4833, n_n4875, n_n4940, n_n4939, n_n4729, n_n4728, wire373, wire374, n_n5132, n_n5128, n_n5016, wire732, n_n4129, n_n5306, n_n5308, n_n3019, n_n5009, n_n5335, n_n4562, n_n4506, n_n4492, n_n4580, n_n4635, wire12047, wire12048, n_n1338, n_n4496, n_n4535, wire12054, n_n1326, n_n4743, wire12067, wire12068, n_n1336, n_n4788, wire12074, wire12075, wire12083, n_n1325, n_n4342, n_n4608, n_n4610, n_n4606, n_n4675, n_n4676, n_n4730, n_n4802, n_n4851, n_n4852, n_n4914, n_n4962, n_n4956, n_n5020, n_n5064, n_n5189, n_n5190, n_n5188, n_n4352, n_n4351, n_n4356, wire67, wire11610, wire11611, n_n1120, n_n4507, n_n4509, n_n4508, wire129, wire308, n_n4622, n_n4621, wire75, n_n3861, n_n5073, n_n5074, n_n5072, n_n4152, n_n4931, wire180, wire382, n_n4978, n_n4980, n_n4897, n_n1985, n_n3815, wire11818, n_n1077, wire264, n_n4349, n_n4348, n_n1002, n_n5172, n_n4419, n_n4605, n_n4655, n_n4683, n_n4689, n_n4697, n_n4703, n_n4712, n_n4763, n_n4915, n_n4989, n_n5011, n_n5061, n_n5070, n_n5076, n_n5135, n_n5157, n_n5201, n_n5207, n_n5237, n_n5252, n_n4353, n_n4456, n_n4671, n_n4747, n_n4772, n_n4773, n_n4771, wire12393, n_n5023, n_n5024, n_n5082, n_n5084, n_n5275, n_n5276, n_n4600, wire45, n_n4775, n_n4204, n_n4065, wire13162, wire13163, wire13166, wire13177, wire13178, wire13181, wire13228, wire13229, wire13233, wire13236, n_n3990, n_n4753, n_n4752, n_n4075, wire13249, wire13250, wire13254, n_n4013, wire47, wire13270, n_n3992, n_n4457, n_n5075, n_n5079, n_n5088, n_n5078, n_n5083, wire123, wire122, wire232, n_n5063, n_n5058, wire160, n_n4891, n_n4836, wire14260, wire14261, n_n3558, wire14267, wire14268, n_n3557, n_n3560, n_n3561, wire14332, n_n3548, n_n4505, n_n5095, n_n5158, n_n5154, n_n3469, n_n5013, n_n5150, n_n5147, wire76, wire196, wire57, wire251, n_n4948, n_n4957, n_n4971, wire342, n_n4471, n_n4490, n_n4479, n_n901, wire14120, n_n3358, wire14126, wire14127, wire14131, n_n3285, n_n4423, n_n4421, wire84, n_n4446, wire470, n_n4630, n_n5065, n_n5287, n_n5281, n_n5268, n_n5261, wire13709, wire13710, n_n4332, n_n4329, n_n4448, n_n4449, n_n4447, n_n5029, n_n4468, n_n3162, n_n4472, n_n4469, n_n4474, wire15423, n_n3001, wire465, n_n4620, n_n5001, n_n2601, n_n2602, wire14904, wire14905, n_n4867, n_n4866, n_n4889, wire12179, n_n2597, n_n4863, n_n2727, wire14927, n_n4965, wire228, n_n2611, wire15011, wire15012, wire15016, wire315, n_n4321, n_n4972, n_n5118, n_n5119, n_n5229, n_n5228, n_n5295, n_n4540, n_n4536, n_n4532, n_n4541, wire416, n_n4681, n_n4679, n_n4677, n_n4678, wire81, wire16404, wire16405, wire414, wire345, wire164, n_n4465, n_n4443, n_n5121, n_n5122, n_n4486, n_n4484, wire199, n_n4893, wire154, wire16784, wire16785, n_n2095, n_n5168, wire16795, wire16796, n_n2091, n_n4973, wire16790, n_n2084, n_n4377, n_n4710, n_n4709, n_n4765, n_n4603, n_n4604, n_n2037, n_n4588, n_n4595, wire16038, n_n1877, wire12309, wire12310, n_n1450, n_n5152, n_n5149, wire195, wire358, wire406, n_n5288, n_n4751, wire12122, wire12123, n_n1333, n_n4435, n_n4626, n_n4627, n_n4625, n_n4660, n_n4719, n_n4954, n_n4955, n_n5133, n_n5138, n_n5139, n_n5309, n_n4387, wire420, n_n4619, wire179, n_n4750, n_n4745, n_n4736, wire293, n_n4722, n_n4721, wire457, n_n5159, n_n5160, wire287, n_n5169, wire33, wire107, wire113, wire254, n_n4658, n_n5108, n_n4510, n_n4424, n_n4498, n_n4591, n_n4663, n_n4698, n_n4705, n_n4805, n_n4841, n_n4944, n_n5068, n_n5187, n_n5199, n_n5260, n_n5272, n_n4405, n_n4406, n_n4462, n_n4501, n_n4684, n_n4222, n_n4741, n_n4740, n_n4819, n_n5077, n_n5221, n_n5220, n_n834, n_n5134, n_n5125, wire336, wire13322, wire13323, wire13325, wire13327, n_n3988, n_n5290, n_n5291, n_n5292, n_n5304, wire13329, wire13347, wire441, wire13365, wire13374, n_n3987, n_n4410, n_n4652, n_n4650, wire14658, wire14659, n_n3681, wire14661, wire14662, wire14667, wire159, n_n5226, n_n5218, wire435, n_n5153, n_n5021, n_n4654, wire140, wire391, n_n4665, wire72, wire418, wire248, n_n4394, wire14168, n_n3363, wire14173, n_n3362, wire14178, wire14179, n_n3287, n_n4279, wire14183, wire363, n_n3370, wire156, wire14163, wire14164, wire14195, n_n3262, n_n4896, n_n4428, wire403, n_n4499, n_n4545, wire471, n_n4376, n_n3176, n_n4585, n_n4873, n_n4932, n_n4592, n_n5052, wire15601, wire15602, n_n2956, n_n5235, n_n5234, n_n5286, n_n5285, n_n1764, n_n3810, n_n2304, n_n5256, n_n5253, n_n1139, n_n4414, wire215, wire16691, wire16692, wire16696, n_n5170, wire168, wire16682, wire16683, n_n2214, wire16753, wire16754, wire16758, n_n5333, n_n4429, n_n4813, n_n4815, wire85, wire16811, wire16812, n_n2096, n_n4715, n_n4714, n_n5225, n_n5224, n_n1530, wire437, n_n5279, n_n5277, n_n4708, n_n4706, wire366, n_n4427, n_n4716, n_n4807, n_n1162, n_n5312, n_n5313, n_n4596, wire256, wire11912, n_n1059, wire11914, wire28, n_n4672, n_n4418, n_n4688, n_n4961, n_n5140, n_n5194, n_n5259, n_n5271, n_n4537, n_n4614, wire13202, wire13203, n_n4058, n_n4016, wire13468, n_n3993, n_n4021, wire13520, n_n3995, wire12471, wire55, wire13553, wire13554, n_n4707, n_n4701, n_n4643, n_n4642, wire14393, n_n3716, wire14398, n_n3650, n_n4556, wire455, wire91, wire430, n_n4609, wire14422, wire14423, n_n3718, wire14419, wire14420, wire14436, n_n4358, n_n4493, n_n5148, n_n3461, wire11769, n_n3329, n_n5126, wire13923, wire13924, n_n3307, wire13796, wire13797, n_n4808, wire13803, wire13804, n_n3330, wire13813, n_n3275, n_n2710, wire13855, wire13856, wire13860, n_n3274, wire13867, wire58, wire13844, n_n3257, wire12778, wire456, n_n4799, wire13746, wire13747, wire13753, n_n4685, n_n4520, n_n5008, n_n4623, wire304, wire14894, wire14898, wire14899, wire433, n_n5242, wire320, n_n5264, n_n5270, wire77, wire334, wire149, n_n5315, wire13557, wire267, wire15195, wire15198, wire218, wire385, wire399, wire125, wire16749, wire44, wire332, n_n5080, wire209, wire90, n_n5090, wire13305, wire13306, wire144, wire239, n_n4411, n_n5219, wire12156, n_n1521, n_n4528, n_n4529, n_n5319, wire328, n_n4542, wire201, n_n4549, n_n4691, n_n3849, n_n4692, wire11862, n_n1093, wire299, n_n1050, n_n5269, n_n5257, wire62, wire92, wire409, wire11923, wire11927, n_n1048, wire63, wire200, wire11929, n_n1017, wire11944, wire11946, wire175, n_n4686, n_n4354, n_n5196, n_n5203, n_n5210, n_n5217, wire13566, wire13567, n_n3996, n_n4929, n_n4766, wire447, n_n1592, n_n4742, n_n4527, n_n4713, wire14347, wire14350, wire14351, n_n4657, wire14363, n_n3711, wire14362, n_n3649, n_n3724, wire14453, wire14454, wire14458, n_n3653, n_n3729, wire14522, n_n3655, n_n5144, n_n5143, n_n2685, wire13929, n_n3308, n_n5007, wire211, wire14065, wire14066, wire14068, n_n4953, wire13772, wire13773, n_n4334, wire158, wire380, n_n4874, wire49, wire87, wire182, n_n5215, wire220, wire384, wire454, n_n4534, n_n2630, wire15065, wire15066, wire15075, n_n2558, wire15079, wire15080, n_n2626, wire15094, wire15095, wire15103, wire82, wire783, wire11564, wire224, n_n5248, n_n4412, n_n5280, n_n5195, n_n5197, n_n5209, n_n5208, n_n2291, wire451, n_n4723, n_n4892, n_n5213, n_n1532, wire288, n_n5247, wire446, wire12349, n_n1435, n_n1103, wire181, wire452, n_n5211, n_n1111, wire11511, wire11512, wire11518, wire79, wire11543, n_n3875, wire11602, wire11605, n_n1040, n_n4322, wire11614, wire11618, n_n1041, n_n4695, n_n4826, n_n5151, wire773, n_n4197, wire330, n_n5071, n_n1167, wire14211, n_n2997, n_n5198, wire14615, n_n3037, wire183, wire453, n_n5246, n_n5176, wire80, wire157, wire15239, n_n2579, wire88, wire15245, n_n2541, wire297, wire394, wire15235, wire14838, wire14839, wire14854, wire14855, wire361, wire378, wire341, wire362, wire203, wire205, wire438, n_n4699, n_n4687, wire340, n_n5250, n_n5205, n_n801, wire12255, wire12256, n_n1454, wire12352, wire12353, n_n1436, n_n5330, n_n5331, wire421, wire225, wire11856, wire253, wire12009, n_n1061, wire12014, wire12015, wire12020, n_n1022, wire104, wire12004, n_n4323, wire128, n_n910, n_n4631, wire12595, wire12596, n_n4761, n_n4680, wire343, wire379, wire15444, wire15445, n_n2996, wire431, n_n2670, n_n4402, wire238, wire276, n_n4702, wire12159, n_n4599, wire364, n_n5283, wire333, n_n4632, wire139, wire11646, wire11647, n_n953, wire99, wire11642, wire787, wire13020, n_n725, wire52, wire150, n_n4645, wire310, n_n4696, n_n4762, n_n1952, wire13512, wire407, wire13209, n_n4056, wire42, n_n814, wire141, wire317, n_n5192, wire106, wire375, n_n4558, wire417, wire12449, wire27, wire12207, wire12208, n_n1472, n_n763, wire286, wire12871, wire12872, n_n667, wire12874, n_n761, wire12876, wire12877, wire12881, n_n635, wire12884, n_n777, n_n3772, wire12894, wire12898, n_n637, n_n4559, n_n5227, n_n4694, n_n4700, n_n4219, wire221, wire13244, wire173, wire13246, wire13156, wire12225, wire390, wire13576, n_n3926, wire13585, wire13586, n_n3924, wire13592, n_n3923, wire13598, wire13599, n_n3928, wire13897, n_n2378, n_n4693, n_n3051, wire15507, wire15426, n_n3003, wire14917, wire14918, n_n4910, wire190, wire12458, wire12459, n_n1501, wire12465, n_n1426, wire12316, n_n1409, wire12332, wire12333, n_n1448, wire12327, wire12328, wire12340, n_n1408, wire347, n_n789, wire12902, n_n680, wire12908, n_n639, wire12930, n_n625, n_n4548, wire13531, n_n4099, wire13529, wire445, wire422, wire442, wire386, wire789, n_n3879, n_n2058, wire324, wire305, wire291, wire11507, wire12682, wire12683, n_n554, wire279, wire13445, wire13446, wire13452, wire401, wire14316, wire14317, wire434, wire15511, wire15512, n_n3009, wire11520, n_n3889, wire16388, wire16389, n_n1677, wire12493, wire12234, n_n1467, wire12231, wire11866, wire11867, n_n1091, wire13338, wire124, wire12363, wire12364, wire12368, wire12369, n_n1402, wire12371, wire12372, wire204, wire11666, wire11667, n_n956, n_n951, wire11675, wire11676, wire11690, n_n948, n_n949, wire11734, wire11735, wire13342, wire600, n_n1478, n_n1476, wire12416, n_n5289, wire255, n_n1727, wire15829, wire15830, n_n1712, wire15908, wire15909, n_n1730, wire15914, wire15915, n_n1729, n_n1725, n_n1724, wire15930, wire15931, n_n1711, n_n5282, n_n5298, wire13629, wire13630, wire13635, wire13636, wire261, n_n3694, n_n2761, wire15750, wire466, wire15605, wire15606, n_n2953, wire15609, wire15610, n_n2955, wire15616, wire15617, n_n2915, wire265, wire15633, wire15634, wire15642, n_n2902, wire15405, wire15406, wire15069, n_n1840, wire15950, wire15951, wire15957, n_n1801, wire15961, wire15962, n_n1837, wire15968, n_n1800, wire15977, n_n1842, wire15920, wire12783, wire12784, n_n707, n_n691, wire12966, wire12967, n_n632, n_n700, wire12762, n_n646, wire12753, n_n627, wire683, n_n856, wire12790, wire12791, wire12796, n_n648, wire12814, n_n628, wire12865, wire12866, n_n1760, wire15333, wire15334, wire53, wire16159, n_n1852, wire16164, wire16165, wire16168, n_n1805, wire16158, wire444, wire12403, wire12969, wire12970, n_n662, wire12971, wire12975, n_n661, wire13001, wire14470, wire14471, n_n3736, wire15348, wire15349, wire15008, wire13055, wire16188, wire16189, n_n1862, wire16193, wire16194, wire16198, n_n1808, wire16217, n_n1856, wire16213, wire16214, wire16224, wire15822, wire15823, wire15851, wire15852, n_n1722, wire15858, wire15859, n_n1721, wire13028, n_n722, wire13034, wire13035, wire13039, n_n653, wire13016, wire13017, wire13046, n_n630, wire14544, n_n3664, wire15521, n_n3012, wire15517, wire15769, wire15770, n_n2985, wire15774, wire15775, wire15778, n_n2925, n_n2832, n_n2834, wire15367, wire15368, wire15389, wire15390, wire16099, wire16094, wire16105, wire16233, wire12408, wire12409, wire13073, wire13074, n_n732, wire13070, n_n656, wire13066, n_n631, n_n715, wire13106, wire13107, wire13111, n_n651, wire13124, n_n629, wire14322, wire14323, wire15653, n_n2939, wire15354, wire15355, wire15360, wire15361, wire11873, wire11874, n_n1032, wire11718, wire11719, wire12756, wire12757, wire14752, wire14754, n_n3689, wire14448, wire11725, wire11726, wire13100, wire13101, wire14618, wire14619, n_n3670, wire15663, n_n2937, wire15451, wire15452, wire15870, wire15871, n_n1718, wire15875, n_n1717, wire11680, wire11681, wire16300, wire16305, wire15995, wire14438, wire16034, n_n1879, wire16040, wire16041, wire16048, n_n1872, wire16059, wire11852, wire14517, n_n3699, wire14701, wire14702, n_n3701, wire14708, wire14709, n_n3645, wire16052, wire16053, wire16266, wire16267, n_n1828, wire16272, wire14723, wire14624, wire14625, wire14629, wire14760, wire14761, wire14764, wire15766, wire15767, wire15786, wire266, wire606, wire617, wire636, wire656, wire669, wire671, wire675, wire677, wire679, wire686, wire695, wire706, wire724, wire735, wire743, wire745, wire755, wire761, wire765, wire767, wire771, wire772, wire775, wire11482, wire11483, wire11488, wire11489, wire11491, wire11492, wire11495, wire11496, wire11497, wire11498, wire11505, wire11513, wire11515, wire11516, wire11521, wire11522, wire11523, wire11524, wire11527, wire11529, wire11532, wire11534, wire11535, wire11536, wire11539, wire11547, wire11548, wire11549, wire11553, wire11554, wire11555, wire11558, wire11559, wire11560, wire11562, wire11563, wire11566, wire11567, wire11568, wire11570, wire11571, wire11574, wire11575, wire11578, wire11581, wire11582, wire11583, wire11584, wire11585, wire11586, wire11587, wire11588, wire11589, wire11591, wire11592, wire11593, wire11597, wire11598, wire11599, wire11613, wire11620, wire11625, wire11626, wire11628, wire11630, wire11631, wire11633, wire11634, wire11638, wire11653, wire11654, wire11658, wire11660, wire11661, wire11671, wire11677, wire11687, wire11688, wire11693, wire11694, wire11698, wire11699, wire11703, wire11705, wire11706, wire11707, wire11710, wire11712, wire11713, wire11715, wire11731, wire11732, wire11738, wire11739, wire11743, wire11748, wire11751, wire11752, wire11753, wire11754, wire11756, wire11757, wire11759, wire11761, wire11762, wire11765, wire11766, wire11767, wire11768, wire11772, wire11773, wire11774, wire11776, wire11777, wire11778, wire11781, wire11782, wire11783, wire11785, wire11786, wire11788, wire11790, wire11791, wire11795, wire11797, wire11801, wire11802, wire11803, wire11804, wire11805, wire11807, wire11808, wire11809, wire11810, wire11811, wire11812, wire11814, wire11816, wire11824, wire11825, wire11826, wire11829, wire11834, wire11836, wire11837, wire11839, wire11841, wire11842, wire11846, wire11847, wire11848, wire11855, wire11859, wire11870, wire11877, wire11880, wire11881, wire11886, wire11888, wire11889, wire11891, wire11893, wire11899, wire11900, wire11902, wire11906, wire11907, wire11909, wire11916, wire11917, wire11924, wire11928, wire11939, wire11947, wire11951, wire11952, wire11955, wire11959, wire11964, wire11967, wire11968, wire11970, wire11971, wire11972, wire11973, wire11978, wire11981, wire11982, wire11986, wire11987, wire11992, wire11993, wire11994, wire11995, wire11996, wire11997, wire11999, wire12007, wire12018, wire12023, wire12024, wire12027, wire12033, wire12058, wire12060, wire12061, wire12080, wire12081, wire12089, wire12090, wire12091, wire12092, wire12093, wire12096, wire12097, wire12099, wire12101, wire12102, wire12106, wire12108, wire12109, wire12111, wire12113, wire12114, wire12115, wire12117, wire12118, wire12120, wire12126, wire12128, wire12129, wire12131, wire12134, wire12136, wire12137, wire12141, wire12142, wire12146, wire12147, wire12149, wire12152, wire12162, wire12164, wire12165, wire12167, wire12168, wire12169, wire12170, wire12171, wire12172, wire12175, wire12176, wire12177, wire12181, wire12182, wire12183, wire12186, wire12187, wire12188, wire12191, wire12192, wire12196, wire12202, wire12204, wire12205, wire12210, wire12213, wire12214, wire12217, wire12218, wire12219, wire12220, wire12226, wire12232, wire12239, wire12243, wire12245, wire12253, wire12262, wire12266, wire12268, wire12269, wire12271, wire12272, wire12276, wire12277, wire12278, wire12282, wire12283, wire12285, wire12288, wire12290, wire12292, wire12293, wire12296, wire12297, wire12300, wire12301, wire12304, wire12306, wire12317, wire12318, wire12319, wire12323, wire12326, wire12335, wire12337, wire12342, wire12345, wire12355, wire12356, wire12358, wire12359, wire12361, wire12366, wire12376, wire12380, wire12382, wire12384, wire12386, wire12389, wire12391, wire12392, wire12395, wire12398, wire12399, wire12400, wire12401, wire12413, wire12414, wire12420, wire12421, wire12422, wire12425, wire12426, wire12428, wire12435, wire12436, wire12439, wire12442, wire12445, wire12446, wire12448, wire12451, wire12453, wire12456, wire12461, wire12467, wire12472, wire12475, wire12476, wire12478, wire12479, wire12480, wire12481, wire12485, wire12486, wire12488, wire12490, wire12497, wire12498, wire12499, wire12500, wire12501, wire12502, wire12503, wire12507, wire12508, wire12510, wire12514, wire12518, wire12519, wire12520, wire12521, wire12525, wire12530, wire12531, wire12534, wire12535, wire12539, wire12540, wire12541, wire12543, wire12544, wire12545, wire12546, wire12547, wire12551, wire12552, wire12554, wire12555, wire12556, wire12557, wire12559, wire12560, wire12561, wire12564, wire12566, wire12568, wire12569, wire12570, wire12573, wire12574, wire12577, wire12578, wire12579, wire12582, wire12602, wire12607, wire12608, wire12613, wire12614, wire12615, wire12620, wire12621, wire12626, wire12627, wire12629, wire12630, wire12634, wire12635, wire12638, wire12640, wire12641, wire12642, wire12643, wire12648, wire12649, wire12650, wire12651, wire12653, wire12656, wire12657, wire12658, wire12659, wire12663, wire12664, wire12669, wire12670, wire12672, wire12673, wire12675, wire12678, wire12679, wire12688, wire12689, wire12691, wire12693, wire12694, wire12710, wire12722, wire12724, wire12729, wire12730, wire12732, wire12735, wire12736, wire12740, wire12742, wire12743, wire12744, wire12745, wire12747, wire12748, wire12749, wire12759, wire12760, wire12766, wire12770, wire12771, wire12774, wire12787, wire12788, wire12792, wire12794, wire12799, wire12800, wire12801, wire12802, wire12804, wire12805, wire12810, wire12811, wire12815, wire12819, wire12820, wire12822, wire12826, wire12831, wire12832, wire12833, wire12834, wire12835, wire12838, wire12839, wire12841, wire12843, wire12844, wire12845, wire12848, wire12849, wire12852, wire12853, wire12854, wire12857, wire12858, wire12859, wire12862, wire12875, wire12883, wire12888, wire12889, wire12892, wire12893, wire12904, wire12909, wire12914, wire12917, wire12921, wire12922, wire12924, wire12925, wire12926, wire12931, wire12934, wire12935, wire12936, wire12939, wire12940, wire12941, wire12943, wire12946, wire12949, wire12952, wire12953, wire12954, wire12958, wire12960, wire12961, wire12963, wire12972, wire12976, wire12978, wire12979, wire12981, wire12984, wire12985, wire12986, wire12988, wire12989, wire12991, wire12992, wire12996, wire12998, wire13003, wire13005, wire13006, wire13008, wire13013, wire13015, wire13022, wire13025, wire13026, wire13027, wire13036, wire13044, wire13048, wire13049, wire13050, wire13053, wire13054, wire13057, wire13059, wire13060, wire13062, wire13063, wire13067, wire13078, wire13085, wire13087, wire13090, wire13091, wire13093, wire13095, wire13096, wire13104, wire13105, wire13108, wire13113, wire13114, wire13117, wire13118, wire13119, wire13120, wire13126, wire13127, wire13128, wire13132, wire13140, wire13141, wire13144, wire13146, wire13149, wire13151, wire13153, wire13154, wire13171, wire13172, wire13174, wire13182, wire13183, wire13185, wire13187, wire13193, wire13194, wire13198, wire13199, wire13213, wire13215, wire13216, wire13217, wire13218, wire13222, wire13223, wire13224, wire13234, wire13237, wire13239, wire13240, wire13248, wire13251, wire13256, wire13259, wire13260, wire13261, wire13263, wire13264, wire13265, wire13266, wire13268, wire13272, wire13274, wire13277, wire13283, wire13284, wire13285, wire13287, wire13288, wire13291, wire13292, wire13293, wire13294, wire13296, wire13297, wire13298, wire13301, wire13303, wire13304, wire13308, wire13310, wire13311, wire13313, wire13314, wire13317, wire13318, wire13320, wire13334, wire13350, wire13351, wire13352, wire13354, wire13355, wire13359, wire13360, wire13361, wire13368, wire13370, wire13372, wire13378, wire13380, wire13381, wire13384, wire13385, wire13390, wire13391, wire13392, wire13393, wire13394, wire13397, wire13398, wire13399, wire13400, wire13401, wire13404, wire13405, wire13406, wire13408, wire13409, wire13410, wire13411, wire13413, wire13414, wire13415, wire13417, wire13422, wire13424, wire13425, wire13428, wire13429, wire13430, wire13431, wire13432, wire13436, wire13437, wire13438, wire13439, wire13443, wire13448, wire13450, wire13454, wire13455, wire13457, wire13458, wire13459, wire13461, wire13462, wire13463, wire13465, wire13470, wire13471, wire13473, wire13474, wire13475, wire13479, wire13481, wire13487, wire13488, wire13494, wire13495, wire13497, wire13501, wire13502, wire13503, wire13504, wire13505, wire13506, wire13508, wire13509, wire13510, wire13513, wire13515, wire13516, wire13521, wire13522, wire13523, wire13524, wire13525, wire13526, wire13534, wire13535, wire13538, wire13541, wire13542, wire13543, wire13546, wire13550, wire13552, wire13559, wire13560, wire13561, wire13562, wire13577, wire13601, wire13606, wire13607, wire13611, wire13612, wire13616, wire13617, wire13638, wire13648, wire13650, wire13651, wire13656, wire13657, wire13660, wire13662, wire13663, wire13666, wire13670, wire13673, wire13681, wire13683, wire13689, wire13690, wire13694, wire13696, wire13697, wire13698, wire13703, wire13704, wire13713, wire13717, wire13719, wire13720, wire13725, wire13726, wire13735, wire13736, wire13741, wire13742, wire13755, wire13756, wire13765, wire13776, wire13777, wire13779, wire13788, wire13789, wire13790, wire13791, wire13792, wire13798, wire13800, wire13807, wire13810, wire13815, wire13816, wire13823, wire13824, wire13827, wire13833, wire13834, wire13836, wire13837, wire13840, wire13841, wire13854, wire13857, wire13865, wire13866, wire13870, wire13872, wire13873, wire13874, wire13877, wire13880, wire13881, wire13883, wire13884, wire13885, wire13887, wire13888, wire13891, wire13892, wire13893, wire13895, wire13896, wire13900, wire13902, wire13903, wire13905, wire13906, wire13910, wire13911, wire13913, wire13914, wire13915, wire13918, wire13919, wire13920, wire13931, wire13932, wire13934, wire13935, wire13938, wire13940, wire13942, wire13943, wire13944, wire13947, wire13948, wire13952, wire13955, wire13957, wire13960, wire13961, wire13962, wire13963, wire13964, wire13966, wire13967, wire13968, wire13969, wire13971, wire13972, wire13975, wire13977, wire13978, wire13979, wire13981, wire13982, wire13985, wire13989, wire13990, wire13991, wire13992, wire13995, wire13996, wire13997, wire13999, wire14000, wire14001, wire14003, wire14006, wire14007, wire14009, wire14010, wire14011, wire14012, wire14015, wire14016, wire14018, wire14021, wire14023, wire14025, wire14027, wire14028, wire14029, wire14031, wire14033, wire14034, wire14036, wire14037, wire14040, wire14042, wire14043, wire14045, wire14046, wire14047, wire14049, wire14050, wire14055, wire14056, wire14058, wire14061, wire14062, wire14079, wire14080, wire14094, wire14097, wire14099, wire14103, wire14105, wire14106, wire14111, wire14112, wire14128, wire14133, wire14134, wire14138, wire14139, wire14141, wire14142, wire14143, wire14144, wire14148, wire14149, wire14150, wire14153, wire14154, wire14155, wire14157, wire14158, wire14159, wire14160, wire14171, wire14177, wire14192, wire14198, wire14199, wire14200, wire14202, wire14203, wire14205, wire14208, wire14213, wire14214, wire14218, wire14219, wire14226, wire14227, wire14232, wire14233, wire14238, wire14239, wire14240, wire14241, wire14245, wire14246, wire14252, wire14253, wire14254, wire14256, wire14272, wire14273, wire14275, wire14277, wire14278, wire14280, wire14281, wire14283, wire14284, wire14285, wire14290, wire14291, wire14293, wire14295, wire14296, wire14301, wire14302, wire14307, wire14308, wire14311, wire14320, wire14329, wire14330, wire14334, wire14338, wire14340, wire14343, wire14344, wire14349, wire14355, wire14356, wire14365, wire14367, wire14373, wire14375, wire14376, wire14377, wire14378, wire14380, wire14381, wire14385, wire14387, wire14396, wire14401, wire14403, wire14404, wire14408, wire14409, wire14410, wire14413, wire14414, wire14415, wire14416, wire14426, wire14428, wire14429, wire14430, wire14432, wire14434, wire14439, wire14440, wire14441, wire14442, wire14443, wire14444, wire14445, wire14446, wire14452, wire14455, wire14461, wire14464, wire14466, wire14467, wire14468, wire14476, wire14479, wire14480, wire14484, wire14485, wire14486, wire14489, wire14490, wire14492, wire14493, wire14495, wire14496, wire14498, wire14499, wire14500, wire14503, wire14505, wire14507, wire14508, wire14510, wire14511, wire14519, wire14520, wire14523, wire14524, wire14526, wire14533, wire14534, wire14536, wire14537, wire14542, wire14550, wire14551, wire14552, wire14554, wire14555, wire14557, wire14558, wire14560, wire14561, wire14563, wire14564, wire14566, wire14567, wire14570, wire14572, wire14573, wire14577, wire14578, wire14579, wire14580, wire14582, wire14583, wire14587, wire14588, wire14591, wire14592, wire14594, wire14595, wire14598, wire14599, wire14601, wire14603, wire14605, wire14606, wire14609, wire14610, wire14621, wire14622, wire14623, wire14631, wire14635, wire14637, wire14641, wire14644, wire14645, wire14646, wire14648, wire14649, wire14652, wire14656, wire14665, wire14669, wire14671, wire14672, wire14673, wire14674, wire14675, wire14678, wire14680, wire14681, wire14683, wire14690, wire14691, wire14692, wire14695, wire14706, wire14714, wire14715, wire14718, wire14719, wire14724, wire14726, wire14730, wire14735, wire14738, wire14739, wire14740, wire14742, wire14743, wire14745, wire14747, wire14748, wire14756, wire14759, wire14762, wire14766, wire14768, wire14770, wire14774, wire14775, wire14782, wire14784, wire14785, wire14790, wire14791, wire14795, wire14796, wire14797, wire14808, wire14816, wire14817, wire14825, wire14826, wire14829, wire14830, wire14831, wire14836, wire14843, wire14845, wire14846, wire14859, wire14867, wire14868, wire14873, wire14886, wire14887, wire14890, wire14892, wire14896, wire14903, wire14909, wire14910, wire14911, wire14914, wire14915, wire14920, wire14924, wire14931, wire14933, wire14937, wire14938, wire14939, wire14940, wire14942, wire14943, wire14944, wire14946, wire14948, wire14949, wire14954, wire14955, wire14956, wire14957, wire14960, wire14961, wire14962, wire14964, wire14965, wire14967, wire14969, wire14970, wire14971, wire14974, wire14975, wire14978, wire14979, wire14980, wire14982, wire14983, wire14985, wire14986, wire14987, wire14988, wire14990, wire14991, wire14992, wire14993, wire14995, wire14996, wire14999, wire15000, wire15001, wire15002, wire15007, wire15020, wire15021, wire15024, wire15035, wire15038, wire15042, wire15043, wire15046, wire15052, wire15057, wire15058, wire15059, wire15061, wire15062, wire15063, wire15071, wire15077, wire15082, wire15083, wire15084, wire15085, wire15089, wire15090, wire15091, wire15097, wire15099, wire15101, wire15108, wire15109, wire15111, wire15112, wire15113, wire15115, wire15117, wire15120, wire15121, wire15122, wire15123, wire15125, wire15126, wire15127, wire15130, wire15131, wire15132, wire15133, wire15135, wire15136, wire15137, wire15140, wire15141, wire15142, wire15143, wire15144, wire15145, wire15149, wire15153, wire15154, wire15155, wire15159, wire15160, wire15162, wire15163, wire15165, wire15166, wire15174, wire15175, wire15178, wire15179, wire15180, wire15184, wire15185, wire15186, wire15188, wire15189, wire15192, wire15200, wire15203, wire15208, wire15211, wire15212, wire15216, wire15217, wire15218, wire15221, wire15222, wire15223, wire15224, wire15226, wire15227, wire15230, wire15231, wire15241, wire15243, wire15247, wire15252, wire15254, wire15255, wire15257, wire15258, wire15261, wire15263, wire15266, wire15269, wire15270, wire15273, wire15274, wire15275, wire15278, wire15279, wire15280, wire15284, wire15285, wire15288, wire15289, wire15290, wire15292, wire15294, wire15296, wire15304, wire15310, wire15312, wire15315, wire15316, wire15326, wire15340, wire15341, wire15375, wire15376, wire15382, wire15383, wire15385, wire15396, wire15397, wire15416, wire15421, wire15428, wire15431, wire15432, wire15434, wire15435, wire15448, wire15456, wire15459, wire15460, wire15468, wire15469, wire15472, wire15474, wire15475, wire15478, wire15479, wire15481, wire15482, wire15483, wire15485, wire15488, wire15489, wire15490, wire15493, wire15495, wire15498, wire15499, wire15509, wire15525, wire15526, wire15529, wire15532, wire15533, wire15534, wire15536, wire15537, wire15538, wire15539, wire15542, wire15546, wire15551, wire15554, wire15555, wire15557, wire15559, wire15560, wire15562, wire15565, wire15569, wire15570, wire15573, wire15574, wire15575, wire15576, wire15579, wire15582, wire15583, wire15586, wire15587, wire15589, wire15591, wire15593, wire15595, wire15596, wire15597, wire15598, wire15612, wire15614, wire15620, wire15621, wire15623, wire15624, wire15626, wire15627, wire15628, wire15629, wire15639, wire15647, wire15648, wire15649, wire15651, wire15658, wire15659, wire15660, wire15666, wire15667, wire15671, wire15672, wire15675, wire15677, wire15678, wire15680, wire15681, wire15683, wire15684, wire15685, wire15686, wire15688, wire15689, wire15693, wire15695, wire15696, wire15697, wire15698, wire15700, wire15701, wire15702, wire15704, wire15705, wire15707, wire15709, wire15710, wire15712, wire15715, wire15718, wire15719, wire15721, wire15723, wire15724, wire15725, wire15729, wire15733, wire15734, wire15738, wire15739, wire15741, wire15747, wire15748, wire15754, wire15756, wire15757, wire15758, wire15760, wire15761, wire15763, wire15773, wire15776, wire15781, wire15784, wire15790, wire15791, wire15792, wire15794, wire15795, wire15798, wire15799, wire15800, wire15802, wire15805, wire15807, wire15811, wire15813, wire15819, wire15834, wire15836, wire15837, wire15841, wire15842, wire15843, wire15844, wire15845, wire15848, wire15864, wire15865, wire15873, wire15876, wire15880, wire15885, wire15886, wire15887, wire15892, wire15894, wire15895, wire15897, wire15898, wire15899, wire15901, wire15902, wire15903, wire15922, wire15927, wire15937, wire15938, wire15941, wire15943, wire15947, wire15952, wire15954, wire15964, wire15970, wire15972, wire15975, wire15980, wire15982, wire15983, wire15985, wire15987, wire15989, wire15991, wire15993, wire15999, wire16001, wire16002, wire16003, wire16004, wire16007, wire16008, wire16009, wire16011, wire16012, wire16014, wire16015, wire16016, wire16018, wire16019, wire16020, wire16022, wire16023, wire16031, wire16032, wire16045, wire16046, wire16056, wire16057, wire16064, wire16069, wire16075, wire16077, wire16078, wire16081, wire16082, wire16083, wire16088, wire16091, wire16093, wire16102, wire16103, wire16109, wire16110, wire16112, wire16119, wire16120, wire16121, wire16124, wire16125, wire16130, wire16131, wire16132, wire16134, wire16135, wire16139, wire16140, wire16141, wire16144, wire16145, wire16146, wire16148, wire16149, wire16152, wire16153, wire16155, wire16166, wire16171, wire16174, wire16175, wire16179, wire16182, wire16184, wire16185, wire16186, wire16192, wire16195, wire16201, wire16203, wire16204, wire16206, wire16207, wire16211, wire16215, wire16222, wire16229, wire16236, wire16238, wire16245, wire16246, wire16248, wire16249, wire16251, wire16253, wire16254, wire16256, wire16257, wire16258, wire16259, wire16270, wire16278, wire16279, wire16282, wire16286, wire16288, wire16293, wire16294, wire16297, wire16306, wire16308, wire16309, wire16310, wire16312, wire16313, wire16320, wire16339, wire16340, wire16345, wire16346, wire16347, wire16349, wire16350, wire16360, wire16366, wire16367, wire16368, wire16373, wire16378, wire16379, wire16382, wire16383, wire16385, wire16386, wire16396, wire16408, wire16409, wire16412, wire16420, wire16421, wire16427, wire16430, wire16431, wire16435, wire16436, wire16438, wire16442, wire16443, wire16447, wire16448, wire16453, wire16454, wire16461, wire16462, wire16463, wire16465, wire16468, wire16470, wire16479, wire16480, wire16482, wire16483, wire16487, wire16488, wire16490, wire16498, wire16500, wire16506, wire16514, wire16518, wire16531, wire16537, wire16538, wire16539, wire16544, wire16548, wire16549, wire16551, wire16552, wire16556, wire16560, wire16562, wire16563, wire16566, wire16567, wire16568, wire16570, wire16571, wire16572, wire16574, wire16578, wire16580, wire16581, wire16585, wire16586, wire16587, wire16590, wire16591, wire16593, wire16594, wire16596, wire16598, wire16599, wire16601, wire16602, wire16603, wire16605, wire16606, wire16609, wire16611, wire16612, wire16617, wire16618, wire16621, wire16623, wire16627, wire16628, wire16629, wire16631, wire16632, wire16633, wire16635, wire16636, wire16638, wire16641, wire16642, wire16644, wire16645, wire16646, wire16656, wire16657, wire16658, wire16662, wire16663, wire16666, wire16670, wire16673, wire16674, wire16676, wire16677, wire16678, wire16679, wire16690, wire16693, wire16698, wire16699, wire16702, wire16704, wire16709, wire16710, wire16711, wire16715, wire16716, wire16717, wire16718, wire16719, wire16721, wire16723, wire16724, wire16728, wire16730, wire16731, wire16739, wire16740, wire16742, wire16755, wire16760, wire16761, wire16769, wire16770, wire16773, wire16788, wire16798, wire16799, wire16804, wire16818, wire16819, wire16820, wire16823, wire16825, wire16827, wire16829, _38, _64, _72, _90, _120, _144, _172, _198, _204, _206, _220, _226, _230, _298, _348, _356, _362, _364, _388, _462, _514, _560, _564, _600, _660, _664, _670, _672, _690, _708, _778, _904, _930, _932, _1018, _1050, _1120, _1152, _1160, _1176, _1190, _1204, _1230, _1240, _1244, _1366, _1394, _1428, _1490, _1514, _1694, _22059, _22066, _22147, _22149, _22150, _22151, _22193, _22194, _22212, _22253, _22279, _22321, _22359, _22360, _22415, _22416, _22433, _22464, _22478, _22494, _22495, _22502, _22511, _22549, _22550, _22551, _22552, _22574, _22575, _22614, _22691, _22692, _22732, _22733, _22749, _22752, _22800, _22801, _22829, _22846, _22891, _22972, _22973, _22987, _23016, _23017, _23150, _23316, _23327, _23360, _23446, _23478, _23479, _23490, _23507, _23508, _23538, _23540, _23541, _23543, _23548, _23567, _23568, _23569, _23648, _23670, _23708, _23747, _23753, _23780, _23821, _23822, _23853, _23965, _23986, _23987, _24115, _24138, _24139, _24226, _24227, _24250, _24258, _24270, _24285, _24286, _24317, _24320, _24373, _24405, _24444, _24445, _24448, _24456, _24460, _24477, _24485, _24486, _24493, _24526, _24527, _24555, _24594, _24595, _24602, _24620, _24621, _24749, _24750, _24759, _24803, _24805, _24806, _24831, _24874, _24885, _24886, _24893, _24946, _24947, _24948, _24968, _24971, _24973, _24974, _24978, _24983, _25017, _25018, _25047, _25048, _25076, _25084, _25085, _25094, _25187, _25250, _25251, _25252, _25280, _25314, _25315, _25322, _25336, _25337, _25342, _25369, _25381, _25382, _25401, _25431, _25432, _25436, _25438, _25451, _25538, _25555, _25558, _25595, _25596, _25597, _25598, _25613, _25616, _25630, _25638, _25639, _25642, _25663, _25671, _25724, _25725, _25791, _25808, _25813, _25815, _25818, _25825, _25826, _25832, _25847, _25860, _25862, _25892, _25931, _25940, _25945, _25967, _25970, _25975, _25978, _25980, _26007, _26036, _26043, _26064, _26108, _26110, _26122, _26133, _26177, _26195, _26246, _26247, _26248, _26253, _26270, _26291, _26294, _26299, _26304, _26306, _26307, _26324, _26339, _26353, _26354, _26367, _26379, _26416, _26417, _26451, _26476, _26486, _26498, _26499, _26500, _26515, _26519, _26573, _26577, _26585, _26606, _26631, _26646, _26648, _26776, _26794, _26795, _26796, _26834, _26840, _26875, _26878, _26879, _26880, _26883, _26907, _26926, _26929, _26931, _26964, _27049, _27085, _27086, _27110, _27137, _27138, _27142, _27156, _27192, _27197, _27206, _27223, _27224, _27225, _27243, _27245, _27260, _27356, _27364, _27368, _27369, _27388, _27389, _27390, _27424, _27425, _27427, _27452, _27453, _27469, _27470, _27472, _27475, _27476, _27478, _27489, _27498, _27515, _27519, _27547, _27548, _27572, _27574, _27575, _27581, _27582, _27584, _27589, _27591, _27623, _27671, _27702, _27703, _27731, _27741, _27832, _27833, _27835, _27854, _27859, _27861, _27868, _27885, _27896, _27897, _27906, _27910, _27917, _27951, _27952, _27996, _28000, _28058, _28071, _28106, _28114, _28116, _28124, _28137, _28144, _28151, _28172, _28175, _28185, _28238, _28239, _28262, _28268, _28280, _28289, _28301, _28305, _28312, _28313, _28320, _28341, _28352, _28355, _28357, _28359, _28361, _28362, _28370, _28382, _28406, _28412, _28413, _28416, _28422, _28424, _28427, _28441, _28496, _28538, _28546, _28573, _28574, _28575, _28577, _28581, _28589, _28605, _28607, _28618, _28636, _28637, _28642, _28665, _28666, _28668, _28669, _28677, _28704, _28709, _28710, _28731, _28734, _28735, _28741, _28749, _28750, _28753, _28757, _28767, _28771, _28786, _28787, _28790, _28794, _28812, _28817, _28838, _28839, _28844, _28847, _28857, _28879, _28882, _28884, _28885, _28888, _28895, _28900, _28912, _28923, _28927, _28931, _28934, _28935, _28949, _28951, _28952, _29002, _29003, _29004, _29006, _29007, _29028, _29029, _29041, _29050, _29051, _29082, _29086, _29091, _29098, _29100, _29196, _29216, _29219, _29241, _29242, _29247, _29258, _29270, _29306, _29324, _29335;

assign o_1_ = ( n_n1005 ) | ( n_n1004 ) | ( wire12040 ) | ( wire12041 ) ;
 assign o_2_ = ( wire12585 ) | ( wire12586 ) | ( wire12588 ) | ( wire12589 ) ;
 assign o_0_ = ( n_n621 ) | ( n_n620 ) | ( wire13136 ) | ( wire13147 ) ;
 assign o_9_ = ( n_n3986 ) | ( wire13573 ) | ( _25980 ) ;
 assign o_7_ = ( n_n3253 ) | ( wire14216 ) | ( _26631 ) ;
 assign o_8_ = ( n_n3622 ) | ( wire14777 ) | ( wire14778 ) | ( wire14779 ) ;
 assign o_5_ = ( n_n2525 ) | ( n_n2523 ) | ( wire15299 ) | ( wire15300 ) ;
 assign o_6_ = ( n_n2898 ) | ( wire15816 ) | ( wire15817 ) ;
 assign o_3_ = ( n_n1784 ) | ( wire16323 ) | ( wire16324 ) ;
 assign o_4_ = ( wire16830 ) | ( wire16831 ) | ( _28951 ) | ( _28952 ) ;
 assign n_n1005 = ( n_n1012 ) | ( wire11893 ) | ( _22415 ) | ( _22416 ) ;
 assign n_n1004 = ( n_n1007 ) | ( n_n1009 ) | ( wire12036 ) | ( wire12037 ) ;
 assign wire12040 = ( n_n1014 ) | ( wire11581 ) | ( wire11582 ) ;
 assign wire12041 = ( n_n4309 ) | ( n_n1040 ) | ( n_n1041 ) | ( wire11634 ) ;
 assign wire12585 = ( n_n1426 ) | ( wire12582 ) | ( _23540 ) | ( _23541 ) ;
 assign wire12586 = ( wire12518 ) | ( wire12568 ) | ( _23747 ) ;
 assign wire12588 = ( n_n1398 ) | ( n_n1326 ) | ( n_n1325 ) | ( wire12152 ) ;
 assign wire12589 = ( n_n1396 ) | ( n_n1397 ) | ( wire12391 ) | ( wire12392 ) ;
 assign n_n621 = ( n_n627 ) | ( n_n628 ) | ( wire12865 ) | ( wire12866 ) ;
 assign n_n620 = ( n_n635 ) | ( n_n637 ) | ( n_n625 ) | ( wire13001 ) ;
 assign wire13136 = ( n_n630 ) | ( n_n631 ) | ( n_n629 ) ;
 assign wire13147 = ( wire12693 ) | ( wire12694 ) | ( wire13146 ) ;
 assign n_n3986 = ( n_n3993 ) | ( n_n3995 ) | ( wire13553 ) | ( wire13554 ) ;
 assign wire13572 = ( wire13424 ) | ( _25596 ) | ( _25597 ) | ( _25598 ) ;
 assign wire13573 = ( n_n3990 ) | ( n_n3992 ) | ( n_n3988 ) | ( n_n3987 ) ;
 assign n_n3253 = ( n_n3260 ) | ( n_n3262 ) | ( wire14211 ) ;
 assign wire14216 = ( n_n3257 ) | ( wire13919 ) | ( wire13920 ) | ( wire14214 ) ;
 assign wire14222 = ( n_n3187 ) | ( n_n3192 ) | ( n_n3191 ) | ( wire14219 ) ;
 assign n_n3622 = ( n_n3629 ) | ( wire14513 ) | ( wire14514 ) | ( wire14540 ) ;
 assign wire14777 = ( n_n3639 ) | ( wire14684 ) | ( _26875 ) | ( _26931 ) ;
 assign wire14778 = ( n_n3626 ) | ( wire14277 ) | ( wire14278 ) | ( wire14343 ) ;
 assign wire14779 = ( n_n3624 ) | ( wire14591 ) | ( wire14592 ) | ( wire14775 ) ;
 assign n_n2525 = ( n_n2533 ) | ( wire15150 ) | ( wire15151 ) | ( wire15169 ) ;
 assign n_n2523 = ( n_n2528 ) | ( wire15296 ) | ( _27547 ) | ( _27548 ) ;
 assign wire15299 = ( n_n2530 ) | ( wire14979 ) | ( wire14980 ) | ( wire14982 ) ;
 assign wire15300 = ( n_n2531 ) | ( wire14829 ) | ( wire14830 ) | ( wire14892 ) ;
 assign n_n2898 = ( n_n2905 ) | ( wire15807 ) | ( _27951 ) | ( _27952 ) ;
 assign wire15816 = ( n_n2821 ) | ( n_n2907 ) | ( wire15813 ) ;
 assign wire15817 = ( n_n2906 ) | ( n_n2908 ) | ( n_n2902 ) | ( wire15677 ) ;
 assign n_n1784 = ( n_n1789 ) | ( n_n1790 ) | ( wire16240 ) | ( wire16241 ) ;
 assign wire16323 = ( wire15902 ) | ( wire15903 ) | ( wire15943 ) | ( wire16320 ) ;
 assign wire16324 = ( n_n1793 ) | ( n_n1792 ) | ( n_n1794 ) | ( n_n1787 ) ;
 assign wire16830 = ( n_n2087 ) | ( n_n2086 ) | ( n_n2166 ) | ( wire16827 ) ;
 assign wire16831 = ( n_n2162 ) | ( n_n2163 ) | ( wire16470 ) | ( wire16829 ) ;
 assign n_n1038 = ( n_n1111 ) | ( wire11511 ) | ( wire11512 ) | ( wire11518 ) ;
 assign wire11502 = ( wire11491 ) | ( wire11492 ) | ( wire11496 ) | ( wire11497 ) ;
 assign n_n1014 = ( n_n1038 ) | ( wire11529 ) | ( _22972 ) | ( _22973 ) ;
 assign n_n942 = ( n_n953 ) | ( wire11653 ) | ( wire11654 ) | ( _23150 ) ;
 assign n_n941 = ( n_n951 ) | ( wire11675 ) | ( wire11676 ) | ( wire11690 ) ;
 assign n_n937 = ( n_n948 ) | ( n_n949 ) | ( wire11734 ) | ( wire11735 ) ;
 assign wire11745 = ( n_n956 ) | ( wire11660 ) | ( wire11661 ) | ( wire11743 ) ;
 assign n_n4309 = ( n_n942 ) | ( n_n941 ) | ( n_n937 ) | ( wire11745 ) ;
 assign n_n1012 = ( n_n1032 ) | ( _22149 ) | ( _22150 ) | ( _22151 ) ;
 assign wire11832 = ( n_n1077 ) | ( wire11829 ) | ( _22193 ) | ( _22194 ) ;
 assign n_n1007 = ( n_n1017 ) | ( _22550 ) | ( _22551 ) | ( _22552 ) ;
 assign n_n1009 = ( n_n1022 ) | ( wire12027 ) | ( _22691 ) | ( _22692 ) ;
 assign wire12036 = ( n_n1059 ) | ( wire12033 ) | ( _22732 ) | ( _22733 ) ;
 assign wire12037 = ( wire11909 ) | ( wire11978 ) | ( _22829 ) ;
 assign n_n1456 = ( n_n4983 ) | ( n_n4984 ) | ( wire57 ) | ( wire12156 ) ;
 assign n_n1455 = ( n_n4991 ) | ( n_n1576 ) | ( n_n5000 ) | ( wire12159 ) ;
 assign wire12197 = ( wire228 ) | ( wire362 ) | ( wire12196 ) ;
 assign wire12200 = ( wire12176 ) | ( wire12177 ) | ( wire12191 ) | ( wire12192 ) ;
 assign n_n1396 = ( n_n1456 ) | ( n_n1455 ) | ( wire12197 ) | ( wire12200 ) ;
 assign n_n1415 = ( n_n1467 ) | ( wire12239 ) | ( _24138 ) | ( _24139 ) ;
 assign wire12223 = ( n_n1985 ) | ( n_n3815 ) | ( wire12220 ) ;
 assign wire12224 = ( wire12213 ) | ( wire12214 ) | ( wire12218 ) | ( wire12219 ) ;
 assign wire12247 = ( n_n1472 ) | ( wire12204 ) | ( wire12205 ) | ( wire12245 ) ;
 assign n_n1397 = ( n_n1415 ) | ( wire12223 ) | ( wire12224 ) | ( wire12247 ) ;
 assign n_n1418 = ( n_n1478 ) | ( n_n1476 ) | ( wire12416 ) ;
 assign wire12432 = ( wire12420 ) | ( wire12421 ) | ( wire12425 ) | ( wire12426 ) ;
 assign n_n1398 = ( n_n1418 ) | ( wire12439 ) | ( _23821 ) | ( _23822 ) ;
 assign wire25 = ( (~ i_9_)  &  i_7_  &  i_8_  &  i_6_ ) ;
 assign n_n473 = ( i_5_  &  (~ i_3_)  &  (~ i_4_) ) ;
 assign n_n65 = ( (~ i_1_)  &  (~ i_2_)  &  (~ i_0_) ) ;
 assign n_n5305 = ( wire25  &  n_n473  &  n_n65 ) ;
 assign wire15 = ( (~ i_9_)  &  (~ i_7_)  &  i_8_  &  i_6_ ) ;
 assign n_n482 = ( (~ i_5_)  &  (~ i_3_)  &  i_4_ ) ;
 assign n_n5293 = ( n_n65  &  wire15  &  n_n482 ) ;
 assign wire19 = ( i_9_  &  (~ i_1_)  &  (~ i_2_)  &  (~ i_0_) ) ;
 assign n_n526 = ( i_7_  &  i_8_  &  (~ i_6_) ) ;
 assign n_n5296 = ( n_n482  &  wire19  &  n_n526 ) ;
 assign n_n522 = ( (~ i_7_)  &  i_8_  &  (~ i_6_) ) ;
 assign n_n491 = ( i_5_  &  (~ i_3_)  &  i_4_ ) ;
 assign n_n5284 = ( wire19  &  n_n522  &  n_n491 ) ;
 assign n_n559 = ( n_n4585 ) | ( n_n4592 ) | ( wire12595 ) | ( wire12596 ) ;
 assign wire12601 = ( n_n4648 ) | ( n_n4635 ) | ( wire140 ) | ( n_n4645 ) ;
 assign n_n543 = ( n_n559 ) | ( wire12607 ) | ( wire12608 ) | ( _25187 ) ;
 assign n_n4379 = ( n_n491  &  n_n536  &  wire24 ) ;
 assign n_n4399 = ( n_n482  &  n_n536  &  wire11 ) ;
 assign wire12699 = ( n_n4417 ) | ( n_n4371 ) | ( n_n4442 ) ;
 assign wire12700 = ( n_n4404 ) | ( n_n4441 ) | ( n_n4437 ) | ( n_n4384 ) ;
 assign n_n562 = ( n_n4379 ) | ( n_n4399 ) | ( wire12699 ) | ( wire12700 ) ;
 assign n_n4458 = ( n_n518  &  wire13  &  n_n532 ) ;
 assign n_n4488 = ( wire13  &  n_n534  &  n_n500 ) ;
 assign wire12706 = ( n_n4512 ) | ( n_n4453 ) | ( n_n4471 ) ;
 assign wire12707 = ( n_n4450 ) | ( n_n4460 ) | ( n_n4473 ) | ( n_n4506 ) ;
 assign n_n561 = ( n_n4458 ) | ( n_n4488 ) | ( wire12706 ) | ( wire12707 ) ;
 assign n_n4350 = ( wire16  &  n_n509  &  n_n528 ) ;
 assign n_n4331 = ( n_n518  &  n_n536  &  wire24 ) ;
 assign wire12713 = ( n_n4338 ) | ( n_n4327 ) | ( n_n4326 ) ;
 assign wire12714 = ( n_n4320 ) | ( n_n4315 ) | ( wire12710 ) ;
 assign n_n563 = ( n_n4350 ) | ( n_n4331 ) | ( wire12713 ) | ( wire12714 ) ;
 assign wire22 = ( (~ i_9_)  &  i_7_  &  i_8_  &  (~ i_6_) ) ;
 assign n_n5297 = ( n_n65  &  n_n482  &  wire22 ) ;
 assign n_n4378 = ( n_n491  &  wire16  &  n_n532 ) ;
 assign n_n4408 = ( n_n473  &  wire16  &  n_n534 ) ;
 assign wire13622 = ( n_n4388 ) | ( n_n4407 ) | ( n_n4402 ) ;
 assign wire13623 = ( n_n4399 ) | ( n_n4391 ) | ( n_n4371 ) | ( n_n4392 ) ;
 assign n_n3936 = ( n_n4378 ) | ( n_n4408 ) | ( wire13622 ) | ( wire13623 ) ;
 assign n_n3931 = ( n_n4701 ) | ( n_n4692 ) | ( wire13629 ) | ( wire13630 ) ;
 assign n_n3929 = ( n_n4901 ) | ( n_n4904 ) | ( wire13635 ) | ( wire13636 ) ;
 assign wire13643 = ( n_n4748 ) | ( n_n4725 ) | ( n_n4788 ) | ( n_n4802 ) ;
 assign wire13644 = ( n_n4765 ) | ( n_n4808 ) | ( n_n4742 ) | ( wire13638 ) ;
 assign n_n3920 = ( n_n3931 ) | ( n_n3929 ) | ( wire13643 ) | ( wire13644 ) ;
 assign n_n4362 = ( wire16  &  n_n532  &  n_n500 ) ;
 assign n_n4312 = ( wire16  &  n_n534  &  n_n535 ) ;
 assign wire13674 = ( wire15  &  n_n536  &  n_n535 ) | ( n_n536  &  n_n535  &  wire20 ) ;
 assign wire13679 = ( n_n4368 ) | ( n_n4358 ) | ( n_n4354 ) | ( wire124 ) ;
 assign n_n3194 = ( n_n5281 ) | ( n_n5268 ) | ( wire13709 ) | ( wire13710 ) ;
 assign wire13714 = ( wire13703 ) | ( wire13704 ) | ( wire13713 ) ;
 assign wire13728 = ( n_n5033 ) | ( n_n5051 ) | ( wire13725 ) | ( wire13726 ) ;
 assign wire13729 = ( wire13696 ) | ( wire13697 ) | ( wire13719 ) | ( wire13720 ) ;
 assign n_n3187 = ( n_n3194 ) | ( wire13714 ) | ( wire13728 ) | ( wire13729 ) ;
 assign n_n3202 = ( n_n4767 ) | ( n_n4752 ) | ( wire13746 ) | ( wire13747 ) ;
 assign wire13760 = ( n_n4663 ) | ( n_n4685 ) | ( n_n4696 ) | ( wire13755 ) ;
 assign n_n3192 = ( n_n3202 ) | ( wire13753 ) | ( _26577 ) | ( _26585 ) ;
 assign n_n3201 = ( n_n4839 ) | ( n_n4844 ) | ( wire13772 ) | ( wire13773 ) ;
 assign wire13767 = ( n_n4977 ) | ( n_n4920 ) | ( n_n4922 ) | ( n_n4959 ) ;
 assign wire13768 = ( n_n4913 ) | ( n_n4914 ) | ( n_n4953 ) | ( wire13765 ) ;
 assign wire13782 = ( wire13776 ) | ( wire13777 ) | ( wire13779 ) | ( _26606 ) ;
 assign n_n3191 = ( n_n3201 ) | ( wire13767 ) | ( wire13768 ) | ( wire13782 ) ;
 assign n_n3629 = ( n_n3650 ) | ( wire14419 ) | ( wire14420 ) | ( wire14436 ) ;
 assign wire14513 = ( n_n3736 ) | ( wire14466 ) | ( wire14467 ) | ( wire14511 ) ;
 assign wire14514 = ( wire14489 ) | ( wire14490 ) | ( wire14507 ) | ( wire14508 ) ;
 assign wire14540 = ( n_n3653 ) | ( n_n3655 ) | ( wire14536 ) | ( wire14537 ) ;
 assign n_n3635 = ( n_n3670 ) | ( wire14624 ) | ( wire14625 ) | ( wire14629 ) ;
 assign wire14614 = ( n_n3051 ) | ( wire14605 ) | ( wire14606 ) | ( wire14609 ) ;
 assign n_n3624 = ( n_n3635 ) | ( wire14637 ) | ( _27137 ) | ( _27138 ) ;
 assign n_n3639 = ( n_n3681 ) | ( wire14661 ) | ( wire14662 ) | ( wire14667 ) ;
 assign wire14655 = ( wire14644 ) | ( wire14645 ) | ( wire14648 ) | ( wire14649 ) ;
 assign wire14684 = ( wire14680 ) | ( wire14681 ) | ( wire14683 ) ;
 assign n_n3641 = ( n_n3689 ) | ( wire14760 ) | ( wire14761 ) | ( wire14764 ) ;
 assign wire14750 = ( n_n4917 ) | ( n_n4914 ) | ( wire14747 ) | ( wire14748 ) ;
 assign wire14751 = ( wire12168 ) | ( wire12169 ) | ( wire14742 ) | ( wire14743 ) ;
 assign wire14772 = ( n_n3694 ) | ( wire14738 ) | ( wire14739 ) | ( wire14770 ) ;
 assign n_n3626 = ( n_n3641 ) | ( wire14750 ) | ( wire14751 ) | ( wire14772 ) ;
 assign n_n524 = ( i_7_  &  (~ i_8_)  &  (~ i_6_) ) ;
 assign n_n464 = ( (~ i_5_)  &  (~ i_3_)  &  (~ i_4_) ) ;
 assign wire148 = ( i_9_  &  n_n65  &  n_n524  &  n_n464 ) | ( (~ i_9_)  &  n_n65  &  n_n524  &  n_n464 ) ;
 assign n_n2548 = ( n_n2601 ) | ( n_n2602 ) | ( wire14904 ) | ( wire14905 ) ;
 assign wire14935 = ( n_n2597 ) | ( wire14910 ) | ( wire14911 ) | ( wire14933 ) ;
 assign n_n2530 = ( n_n2548 ) | ( wire14935 ) | ( wire14927 ) | ( _27582 ) ;
 assign n_n2551 = ( n_n2611 ) | ( wire15011 ) | ( wire15012 ) | ( wire15016 ) ;
 assign wire15006 = ( wire14995 ) | ( wire14996 ) | ( wire15000 ) | ( wire15001 ) ;
 assign n_n2531 = ( n_n2551 ) | ( wire15024 ) | ( _27702 ) | ( _27703 ) ;
 assign n_n2533 = ( n_n2558 ) | ( wire15094 ) | ( wire15095 ) | ( wire15103 ) ;
 assign wire15150 = ( wire82 ) | ( wire224 ) | ( wire15143 ) | ( wire15149 ) ;
 assign wire15151 = ( wire15121 ) | ( wire15122 ) | ( wire15140 ) | ( wire15141 ) ;
 assign wire15169 = ( n_n2560 ) | ( n_n2559 ) | ( wire15165 ) | ( wire15166 ) ;
 assign n_n2528 = ( n_n2541 ) | ( wire15263 ) | ( _27452 ) | ( _27453 ) ;
 assign wire15206 = ( wire15192 ) | ( wire15203 ) | ( _27469 ) | ( _27470 ) ;
 assign n_n4436 = ( n_n522  &  n_n464  &  wire16 ) ;
 assign n_n4417 = ( n_n473  &  wire22  &  n_n536 ) ;
 assign wire15307 = ( n_n4371 ) | ( n_n4431 ) | ( n_n4424 ) ;
 assign wire15308 = ( n_n4384 ) | ( n_n4397 ) | ( wire15304 ) ;
 assign n_n2845 = ( n_n4436 ) | ( n_n4417 ) | ( wire15307 ) | ( wire15308 ) ;
 assign n_n4355 = ( wire21  &  n_n536  &  n_n509 ) ;
 assign n_n4335 = ( n_n518  &  n_n536  &  wire11 ) ;
 assign wire15321 = ( n_n4316 ) | ( n_n4345 ) | ( n_n4319 ) ;
 assign wire15322 = ( n_n4320 ) | ( n_n4357 ) | ( n_n4315 ) | ( n_n4348 ) ;
 assign n_n2846 = ( n_n4355 ) | ( n_n4335 ) | ( wire15321 ) | ( wire15322 ) ;
 assign n_n2841 = ( n_n4691 ) | ( n_n4686 ) | ( wire15333 ) | ( wire15334 ) ;
 assign wire15328 = ( n_n4598 ) | ( n_n4570 ) | ( n_n4612 ) | ( n_n4572 ) ;
 assign n_n2827 = ( n_n2841 ) | ( wire15340 ) | ( wire15341 ) | ( _28058 ) ;
 assign n_n2837 = ( wire15348 ) | ( wire15349 ) ;
 assign n_n2824 = ( n_n2832 ) | ( n_n2834 ) | ( wire15367 ) | ( wire15368 ) ;
 assign n_n2835 = ( n_n4986 ) | ( n_n4980 ) | ( wire15389 ) | ( wire15390 ) ;
 assign wire15400 = ( wire15385 ) | ( wire15396 ) | ( wire15397 ) | ( _27996 ) ;
 assign n_n2821 = ( n_n2837 ) | ( n_n2824 ) | ( n_n2835 ) | ( wire15400 ) ;
 assign n_n2839 = ( n_n4778 ) | ( n_n4745 ) | ( wire15405 ) | ( wire15406 ) ;
 assign wire15412 = ( n_n4854 ) | ( n_n4843 ) | ( wire150 ) ;
 assign wire15413 = ( wire40 ) | ( n_n4872 ) | ( n_n4852 ) | ( n_n4826 ) ;
 assign wire15418 = ( n_n4718 ) | ( n_n4700 ) | ( n_n1760 ) | ( wire15416 ) ;
 assign n_n2826 = ( n_n2839 ) | ( wire15412 ) | ( wire15413 ) | ( wire15418 ) ;
 assign n_n2929 = ( n_n2997 ) | ( n_n2996 ) | ( wire15451 ) | ( wire15452 ) ;
 assign wire15437 = ( n_n4510 ) | ( wire14200 ) | ( wire15434 ) | ( wire15435 ) ;
 assign wire15438 = ( wire11511 ) | ( wire11512 ) | ( wire15431 ) | ( wire15432 ) ;
 assign wire15463 = ( n_n3001 ) | ( n_n3003 ) | ( wire15459 ) | ( wire15460 ) ;
 assign n_n2907 = ( n_n2929 ) | ( wire15437 ) | ( wire15438 ) | ( wire15463 ) ;
 assign wire15501 = ( n_n4561 ) | ( n_n4556 ) | ( wire15498 ) | ( wire15499 ) ;
 assign wire15502 = ( wire15474 ) | ( wire15475 ) | ( wire15478 ) | ( wire15479 ) ;
 assign wire15504 = ( wire15472 ) | ( wire15495 ) | ( _28137 ) ;
 assign n_n2906 = ( wire15501 ) | ( wire15502 ) | ( wire15504 ) ;
 assign n_n2934 = ( n_n3012 ) | ( wire15525 ) | ( wire15526 ) | ( _28151 ) ;
 assign wire15543 = ( n_n4409 ) | ( n_n4410 ) | ( wire15538 ) | ( wire15542 ) ;
 assign wire15544 = ( wire15532 ) | ( wire15533 ) | ( wire15536 ) | ( wire15537 ) ;
 assign wire15549 = ( wire15507 ) | ( n_n3009 ) | ( _28175 ) | ( _28185 ) ;
 assign n_n2908 = ( n_n2934 ) | ( wire15543 ) | ( wire15544 ) | ( wire15549 ) ;
 assign n_n2905 = ( n_n2925 ) | ( wire15766 ) | ( wire15767 ) | ( wire15786 ) ;
 assign wire15743 = ( wire15715 ) | ( wire15729 ) | ( _27906 ) ;
 assign wire16025 = ( n_n4500 ) | ( n_n4508 ) | ( wire16022 ) | ( wire16023 ) ;
 assign wire16028 = ( wire16007 ) | ( wire16008 ) | ( wire16018 ) | ( wire16019 ) ;
 assign n_n1793 = ( wire16025 ) | ( wire16028 ) | ( _28704 ) ;
 assign n_n1813 = ( n_n1877 ) | ( wire16040 ) | ( wire16041 ) | ( wire16048 ) ;
 assign n_n1812 = ( n_n1872 ) | ( wire16064 ) | ( _28734 ) | ( _28735 ) ;
 assign wire16072 = ( n_n1879 ) | ( wire16069 ) | ( _28749 ) | ( _28750 ) ;
 assign n_n1792 = ( n_n1813 ) | ( n_n1812 ) | ( wire16072 ) ;
 assign n_n1818 = ( wire16099 ) | ( wire16105 ) | ( _28757 ) | ( _28767 ) ;
 assign wire16086 = ( n_n4329 ) | ( wire16083 ) | ( _25342 ) | ( _28771 ) ;
 assign wire16087 = ( wire16077 ) | ( wire16078 ) | ( wire16081 ) | ( wire16082 ) ;
 assign wire16114 = ( wire16112 ) | ( _28786 ) | ( _28787 ) | ( _28794 ) ;
 assign n_n1794 = ( n_n1818 ) | ( wire16086 ) | ( wire16087 ) | ( wire16114 ) ;
 assign n_n1789 = ( n_n1805 ) | ( wire16179 ) | ( _28361 ) | ( _28362 ) ;
 assign n_n1790 = ( n_n1808 ) | ( wire16213 ) | ( wire16214 ) | ( wire16224 ) ;
 assign wire16240 = ( wire16233 ) | ( wire16238 ) | ( _28416 ) | ( _28422 ) ;
 assign wire16241 = ( wire16130 ) | ( wire16131 ) | ( wire16144 ) | ( wire16145 ) ;
 assign n_n1797 = ( n_n1828 ) | ( wire16278 ) | ( wire16279 ) | ( _28812 ) ;
 assign wire16263 = ( wire16253 ) | ( wire16254 ) | ( wire16257 ) | ( wire16258 ) ;
 assign n_n1787 = ( n_n1797 ) | ( wire16288 ) | ( _28838 ) | ( _28839 ) ;
 assign wire16316 = ( wire16297 ) | ( wire16312 ) | ( _28589 ) ;
 assign wire16318 = ( wire117 ) | ( wire16308 ) | ( wire16309 ) | ( wire16313 ) ;
 assign n_n1786 = ( wire16316 ) | ( wire16318 ) | ( _28605 ) ;
 assign n_n4404 = ( n_n482  &  n_n522  &  wire16 ) ;
 assign n_n4413 = ( n_n473  &  wire15  &  n_n536 ) ;
 assign wire16475 = ( n_n4416 ) | ( n_n4405 ) | ( n_n4406 ) ;
 assign wire16476 = ( n_n4400 ) | ( n_n4389 ) | ( n_n4420 ) | ( n_n4407 ) ;
 assign n_n2104 = ( n_n4404 ) | ( n_n4413 ) | ( wire16475 ) | ( wire16476 ) ;
 assign wire16492 = ( _90 ) | ( wire15  &  n_n464  &  n_n455 ) ;
 assign wire16493 = ( n_n4571 ) | ( n_n4523 ) | ( n_n4553 ) ;
 assign wire16494 = ( n_n4521 ) | ( n_n4544 ) | ( wire16490 ) ;
 assign wire16497 = ( wire16482 ) | ( wire16483 ) | ( wire16487 ) | ( wire16488 ) ;
 assign n_n2087 = ( wire16492 ) | ( wire16493 ) | ( wire16494 ) | ( wire16497 ) ;
 assign n_n2099 = ( n_n4674 ) | ( n_n4661 ) | ( wire16508 ) | ( wire16509 ) ;
 assign wire16503 = ( n_n4710 ) | ( n_n4719 ) | ( wire16500 ) ;
 assign wire16504 = ( n_n4706 ) | ( n_n4699 ) | ( n_n4687 ) | ( wire16498 ) ;
 assign wire16516 = ( n_n2130 ) | ( n_n4811 ) | ( n_n4781 ) | ( wire16514 ) ;
 assign n_n2086 = ( n_n2099 ) | ( wire16503 ) | ( wire16504 ) | ( wire16516 ) ;
 assign n_n2190 = ( n_n2263 ) | ( wire16531 ) | ( _29006 ) | ( _29007 ) ;
 assign wire16545 = ( n_n2446 ) | ( n_n2443 ) | ( n_n2445 ) | ( wire16539 ) ;
 assign n_n2166 = ( n_n2190 ) | ( wire16556 ) | ( _29028 ) | ( _29029 ) ;
 assign n_n4367 = ( n_n536  &  wire11  &  n_n500 ) ;
 assign n_n4374 = ( wire16  &  n_n520  &  n_n500 ) ;
 assign wire16651 = ( n_n4338 ) | ( n_n4325 ) | ( n_n4380 ) | ( n_n4345 ) ;
 assign wire16745 = ( wire16715 ) | ( wire16716 ) | ( wire16730 ) | ( wire16731 ) ;
 assign wire16763 = ( wire16758 ) | ( wire16662 ) | ( _28934 ) | ( _28949 ) ;
 assign wire16 = ( i_9_  &  i_1_  &  i_2_  &  i_0_ ) ;
 assign n_n518 = ( (~ i_5_)  &  i_3_  &  i_4_ ) ;
 assign n_n4338 = ( n_n524  &  wire16  &  n_n518 ) ;
 assign wire21 = ( (~ i_9_)  &  i_7_  &  (~ i_8_)  &  (~ i_6_) ) ;
 assign n_n536 = ( i_1_  &  i_2_  &  i_0_ ) ;
 assign n_n4339 = ( n_n518  &  wire21  &  n_n536 ) ;
 assign n_n4337 = ( wire22  &  n_n518  &  n_n536 ) ;
 assign n_n4401 = ( n_n482  &  wire22  &  n_n536 ) ;
 assign n_n4403 = ( n_n482  &  wire21  &  n_n536 ) ;
 assign n_n4400 = ( n_n482  &  n_n526  &  wire16 ) ;
 assign wire13 = ( i_9_  &  i_1_  &  (~ i_2_)  &  i_0_ ) ;
 assign n_n4464 = ( n_n526  &  n_n518  &  wire13 ) ;
 assign n_n455 = ( i_1_  &  (~ i_2_)  &  i_0_ ) ;
 assign n_n4467 = ( n_n518  &  wire21  &  n_n455 ) ;
 assign wire11 = ( (~ i_9_)  &  (~ i_7_)  &  (~ i_8_)  &  i_6_ ) ;
 assign n_n4463 = ( n_n518  &  n_n455  &  wire11 ) ;
 assign wire10 = ( i_9_  &  (~ i_1_)  &  i_2_  &  i_0_ ) ;
 assign n_n532 = ( i_7_  &  (~ i_8_)  &  i_6_ ) ;
 assign n_n4666 = ( n_n473  &  wire10  &  n_n532 ) ;
 assign wire24 = ( (~ i_9_)  &  i_7_  &  (~ i_8_)  &  i_6_ ) ;
 assign n_n390 = ( (~ i_1_)  &  i_2_  &  i_0_ ) ;
 assign n_n4667 = ( n_n473  &  wire24  &  n_n390 ) ;
 assign n_n534 = ( i_7_  &  i_8_  &  i_6_ ) ;
 assign n_n4664 = ( n_n473  &  wire10  &  n_n534 ) ;
 assign n_n509 = ( i_5_  &  i_3_  &  (~ i_4_) ) ;
 assign n_n325 = ( (~ i_1_)  &  (~ i_2_)  &  i_0_ ) ;
 assign n_n4737 = ( wire22  &  n_n509  &  n_n325 ) ;
 assign wire14 = ( i_9_  &  (~ i_1_)  &  (~ i_2_)  &  i_0_ ) ;
 assign n_n4738 = ( n_n524  &  n_n509  &  wire14 ) ;
 assign n_n4735 = ( wire11  &  n_n509  &  n_n325 ) ;
 assign n_n528 = ( (~ i_7_)  &  (~ i_8_)  &  i_6_ ) ;
 assign n_n4782 = ( n_n482  &  wire14  &  n_n528 ) ;
 assign n_n4784 = ( n_n482  &  n_n526  &  wire14 ) ;
 assign n_n4779 = ( n_n482  &  wire24  &  n_n325 ) ;
 assign wire17 = ( i_9_  &  i_1_  &  i_2_  &  (~ i_0_) ) ;
 assign n_n535 = ( i_5_  &  i_3_  &  i_4_ ) ;
 assign n_n4830 = ( n_n528  &  wire17  &  n_n535 ) ;
 assign n_n260 = ( i_1_  &  i_2_  &  (~ i_0_) ) ;
 assign n_n4831 = ( wire11  &  n_n535  &  n_n260 ) ;
 assign n_n4900 = ( n_n522  &  n_n491  &  wire17 ) ;
 assign n_n520 = ( (~ i_7_)  &  (~ i_8_)  &  (~ i_6_) ) ;
 assign n_n4902 = ( n_n491  &  wire17  &  n_n520 ) ;
 assign n_n4898 = ( n_n491  &  n_n524  &  wire17 ) ;
 assign wire18 = ( i_9_  &  i_1_  &  (~ i_2_)  &  (~ i_0_) ) ;
 assign n_n4976 = ( n_n526  &  n_n518  &  wire18 ) ;
 assign n_n195 = ( i_1_  &  (~ i_2_)  &  (~ i_0_) ) ;
 assign n_n4977 = ( wire22  &  n_n518  &  n_n195 ) ;
 assign n_n4975 = ( n_n518  &  wire11  &  n_n195 ) ;
 assign n_n5038 = ( n_n482  &  n_n528  &  wire18 ) ;
 assign n_n5040 = ( n_n482  &  n_n526  &  wire18 ) ;
 assign n_n5034 = ( n_n482  &  n_n532  &  wire18 ) ;
 assign wire12 = ( i_9_  &  (~ i_1_)  &  i_2_  &  (~ i_0_) ) ;
 assign n_n5092 = ( n_n522  &  n_n535  &  wire12 ) ;
 assign wire20 = ( (~ i_9_)  &  (~ i_7_)  &  i_8_  &  (~ i_6_) ) ;
 assign n_n130 = ( (~ i_1_)  &  i_2_  &  (~ i_0_) ) ;
 assign n_n5093 = ( n_n535  &  wire20  &  n_n130 ) ;
 assign n_n5091 = ( wire21  &  n_n535  &  n_n130 ) ;
 assign n_n4440 = ( wire13  &  n_n534  &  n_n535 ) ;
 assign n_n4434 = ( n_n524  &  n_n464  &  wire16 ) ;
 assign n_n4432 = ( n_n526  &  n_n464  &  wire16 ) ;
 assign wire98 = ( wire22  &  n_n464  &  n_n536 ) | ( n_n464  &  n_n536  &  wire11 ) ;
 assign wire233 = ( i_9_  &  n_n464  &  n_n536  &  n_n520 ) | ( (~ i_9_)  &  n_n464  &  n_n536  &  n_n520 ) ;
 assign wire236 = ( i_9_  &  n_n522  &  n_n464  &  n_n536 ) | ( (~ i_9_)  &  n_n522  &  n_n464  &  n_n536 ) ;
 assign n_n4720 = ( n_n526  &  n_n518  &  wire14 ) ;
 assign n_n4718 = ( n_n518  &  wire14  &  n_n528 ) ;
 assign n_n4717 = ( wire15  &  n_n518  &  n_n325 ) ;
 assign n_n4857 = ( wire25  &  n_n509  &  n_n260 ) ;
 assign n_n4862 = ( n_n509  &  n_n528  &  wire17 ) ;
 assign n_n4856 = ( n_n534  &  n_n509  &  wire17 ) ;
 assign wire40 = ( wire22  &  n_n509  &  n_n260 ) | ( wire11  &  n_n509  &  n_n260 ) ;
 assign wire102 = ( i_9_  &  n_n518  &  n_n260  &  n_n520 ) | ( (~ i_9_)  &  n_n518  &  n_n260  &  n_n520 ) ;
 assign wire245 = ( i_9_  &  n_n532  &  n_n509  &  n_n260 ) | ( (~ i_9_)  &  n_n532  &  n_n509  &  n_n260 ) ;
 assign n_n4991 = ( wire11  &  n_n509  &  n_n195 ) ;
 assign n_n4996 = ( n_n522  &  n_n509  &  wire18 ) ;
 assign n_n4992 = ( n_n526  &  n_n509  &  wire18 ) ;
 assign n_n4995 = ( wire21  &  n_n509  &  n_n195 ) ;
 assign n_n4990 = ( n_n509  &  n_n528  &  wire18 ) ;
 assign n_n4998 = ( n_n509  &  n_n520  &  wire18 ) ;
 assign wire23 = ( (~ i_9_)  &  (~ i_7_)  &  (~ i_8_)  &  (~ i_6_) ) ;
 assign n_n4999 = ( n_n509  &  n_n195  &  wire23 ) ;
 assign n_n500 = ( (~ i_5_)  &  i_3_  &  (~ i_4_) ) ;
 assign wire103 = ( i_9_  &  n_n534  &  n_n195  &  n_n500 ) | ( (~ i_9_)  &  n_n534  &  n_n195  &  n_n500 ) ;
 assign n_n4617 = ( wire25  &  n_n390  &  n_n500 ) ;
 assign n_n4637 = ( wire15  &  n_n491  &  n_n390 ) ;
 assign n_n4613 = ( n_n390  &  n_n509  &  wire20 ) ;
 assign n_n4927 = ( n_n473  &  wire11  &  n_n260 ) ;
 assign n_n4958 = ( n_n528  &  n_n535  &  wire18 ) ;
 assign n_n4920 = ( n_n473  &  n_n534  &  wire17 ) ;
 assign n_n4325 = ( n_n536  &  n_n535  &  wire20 ) ;
 assign n_n4327 = ( n_n536  &  n_n535  &  wire23 ) ;
 assign n_n4324 = ( n_n522  &  wire16  &  n_n535 ) ;
 assign n_n4382 = ( n_n491  &  wire16  &  n_n528 ) ;
 assign n_n4383 = ( n_n491  &  n_n536  &  wire11 ) ;
 assign n_n530 = ( (~ i_7_)  &  i_8_  &  i_6_ ) ;
 assign n_n4380 = ( n_n491  &  wire16  &  n_n530 ) ;
 assign n_n4923 = ( n_n473  &  wire24  &  n_n260 ) ;
 assign n_n4924 = ( n_n473  &  wire17  &  n_n530 ) ;
 assign n_n4921 = ( wire25  &  n_n473  &  n_n260 ) ;
 assign n_n4982 = ( n_n518  &  n_n520  &  wire18 ) ;
 assign n_n4983 = ( n_n518  &  n_n195  &  wire23 ) ;
 assign n_n4981 = ( n_n518  &  n_n195  &  wire20 ) ;
 assign n_n5035 = ( n_n482  &  wire24  &  n_n195 ) ;
 assign n_n5032 = ( n_n482  &  n_n534  &  wire18 ) ;
 assign n_n5111 = ( n_n518  &  n_n130  &  wire23 ) ;
 assign n_n5112 = ( n_n534  &  n_n509  &  wire12 ) ;
 assign n_n5109 = ( n_n518  &  wire20  &  n_n130 ) ;
 assign n_n5171 = ( n_n482  &  wire21  &  n_n130 ) ;
 assign n_n5174 = ( n_n482  &  n_n520  &  wire12 ) ;
 assign n_n5167 = ( n_n482  &  wire11  &  n_n130 ) ;
 assign n_n4597 = ( n_n518  &  n_n390  &  wire20 ) ;
 assign n_n4598 = ( n_n518  &  wire10  &  n_n520 ) ;
 assign n_n4602 = ( wire10  &  n_n532  &  n_n509 ) ;
 assign n_n4593 = ( wire22  &  n_n518  &  n_n390 ) ;
 assign n_n4601 = ( wire25  &  n_n390  &  n_n509 ) ;
 assign wire108 = ( i_9_  &  n_n390  &  n_n509  &  n_n530 ) | ( (~ i_9_)  &  n_n390  &  n_n509  &  n_n530 ) ;
 assign n_n4744 = ( n_n534  &  wire14  &  n_n500 ) ;
 assign n_n4754 = ( n_n524  &  wire14  &  n_n500 ) ;
 assign n_n4757 = ( n_n325  &  wire20  &  n_n500 ) ;
 assign n_n4749 = ( wire15  &  n_n325  &  n_n500 ) ;
 assign n_n4756 = ( n_n522  &  wire14  &  n_n500 ) ;
 assign wire109 = ( i_9_  &  n_n325  &  n_n528  &  n_n500 ) | ( (~ i_9_)  &  n_n325  &  n_n528  &  n_n500 ) ;
 assign n_n4887 = ( n_n260  &  wire23  &  n_n500 ) ;
 assign n_n4888 = ( n_n491  &  n_n534  &  wire17 ) ;
 assign n_n4885 = ( n_n260  &  wire20  &  n_n500 ) ;
 assign n_n3450 = ( n_n4887 ) | ( n_n4888 ) | ( n_n4885 ) ;
 assign n_n4882 = ( n_n524  &  wire17  &  n_n500 ) ;
 assign n_n4884 = ( n_n522  &  wire17  &  n_n500 ) ;
 assign n_n4883 = ( wire21  &  n_n260  &  n_n500 ) ;
 assign n_n5026 = ( n_n491  &  n_n524  &  wire18 ) ;
 assign n_n5027 = ( n_n491  &  wire21  &  n_n195 ) ;
 assign n_n5025 = ( n_n491  &  wire22  &  n_n195 ) ;
 assign wire114 = ( i_9_  &  n_n473  &  n_n532  &  n_n130 ) | ( (~ i_9_)  &  n_n473  &  n_n532  &  n_n130 ) ;
 assign n_n5181 = ( n_n473  &  wire15  &  n_n130 ) ;
 assign n_n5184 = ( n_n473  &  n_n526  &  wire12 ) ;
 assign n_n5183 = ( n_n473  &  wire11  &  n_n130 ) ;
 assign wire112 = ( i_9_  &  n_n473  &  n_n524  &  n_n130 ) | ( (~ i_9_)  &  n_n473  &  n_n524  &  n_n130 ) ;
 assign n_n5318 = ( n_n473  &  wire19  &  n_n520 ) ;
 assign n_n5314 = ( n_n473  &  wire19  &  n_n524 ) ;
 assign n_n5320 = ( wire19  &  n_n464  &  n_n534 ) ;
 assign wire459 = ( i_9_  &  n_n473  &  n_n65  &  n_n526 ) | ( (~ i_9_)  &  n_n473  &  n_n65  &  n_n526 ) ;
 assign n_n4615 = ( n_n390  &  n_n509  &  wire23 ) ;
 assign n_n4616 = ( wire10  &  n_n534  &  n_n500 ) ;
 assign n_n4607 = ( wire11  &  n_n390  &  n_n509 ) ;
 assign wire396 = ( n_n526  &  wire10  &  n_n509 ) | ( wire10  &  n_n509  &  n_n528 ) ;
 assign wire14071 = ( n_n4607 ) | ( n_n4612 ) | ( n_n4609 ) ;
 assign wire14072 = ( n_n4617 ) | ( n_n4613 ) | ( wire396 ) ;
 assign n_n3346 = ( n_n4615 ) | ( n_n4616 ) | ( wire14071 ) | ( wire14072 ) ;
 assign n_n4641 = ( n_n491  &  wire22  &  n_n390 ) ;
 assign n_n4634 = ( n_n491  &  wire10  &  n_n532 ) ;
 assign n_n4648 = ( n_n482  &  wire10  &  n_n534 ) ;
 assign n_n4618 = ( wire10  &  n_n532  &  n_n500 ) ;
 assign n_n4628 = ( n_n522  &  wire10  &  n_n500 ) ;
 assign wire26 = ( i_9_  &  n_n491  &  n_n390  &  n_n530 ) | ( (~ i_9_)  &  n_n491  &  n_n390  &  n_n530 ) ;
 assign wire118 = ( wire15  &  n_n390  &  n_n500 ) | ( wire24  &  n_n390  &  n_n500 ) ;
 assign wire309 = ( n_n491  &  wire21  &  n_n390 ) | ( n_n491  &  n_n390  &  wire20 ) ;
 assign wire14078 = ( n_n4639 ) | ( n_n4642 ) | ( n_n4631 ) | ( n_n4632 ) ;
 assign n_n3281 = ( n_n3346 ) | ( wire14079 ) | ( wire14080 ) | ( _26195 ) ;
 assign n_n5050 = ( n_n473  &  n_n532  &  wire18 ) ;
 assign n_n5060 = ( n_n473  &  n_n522  &  wire18 ) ;
 assign n_n5055 = ( n_n473  &  wire11  &  n_n195 ) ;
 assign n_n5054 = ( n_n473  &  n_n528  &  wire18 ) ;
 assign n_n5059 = ( n_n473  &  wire21  &  n_n195 ) ;
 assign n_n5048 = ( n_n473  &  n_n534  &  wire18 ) ;
 assign n_n5028 = ( n_n522  &  n_n491  &  wire18 ) ;
 assign n_n5036 = ( n_n482  &  wire18  &  n_n530 ) ;
 assign wire50 = ( i_9_  &  n_n491  &  n_n520  &  n_n195 ) | ( (~ i_9_)  &  n_n491  &  n_n520  &  n_n195 ) ;
 assign n_n5039 = ( n_n482  &  wire11  &  n_n195 ) ;
 assign wire97 = ( i_9_  &  n_n482  &  n_n526  &  n_n195 ) | ( (~ i_9_)  &  n_n482  &  n_n526  &  n_n195 ) ;
 assign wire13983 = ( n_n482  &  n_n524  &  wire18 ) | ( n_n482  &  n_n528  &  wire18 ) ;
 assign wire231 = ( i_9_  &  n_n482  &  n_n532  &  n_n195 ) | ( (~ i_9_)  &  n_n482  &  n_n532  &  n_n195 ) ;
 assign wire356 = ( n_n482  &  n_n522  &  wire18 ) | ( n_n482  &  n_n520  &  wire18 ) ;
 assign n_n4571 = ( wire24  &  n_n390  &  n_n535 ) ;
 assign n_n4578 = ( n_n524  &  wire10  &  n_n535 ) ;
 assign n_n4570 = ( wire10  &  n_n532  &  n_n535 ) ;
 assign n_n4849 = ( wire22  &  n_n518  &  n_n260 ) ;
 assign n_n4853 = ( n_n518  &  n_n260  &  wire20 ) ;
 assign n_n4847 = ( n_n518  &  wire11  &  n_n260 ) ;
 assign n_n5096 = ( n_n518  &  n_n534  &  wire12 ) ;
 assign n_n5099 = ( n_n518  &  wire24  &  n_n130 ) ;
 assign n_n5085 = ( wire15  &  n_n535  &  n_n130 ) ;
 assign n_n4314 = ( wire16  &  n_n532  &  n_n535 ) ;
 assign n_n4389 = ( n_n491  &  n_n536  &  wire20 ) ;
 assign n_n4369 = ( wire22  &  n_n536  &  n_n500 ) ;
 assign n_n4381 = ( wire15  &  n_n491  &  n_n536 ) ;
 assign n_n4340 = ( n_n522  &  wire16  &  n_n518 ) ;
 assign wire280 = ( i_9_  &  n_n491  &  n_n536  &  n_n532 ) | ( (~ i_9_)  &  n_n491  &  n_n536  &  n_n532 ) ;
 assign n_n5101 = ( wire15  &  n_n518  &  n_n130 ) ;
 assign n_n5110 = ( n_n518  &  n_n520  &  wire12 ) ;
 assign n_n5142 = ( n_n520  &  wire12  &  n_n500 ) ;
 assign n_n5107 = ( n_n518  &  wire21  &  n_n130 ) ;
 assign n_n5130 = ( n_n532  &  wire12  &  n_n500 ) ;
 assign n_n5123 = ( wire21  &  n_n509  &  n_n130 ) ;
 assign n_n5129 = ( wire25  &  n_n130  &  n_n500 ) ;
 assign n_n5156 = ( n_n522  &  n_n491  &  wire12 ) ;
 assign n_n4317 = ( wire15  &  n_n536  &  n_n535 ) ;
 assign n_n4318 = ( wire16  &  n_n528  &  n_n535 ) ;
 assign n_n4388 = ( n_n522  &  n_n491  &  wire16 ) ;
 assign n_n4459 = ( n_n518  &  n_n455  &  wire24 ) ;
 assign n_n4461 = ( wire15  &  n_n518  &  n_n455 ) ;
 assign n_n4455 = ( n_n455  &  n_n535  &  wire23 ) ;
 assign n_n4513 = ( n_n491  &  wire22  &  n_n455 ) ;
 assign n_n4515 = ( n_n491  &  wire21  &  n_n455 ) ;
 assign n_n4512 = ( n_n526  &  n_n491  &  wire13 ) ;
 assign n_n4790 = ( n_n482  &  wire14  &  n_n520 ) ;
 assign n_n4791 = ( n_n482  &  n_n325  &  wire23 ) ;
 assign n_n4787 = ( n_n482  &  wire21  &  n_n325 ) ;
 assign n_n4859 = ( wire24  &  n_n509  &  n_n260 ) ;
 assign n_n4860 = ( n_n509  &  wire17  &  n_n530 ) ;
 assign n_n4858 = ( n_n532  &  n_n509  &  wire17 ) ;
 assign n_n4926 = ( n_n473  &  n_n528  &  wire17 ) ;
 assign n_n4928 = ( n_n473  &  n_n526  &  wire17 ) ;
 assign n_n4925 = ( n_n473  &  wire15  &  n_n260 ) ;
 assign n_n4988 = ( n_n509  &  wire18  &  n_n530 ) ;
 assign n_n4987 = ( wire24  &  n_n509  &  n_n195 ) ;
 assign n_n5041 = ( n_n482  &  wire22  &  n_n195 ) ;
 assign n_n5042 = ( n_n482  &  n_n524  &  wire18 ) ;
 assign n_n5100 = ( n_n518  &  wire12  &  n_n530 ) ;
 assign n_n4724 = ( n_n522  &  n_n518  &  wire14 ) ;
 assign n_n4727 = ( n_n518  &  n_n325  &  wire23 ) ;
 assign n_n4739 = ( wire21  &  n_n509  &  n_n325 ) ;
 assign wire95 = ( i_9_  &  n_n509  &  n_n325  &  n_n528 ) | ( (~ i_9_)  &  n_n509  &  n_n325  &  n_n528 ) ;
 assign wire244 = ( n_n532  &  n_n509  &  wire14 ) | ( n_n534  &  n_n509  &  wire14 ) ;
 assign n_n4864 = ( n_n526  &  n_n509  &  wire17 ) ;
 assign n_n4868 = ( n_n522  &  n_n509  &  wire17 ) ;
 assign n_n5018 = ( n_n491  &  n_n532  &  wire18 ) ;
 assign n_n5022 = ( n_n491  &  n_n528  &  wire18 ) ;
 assign n_n5017 = ( wire25  &  n_n491  &  n_n195 ) ;
 assign wire135 = ( i_9_  &  n_n520  &  n_n195  &  n_n500 ) | ( (~ i_9_)  &  n_n520  &  n_n195  &  n_n500 ) ;
 assign wire296 = ( wire15  &  n_n491  &  n_n195 ) | ( n_n491  &  wire11  &  n_n195 ) ;
 assign n_n4993 = ( wire22  &  n_n509  &  n_n195 ) ;
 assign n_n4994 = ( n_n524  &  n_n509  &  wire18 ) ;
 assign n_n1576 = ( n_n4996 ) | ( n_n4995 ) | ( n_n4994 ) ;
 assign wire134 = ( i_9_  &  n_n509  &  n_n195  &  n_n530 ) | ( (~ i_9_)  &  n_n509  &  n_n195  &  n_n530 ) ;
 assign wire252 = ( n_n522  &  n_n518  &  wire18 ) | ( n_n518  &  n_n520  &  wire18 ) ;
 assign n_n5005 = ( wire15  &  n_n195  &  n_n500 ) ;
 assign n_n5004 = ( wire18  &  n_n500  &  n_n530 ) ;
 assign n_n5000 = ( n_n534  &  wire18  &  n_n500 ) ;
 assign wire136 = ( i_9_  &  n_n528  &  n_n195  &  n_n500 ) | ( (~ i_9_)  &  n_n528  &  n_n195  &  n_n500 ) ;
 assign wire393 = ( i_9_  &  n_n532  &  n_n195  &  n_n500 ) | ( (~ i_9_)  &  n_n532  &  n_n195  &  n_n500 ) ;
 assign n_n4907 = ( n_n482  &  wire24  &  n_n260 ) ;
 assign n_n4913 = ( n_n482  &  wire22  &  n_n260 ) ;
 assign n_n4922 = ( n_n473  &  n_n532  &  wire17 ) ;
 assign n_n4934 = ( n_n473  &  wire17  &  n_n520 ) ;
 assign wire14801 = ( _348 ) | ( n_n482  &  wire19  &  n_n530 ) ;
 assign wire14802 = ( n_n5284 ) | ( n_n5240 ) | ( n_n5248 ) ;
 assign wire14803 = ( n_n5245 ) | ( n_n5278 ) | ( n_n5287 ) | ( n_n5261 ) ;
 assign wire14807 = ( n_n5296 ) | ( n_n5320 ) | ( n_n5324 ) | ( n_n5335 ) ;
 assign n_n2451 = ( wire14801 ) | ( wire14802 ) | ( wire14803 ) | ( wire14807 ) ;
 assign n_n4951 = ( n_n464  &  n_n260  &  wire23 ) ;
 assign n_n5010 = ( n_n524  &  wire18  &  n_n500 ) ;
 assign wire14810 = ( n_n535  &  n_n195  &  wire23 ) | ( n_n195  &  wire23  &  n_n500 ) ;
 assign wire14814 = ( n_n4985 ) | ( n_n4986 ) | ( n_n4962 ) | ( wire14808 ) ;
 assign n_n2462 = ( n_n4951 ) | ( n_n5010 ) | ( wire14810 ) | ( wire14814 ) ;
 assign n_n4886 = ( wire17  &  n_n520  &  n_n500 ) ;
 assign n_n4865 = ( wire22  &  n_n509  &  n_n260 ) ;
 assign wire14819 = ( n_n4847 ) | ( n_n4868 ) | ( n_n4871 ) ;
 assign n_n2464 = ( wire14819 ) | ( wire14816 ) | ( wire14817 ) | ( _27731 ) ;
 assign wire31 = ( i_9_  &  n_n473  &  n_n526  &  n_n260 ) | ( (~ i_9_)  &  n_n473  &  n_n526  &  n_n260 ) ;
 assign n_n4453 = ( n_n455  &  n_n535  &  wire20 ) ;
 assign n_n4420 = ( n_n473  &  n_n522  &  wire16 ) ;
 assign n_n4407 = ( n_n482  &  n_n536  &  wire23 ) ;
 assign n_n2470 = ( n_n4504 ) | ( n_n4525 ) | ( wire14838 ) | ( wire14839 ) ;
 assign wire14833 = ( wire118 ) | ( n_n4631 ) | ( n_n4632 ) ;
 assign wire14834 = ( wire396 ) | ( n_n4629 ) | ( wire14831 ) ;
 assign wire14848 = ( n_n4592 ) | ( n_n4556 ) | ( wire14845 ) | ( wire14846 ) ;
 assign n_n2455 = ( n_n2470 ) | ( wire14833 ) | ( wire14834 ) | ( wire14848 ) ;
 assign n_n2467 = ( n_n4665 ) | ( n_n4708 ) | ( wire14854 ) | ( wire14855 ) ;
 assign wire14861 = ( n_n4735 ) | ( n_n4724 ) | ( n_n4733 ) | ( n_n4725 ) ;
 assign wire14862 = ( n_n4760 ) | ( n_n4758 ) | ( n_n4714 ) | ( wire14859 ) ;
 assign wire14870 = ( n_n4805 ) | ( n_n4766 ) | ( wire14867 ) | ( wire14868 ) ;
 assign n_n2454 = ( n_n2467 ) | ( wire14861 ) | ( wire14862 ) | ( wire14870 ) ;
 assign n_n4391 = ( n_n491  &  n_n536  &  wire23 ) ;
 assign wire14875 = ( n_n4399 ) | ( n_n4396 ) | ( n_n4375 ) ;
 assign wire14876 = ( n_n4403 ) | ( n_n4382 ) | ( wire14873 ) ;
 assign n_n2472 = ( n_n4362 ) | ( n_n4391 ) | ( wire14875 ) | ( wire14876 ) ;
 assign n_n4316 = ( wire16  &  n_n535  &  n_n530 ) ;
 assign n_n4313 = ( wire25  &  n_n536  &  n_n535 ) ;
 assign wire14881 = ( n_n4330 ) | ( n_n4352 ) | ( n_n4351 ) ;
 assign wire14882 = ( n_n4318 ) | ( n_n4344 ) | ( n_n4320 ) | ( n_n4341 ) ;
 assign n_n2473 = ( n_n4316 ) | ( n_n4313 ) | ( wire14881 ) | ( wire14882 ) ;
 assign wire234 = ( wire13  &  n_n534  &  n_n535 ) | ( wire13  &  n_n535  &  n_n530 ) ;
 assign n_n4372 = ( n_n522  &  wire16  &  n_n500 ) ;
 assign n_n4373 = ( n_n536  &  wire20  &  n_n500 ) ;
 assign n_n4371 = ( wire21  &  n_n536  &  n_n500 ) ;
 assign n_n4431 = ( n_n464  &  n_n536  &  wire11 ) ;
 assign n_n4433 = ( wire22  &  n_n464  &  n_n536 ) ;
 assign n_n4430 = ( n_n464  &  wire16  &  n_n528 ) ;
 assign n_n4494 = ( wire13  &  n_n528  &  n_n500 ) ;
 assign n_n4491 = ( n_n455  &  wire24  &  n_n500 ) ;
 assign n_n4834 = ( n_n524  &  wire17  &  n_n535 ) ;
 assign n_n4835 = ( wire21  &  n_n535  &  n_n260 ) ;
 assign n_n4832 = ( n_n526  &  wire17  &  n_n535 ) ;
 assign n_n4909 = ( wire15  &  n_n482  &  n_n260 ) ;
 assign n_n4911 = ( n_n482  &  wire11  &  n_n260 ) ;
 assign n_n4903 = ( n_n491  &  n_n260  &  wire23 ) ;
 assign n_n4979 = ( n_n518  &  wire21  &  n_n195 ) ;
 assign n_n5049 = ( wire25  &  n_n473  &  n_n195 ) ;
 assign n_n5179 = ( n_n473  &  wire24  &  n_n130 ) ;
 assign n_n5239 = ( n_n65  &  n_n518  &  wire23 ) ;
 assign n_n5240 = ( wire19  &  n_n534  &  n_n509 ) ;
 assign n_n5238 = ( wire19  &  n_n518  &  n_n520 ) ;
 assign n_n4514 = ( n_n491  &  n_n524  &  wire13 ) ;
 assign wire791 = ( n_n522  &  n_n491  &  wire13 ) ;
 assign n_n4247 = ( n_n4515 ) | ( n_n4514 ) | ( wire791 ) ;
 assign n_n4646 = ( n_n491  &  wire10  &  n_n520 ) ;
 assign n_n4644 = ( n_n522  &  n_n491  &  wire10 ) ;
 assign n_n4651 = ( n_n482  &  wire24  &  n_n390 ) ;
 assign n_n4649 = ( wire25  &  n_n482  &  n_n390 ) ;
 assign wire311 = ( i_9_  &  n_n482  &  n_n390  &  n_n530 ) | ( (~ i_9_)  &  n_n482  &  n_n390  &  n_n530 ) ;
 assign n_n4952 = ( n_n534  &  n_n535  &  wire18 ) ;
 assign n_n4950 = ( n_n464  &  wire17  &  n_n520 ) ;
 assign n_n3803 = ( n_n4951 ) | ( n_n4952 ) | ( n_n4950 ) ;
 assign n_n4942 = ( n_n464  &  n_n528  &  wire17 ) ;
 assign wire59 = ( wire15  &  n_n464  &  n_n260 ) ;
 assign n_n4945 = ( wire22  &  n_n464  &  n_n260 ) ;
 assign n_n4946 = ( n_n524  &  n_n464  &  wire17 ) ;
 assign n_n4949 = ( n_n464  &  n_n260  &  wire20 ) ;
 assign wire12166 = ( i_9_  &  n_n464  &  n_n528  &  n_n260 ) | ( (~ i_9_)  &  n_n464  &  n_n528  &  n_n260 ) ;
 assign wire16327 = ( n_n4945 ) | ( n_n4946 ) | ( n_n4949 ) ;
 assign n_n2222 = ( n_n3803 ) | ( wire59 ) | ( wire12166 ) | ( wire16327 ) ;
 assign n_n5244 = ( wire19  &  n_n509  &  n_n530 ) ;
 assign n_n5245 = ( n_n65  &  wire15  &  n_n509 ) ;
 assign wire318 = ( i_9_  &  n_n65  &  n_n509  &  n_n528 ) | ( (~ i_9_)  &  n_n65  &  n_n509  &  n_n528 ) ;
 assign wire16686 = ( n_n5239 ) | ( n_n5240 ) | ( wire318 ) ;
 assign n_n4450 = ( n_n524  &  wire13  &  n_n535 ) ;
 assign n_n4445 = ( wire15  &  n_n455  &  n_n535 ) ;
 assign n_n4444 = ( wire13  &  n_n535  &  n_n530 ) ;
 assign n_n4442 = ( wire13  &  n_n532  &  n_n535 ) ;
 assign n_n4441 = ( wire25  &  n_n455  &  n_n535 ) ;
 assign wire368 = ( wire22  &  n_n455  &  n_n535 ) | ( wire21  &  n_n455  &  n_n535 ) ;
 assign n_n4470 = ( n_n518  &  wire13  &  n_n520 ) ;
 assign n_n4460 = ( n_n518  &  wire13  &  n_n530 ) ;
 assign n_n4473 = ( wire25  &  n_n455  &  n_n509 ) ;
 assign n_n4466 = ( n_n524  &  n_n518  &  wire13 ) ;
 assign n_n4895 = ( n_n491  &  wire11  &  n_n260 ) ;
 assign n_n4890 = ( n_n491  &  n_n532  &  wire17 ) ;
 assign wire260 = ( i_9_  &  n_n260  &  n_n520  &  n_n500 ) | ( (~ i_9_)  &  n_n260  &  n_n520  &  n_n500 ) ;
 assign wire16331 = ( n_n4888 ) | ( n_n4885 ) | ( wire260 ) ;
 assign n_n4850 = ( n_n524  &  n_n518  &  wire17 ) ;
 assign wire277 = ( i_9_  &  n_n522  &  n_n518  &  n_n260 ) | ( (~ i_9_)  &  n_n522  &  n_n518  &  n_n260 ) ;
 assign wire295 = ( n_n522  &  n_n509  &  wire17 ) | ( n_n524  &  n_n509  &  wire17 ) ;
 assign wire16334 = ( n_n4862 ) | ( n_n4850 ) | ( n_n4861 ) ;
 assign n_n2228 = ( wire277 ) | ( wire295 ) | ( wire16334 ) | ( _29100 ) ;
 assign n_n4881 = ( wire22  &  n_n260  &  n_n500 ) ;
 assign n_n4878 = ( n_n528  &  wire17  &  n_n500 ) ;
 assign n_n4880 = ( n_n526  &  wire17  &  n_n500 ) ;
 assign n_n4869 = ( n_n509  &  n_n260  &  wire20 ) ;
 assign n_n4877 = ( wire15  &  n_n260  &  n_n500 ) ;
 assign wire174 = ( wire25  &  n_n260  &  n_n500 ) | ( wire24  &  n_n260  &  n_n500 ) ;
 assign wire16342 = ( n_n4880 ) | ( n_n4869 ) | ( wire16339 ) | ( wire16340 ) ;
 assign n_n2178 = ( wire16331 ) | ( n_n2228 ) | ( wire16342 ) | ( _29098 ) ;
 assign n_n5321 = ( wire25  &  n_n65  &  n_n464 ) ;
 assign n_n5323 = ( n_n65  &  n_n464  &  wire24 ) ;
 assign n_n5324 = ( wire19  &  n_n464  &  n_n530 ) ;
 assign n_n5322 = ( wire19  &  n_n464  &  n_n532 ) ;
 assign n_n2274 = ( n_n5323 ) | ( n_n5324 ) | ( n_n5322 ) ;
 assign n_n5307 = ( n_n473  &  n_n65  &  wire24 ) ;
 assign n_n5326 = ( wire19  &  n_n464  &  n_n528 ) ;
 assign n_n5325 = ( n_n65  &  wire15  &  n_n464 ) ;
 assign n_n5332 = ( wire19  &  n_n522  &  n_n464 ) ;
 assign n_n5329 = ( n_n65  &  wire22  &  n_n464 ) ;
 assign wire115 = ( i_9_  &  n_n473  &  n_n65  &  n_n522 ) | ( (~ i_9_)  &  n_n473  &  n_n65  &  n_n522 ) ;
 assign wire16291 = ( i_9_  &  n_n473  &  n_n65  &  n_n524 ) | ( (~ i_9_)  &  n_n473  &  n_n65  &  n_n524 ) ;
 assign wire117 = ( wire459 ) | ( wire115 ) | ( wire16291 ) ;
 assign wire269 = ( i_9_  &  n_n473  &  n_n65  &  n_n528 ) | ( (~ i_9_)  &  n_n473  &  n_n65  &  n_n528 ) ;
 assign n_n2230 = ( wire388 ) | ( wire16351 ) | ( wire16352 ) ;
 assign n_n2229 = ( n_n4843 ) | ( n_n4846 ) | ( wire16355 ) | ( wire16356 ) ;
 assign wire16362 = ( n_n4824 ) | ( n_n4822 ) | ( n_n4823 ) | ( n_n4806 ) ;
 assign wire16363 = ( n_n4810 ) | ( wire186 ) | ( wire16360 ) ;
 assign n_n2179 = ( n_n2230 ) | ( n_n2229 ) | ( wire16362 ) | ( wire16363 ) ;
 assign n_n4776 = ( n_n482  &  n_n534  &  wire14 ) ;
 assign n_n4774 = ( n_n491  &  wire14  &  n_n520 ) ;
 assign n_n4786 = ( n_n482  &  n_n524  &  wire14 ) ;
 assign wire131 = ( n_n482  &  wire22  &  n_n325 ) | ( n_n482  &  wire21  &  n_n325 ) ;
 assign wire313 = ( i_9_  &  n_n482  &  n_n522  &  n_n325 ) | ( (~ i_9_)  &  n_n482  &  n_n522  &  n_n325 ) ;
 assign wire16374 = ( n_n4779 ) | ( n_n4790 ) | ( wire313 ) | ( wire16373 ) ;
 assign wire16375 = ( wire16349 ) | ( wire16350 ) | ( wire16367 ) | ( wire16368 ) ;
 assign n_n2162 = ( n_n2178 ) | ( n_n2179 ) | ( wire16374 ) | ( wire16375 ) ;
 assign n_n4755 = ( wire21  &  n_n325  &  n_n500 ) ;
 assign n_n4759 = ( n_n325  &  wire23  &  n_n500 ) ;
 assign n_n4760 = ( n_n491  &  n_n534  &  wire14 ) ;
 assign n_n4758 = ( wire14  &  n_n520  &  n_n500 ) ;
 assign n_n2238 = ( n_n4724 ) | ( n_n4727 ) | ( wire16388 ) | ( wire16389 ) ;
 assign wire16394 = ( n_n4695 ) | ( n_n4696 ) | ( wire173 ) ;
 assign wire16395 = ( n_n4711 ) | ( n_n4712 ) | ( wire442 ) ;
 assign wire16399 = ( n_n4717 ) | ( n_n2378 ) | ( wire16396 ) | ( _25663 ) ;
 assign n_n2182 = ( n_n2238 ) | ( wire16394 ) | ( wire16395 ) | ( wire16399 ) ;
 assign n_n2242 = ( n_n4677 ) | ( n_n4678 ) | ( wire16404 ) | ( wire16405 ) ;
 assign wire16410 = ( wire431 ) | ( n_n482  &  wire22  &  n_n390 ) ;
 assign wire16411 = ( n_n4662 ) | ( n_n4683 ) | ( wire16408 ) ;
 assign wire16415 = ( n_n3849 ) | ( n_n4693 ) | ( wire12422 ) | ( wire16412 ) ;
 assign n_n2183 = ( n_n2242 ) | ( wire16410 ) | ( wire16411 ) | ( wire16415 ) ;
 assign wire16423 = ( n_n4759 ) | ( n_n4760 ) | ( wire16420 ) | ( wire16421 ) ;
 assign wire16424 = ( wire16382 ) | ( wire16383 ) | ( wire16385 ) | ( wire16386 ) ;
 assign n_n2163 = ( n_n2182 ) | ( n_n2183 ) | ( wire16423 ) | ( wire16424 ) ;
 assign n_n4963 = ( wire21  &  n_n535  &  n_n195 ) ;
 assign n_n4959 = ( wire11  &  n_n535  &  n_n195 ) ;
 assign n_n4960 = ( n_n526  &  n_n535  &  wire18 ) ;
 assign n_n4964 = ( n_n522  &  n_n535  &  wire18 ) ;
 assign n_n2223 = ( wire31 ) | ( wire249 ) | ( _38 ) | ( _29196 ) ;
 assign wire16449 = ( n_n4900 ) | ( n_n4899 ) | ( wire16447 ) ;
 assign wire16450 = ( n_n4898 ) | ( n_n4897 ) | ( n_n4896 ) | ( wire16448 ) ;
 assign wire16456 = ( n_n4921 ) | ( n_n4919 ) | ( wire16453 ) | ( wire16454 ) ;
 assign n_n2177 = ( n_n2223 ) | ( wire16449 ) | ( wire16450 ) | ( wire16456 ) ;
 assign wire250 = ( n_n528  &  n_n535  &  wire18 ) | ( n_n535  &  wire18  &  n_n530 ) ;
 assign n_n4817 = ( wire22  &  n_n464  &  n_n325 ) ;
 assign n_n4827 = ( wire24  &  n_n535  &  n_n260 ) ;
 assign n_n4816 = ( n_n526  &  n_n464  &  wire14 ) ;
 assign n_n5097 = ( wire25  &  n_n518  &  n_n130 ) ;
 assign n_n5019 = ( n_n491  &  wire24  &  n_n195 ) ;
 assign n_n4416 = ( n_n473  &  n_n526  &  wire16 ) ;
 assign n_n4523 = ( n_n482  &  n_n455  &  wire24 ) ;
 assign n_n4547 = ( n_n473  &  wire21  &  n_n455 ) ;
 assign n_n4539 = ( n_n473  &  n_n455  &  wire24 ) ;
 assign n_n4521 = ( wire25  &  n_n482  &  n_n455 ) ;
 assign n_n4544 = ( n_n473  &  n_n526  &  wire13 ) ;
 assign n_n4557 = ( wire15  &  n_n464  &  n_n455 ) ;
 assign n_n4560 = ( n_n526  &  n_n464  &  wire13 ) ;
 assign n_n4553 = ( wire25  &  n_n464  &  n_n455 ) ;
 assign n_n4800 = ( n_n473  &  n_n526  &  wire14 ) ;
 assign n_n4777 = ( wire25  &  n_n482  &  n_n325 ) ;
 assign n_n4778 = ( n_n482  &  n_n532  &  wire14 ) ;
 assign n_n4780 = ( n_n482  &  wire14  &  n_n530 ) ;
 assign n_n2130 = ( n_n4777 ) | ( n_n4778 ) | ( n_n4780 ) ;
 assign n_n4803 = ( n_n473  &  wire21  &  n_n325 ) ;
 assign n_n4783 = ( n_n482  &  wire11  &  n_n325 ) ;
 assign n_n4812 = ( n_n464  &  wire14  &  n_n530 ) ;
 assign n_n4811 = ( n_n464  &  wire24  &  n_n325 ) ;
 assign n_n4781 = ( wire15  &  n_n482  &  n_n325 ) ;
 assign n_n4674 = ( n_n473  &  n_n524  &  wire10 ) ;
 assign n_n4661 = ( n_n482  &  n_n390  &  wire20 ) ;
 assign wire16508 = ( n_n4671 ) | ( n_n4672 ) | ( n_n4685 ) ;
 assign wire16509 = ( n_n4647 ) | ( n_n4656 ) | ( wire16506 ) ;
 assign n_n4361 = ( wire25  &  n_n536  &  n_n500 ) ;
 assign n_n4363 = ( n_n536  &  wire24  &  n_n500 ) ;
 assign n_n4359 = ( n_n536  &  n_n509  &  wire23 ) ;
 assign n_n4438 = ( n_n464  &  wire16  &  n_n520 ) ;
 assign n_n4439 = ( n_n464  &  n_n536  &  wire23 ) ;
 assign n_n4437 = ( n_n464  &  n_n536  &  wire20 ) ;
 assign n_n4825 = ( wire25  &  n_n535  &  n_n260 ) ;
 assign n_n4828 = ( wire17  &  n_n535  &  n_n530 ) ;
 assign n_n4824 = ( n_n534  &  wire17  &  n_n535 ) ;
 assign n_n4879 = ( wire11  &  n_n260  &  n_n500 ) ;
 assign n_n4937 = ( wire25  &  n_n464  &  n_n260 ) ;
 assign n_n4938 = ( n_n464  &  n_n532  &  wire17 ) ;
 assign n_n4936 = ( n_n464  &  n_n534  &  wire17 ) ;
 assign n_n5037 = ( wire15  &  n_n482  &  n_n195 ) ;
 assign n_n1570 = ( n_n5038 ) | ( n_n5035 ) | ( n_n5037 ) ;
 assign n_n5043 = ( n_n482  &  wire21  &  n_n195 ) ;
 assign n_n5045 = ( n_n482  &  n_n195  &  wire20 ) ;
 assign n_n5302 = ( n_n482  &  wire19  &  n_n520 ) ;
 assign n_n5294 = ( n_n482  &  wire19  &  n_n528 ) ;
 assign n_n4894 = ( n_n491  &  n_n528  &  wire17 ) ;
 assign n_n4916 = ( n_n482  &  n_n522  &  wire17 ) ;
 assign n_n4930 = ( n_n473  &  n_n524  &  wire17 ) ;
 assign n_n4947 = ( n_n464  &  wire21  &  n_n260 ) ;
 assign wire96 = ( n_n522  &  n_n491  &  wire17 ) | ( n_n491  &  wire17  &  n_n520 ) ;
 assign n_n5131 = ( wire24  &  n_n130  &  n_n500 ) ;
 assign n_n5137 = ( wire22  &  n_n130  &  n_n500 ) ;
 assign n_n5136 = ( n_n526  &  wire12  &  n_n500 ) ;
 assign n_n5200 = ( n_n526  &  n_n464  &  wire12 ) ;
 assign n_n5206 = ( n_n464  &  n_n520  &  wire12 ) ;
 assign n_n5146 = ( n_n491  &  n_n532  &  wire12 ) ;
 assign n_n5204 = ( n_n522  &  n_n464  &  wire12 ) ;
 assign n_n5191 = ( n_n473  &  n_n130  &  wire23 ) ;
 assign n_n5113 = ( wire25  &  n_n509  &  n_n130 ) ;
 assign n_n5081 = ( wire25  &  n_n535  &  n_n130 ) ;
 assign n_n5089 = ( wire22  &  n_n535  &  n_n130 ) ;
 assign n_n5124 = ( n_n522  &  n_n509  &  wire12 ) ;
 assign wire335 = ( n_n532  &  n_n509  &  wire12 ) | ( n_n509  &  wire12  &  n_n530 ) ;
 assign n_n5258 = ( wire19  &  n_n532  &  n_n500 ) ;
 assign n_n5274 = ( wire19  &  n_n491  &  n_n532 ) ;
 assign n_n5232 = ( wire19  &  n_n526  &  n_n518 ) ;
 assign n_n5255 = ( n_n65  &  n_n509  &  wire23 ) ;
 assign n_n5267 = ( n_n65  &  wire21  &  n_n500 ) ;
 assign n_n5222 = ( wire19  &  n_n535  &  n_n520 ) ;
 assign n_n5212 = ( wire19  &  n_n535  &  n_n530 ) ;
 assign n_n4344 = ( wire16  &  n_n534  &  n_n509 ) ;
 assign n_n4345 = ( wire25  &  n_n536  &  n_n509 ) ;
 assign n_n4343 = ( n_n518  &  n_n536  &  wire23 ) ;
 assign n_n4392 = ( n_n482  &  wire16  &  n_n534 ) ;
 assign n_n4393 = ( wire25  &  n_n482  &  n_n536 ) ;
 assign n_n4612 = ( n_n522  &  wire10  &  n_n509 ) ;
 assign n_n4611 = ( wire21  &  n_n390  &  n_n509 ) ;
 assign n_n4669 = ( n_n473  &  wire15  &  n_n390 ) ;
 assign n_n4673 = ( n_n473  &  wire22  &  n_n390 ) ;
 assign n_n4668 = ( n_n473  &  wire10  &  n_n530 ) ;
 assign n_n4734 = ( n_n509  &  wire14  &  n_n528 ) ;
 assign n_n4733 = ( wire15  &  n_n509  &  n_n325 ) ;
 assign n_n4792 = ( n_n473  &  n_n534  &  wire14 ) ;
 assign n_n4854 = ( n_n518  &  wire17  &  n_n520 ) ;
 assign n_n4855 = ( n_n518  &  n_n260  &  wire23 ) ;
 assign n_n4912 = ( n_n482  &  n_n526  &  wire17 ) ;
 assign n_n4908 = ( n_n482  &  wire17  &  n_n530 ) ;
 assign n_n4966 = ( n_n535  &  n_n520  &  wire18 ) ;
 assign n_n4968 = ( n_n518  &  n_n534  &  wire18 ) ;
 assign n_n5014 = ( n_n520  &  wire18  &  n_n500 ) ;
 assign n_n5015 = ( n_n195  &  wire23  &  n_n500 ) ;
 assign n_n5012 = ( n_n522  &  wire18  &  n_n500 ) ;
 assign n_n5067 = ( n_n464  &  wire24  &  n_n195 ) ;
 assign n_n5069 = ( wire15  &  n_n464  &  n_n195 ) ;
 assign n_n5066 = ( n_n464  &  n_n532  &  wire18 ) ;
 assign n_n5241 = ( wire25  &  n_n65  &  n_n509 ) ;
 assign n_n5243 = ( n_n65  &  wire24  &  n_n509 ) ;
 assign n_n5300 = ( n_n482  &  wire19  &  n_n522 ) ;
 assign n_n5299 = ( n_n65  &  n_n482  &  wire21 ) ;
 assign n_n4364 = ( wire16  &  n_n500  &  n_n530 ) ;
 assign n_n3533 = ( n_n4362 ) | ( n_n4363 ) | ( n_n4364 ) ;
 assign n_n4366 = ( wire16  &  n_n528  &  n_n500 ) ;
 assign n_n4365 = ( wire15  &  n_n536  &  n_n500 ) ;
 assign wire11607 = ( i_9_  &  n_n536  &  n_n528  &  n_n500 ) | ( (~ i_9_)  &  n_n536  &  n_n528  &  n_n500 ) ;
 assign n_n1308 = ( wire11607 ) | ( wire15  &  n_n536  &  n_n500 ) ;
 assign n_n4770 = ( n_n491  &  n_n524  &  wire14 ) ;
 assign n_n4769 = ( n_n491  &  wire22  &  n_n325 ) ;
 assign n_n4767 = ( n_n491  &  wire11  &  n_n325 ) ;
 assign n_n4764 = ( n_n491  &  wire14  &  n_n530 ) ;
 assign n_n4905 = ( wire25  &  n_n482  &  n_n260 ) ;
 assign wire352 = ( n_n482  &  n_n532  &  wire17 ) | ( n_n482  &  n_n534  &  wire17 ) ;
 assign n_n5046 = ( n_n482  &  n_n520  &  wire18 ) ;
 assign n_n5056 = ( n_n473  &  n_n526  &  wire18 ) ;
 assign n_n5057 = ( n_n473  &  wire22  &  n_n195 ) ;
 assign wire166 = ( i_9_  &  n_n473  &  n_n195  &  n_n530 ) | ( (~ i_9_)  &  n_n473  &  n_n195  &  n_n530 ) ;
 assign wire292 = ( i_9_  &  n_n482  &  n_n325  &  n_n520 ) | ( (~ i_9_)  &  n_n482  &  n_n325  &  n_n520 ) ;
 assign n_n4843 = ( n_n518  &  wire24  &  n_n260 ) ;
 assign n_n4845 = ( wire15  &  n_n518  &  n_n260 ) ;
 assign n_n4846 = ( n_n518  &  n_n528  &  wire17 ) ;
 assign n_n4848 = ( n_n526  &  n_n518  &  wire17 ) ;
 assign n_n4839 = ( n_n535  &  n_n260  &  wire23 ) ;
 assign n_n4840 = ( n_n518  &  n_n534  &  wire17 ) ;
 assign n_n4838 = ( wire17  &  n_n535  &  n_n520 ) ;
 assign n_n3820 = ( n_n4839 ) | ( n_n4840 ) | ( n_n4838 ) ;
 assign n_n4384 = ( n_n526  &  n_n491  &  wire16 ) ;
 assign n_n4390 = ( n_n491  &  wire16  &  n_n520 ) ;
 assign n_n4638 = ( n_n491  &  wire10  &  n_n528 ) ;
 assign n_n4633 = ( wire25  &  n_n491  &  n_n390 ) ;
 assign n_n5155 = ( n_n491  &  wire21  &  n_n130 ) ;
 assign n_n5161 = ( wire25  &  n_n482  &  n_n130 ) ;
 assign n_n4425 = ( wire25  &  n_n464  &  n_n536 ) ;
 assign n_n4482 = ( n_n524  &  wire13  &  n_n509 ) ;
 assign n_n4489 = ( wire25  &  n_n455  &  n_n500 ) ;
 assign n_n4504 = ( n_n491  &  wire13  &  n_n534 ) ;
 assign n_n4511 = ( n_n491  &  n_n455  &  wire11 ) ;
 assign n_n4526 = ( n_n482  &  wire13  &  n_n528 ) ;
 assign n_n4533 = ( n_n482  &  n_n455  &  wire20 ) ;
 assign n_n4554 = ( n_n464  &  wire13  &  n_n532 ) ;
 assign n_n4561 = ( wire22  &  n_n464  &  n_n455 ) ;
 assign n_n4568 = ( wire10  &  n_n534  &  n_n535 ) ;
 assign n_n4575 = ( wire11  &  n_n390  &  n_n535 ) ;
 assign n_n4590 = ( n_n518  &  wire10  &  n_n528 ) ;
 assign n_n4640 = ( n_n526  &  n_n491  &  wire10 ) ;
 assign n_n4647 = ( n_n491  &  n_n390  &  wire23 ) ;
 assign n_n4662 = ( n_n482  &  wire10  &  n_n520 ) ;
 assign n_n4690 = ( n_n524  &  n_n464  &  wire10 ) ;
 assign n_n4704 = ( n_n526  &  wire14  &  n_n535 ) ;
 assign n_n4711 = ( n_n325  &  n_n535  &  wire23 ) ;
 assign n_n4748 = ( wire14  &  n_n500  &  n_n530 ) ;
 assign n_n4821 = ( n_n464  &  n_n325  &  wire20 ) ;
 assign n_n4901 = ( n_n491  &  n_n260  &  wire20 ) ;
 assign n_n4974 = ( n_n518  &  n_n528  &  wire18 ) ;
 assign n_n5003 = ( wire24  &  n_n195  &  n_n500 ) ;
 assign n_n5047 = ( n_n482  &  n_n195  &  wire23 ) ;
 assign n_n5098 = ( n_n518  &  n_n532  &  wire12 ) ;
 assign n_n5105 = ( wire22  &  n_n518  &  n_n130 ) ;
 assign n_n5120 = ( n_n526  &  n_n509  &  wire12 ) ;
 assign n_n5127 = ( n_n509  &  n_n130  &  wire23 ) ;
 assign n_n5186 = ( n_n473  &  n_n524  &  wire12 ) ;
 assign n_n5193 = ( wire25  &  n_n464  &  n_n130 ) ;
 assign n_n5251 = ( n_n65  &  wire21  &  n_n509 ) ;
 assign n_n5266 = ( wire19  &  n_n524  &  n_n500 ) ;
 assign n_n5273 = ( wire25  &  n_n65  &  n_n491 ) ;
 assign n_n4347 = ( n_n536  &  wire24  &  n_n509 ) ;
 assign n_n4397 = ( wire15  &  n_n482  &  n_n536 ) ;
 assign n_n4398 = ( n_n482  &  wire16  &  n_n528 ) ;
 assign n_n4396 = ( n_n482  &  wire16  &  n_n530 ) ;
 assign n_n4524 = ( n_n482  &  wire13  &  n_n530 ) ;
 assign n_n4522 = ( n_n482  &  wire13  &  n_n532 ) ;
 assign wire170 = ( i_9_  &  n_n482  &  n_n455  &  n_n532 ) | ( (~ i_9_)  &  n_n482  &  n_n455  &  n_n532 ) ;
 assign n_n4246 = ( wire170 ) | ( n_n482  &  wire13  &  n_n530 ) ;
 assign n_n4670 = ( n_n473  &  wire10  &  n_n528 ) ;
 assign n_n4732 = ( n_n509  &  wire14  &  n_n530 ) ;
 assign n_n4789 = ( n_n482  &  n_n325  &  wire20 ) ;
 assign n_n4906 = ( n_n482  &  n_n532  &  wire17 ) ;
 assign n_n4967 = ( n_n535  &  n_n195  &  wire23 ) ;
 assign n_n5086 = ( n_n528  &  n_n535  &  wire12 ) ;
 assign n_n5087 = ( wire11  &  n_n535  &  n_n130 ) ;
 assign n_n4589 = ( wire15  &  n_n518  &  n_n390 ) ;
 assign n_n4587 = ( n_n518  &  wire24  &  n_n390 ) ;
 assign n_n881 = ( n_n4590 ) | ( n_n4589 ) | ( n_n4587 ) ;
 assign n_n4594 = ( n_n524  &  n_n518  &  wire10 ) ;
 assign n_n4083 = ( n_n881 ) | ( _25250 ) | ( _25251 ) | ( _25252 ) ;
 assign n_n4639 = ( n_n491  &  wire11  &  n_n390 ) ;
 assign n_n4904 = ( n_n482  &  n_n534  &  wire17 ) ;
 assign n_n4319 = ( n_n536  &  wire11  &  n_n535 ) ;
 assign n_n4320 = ( n_n526  &  wire16  &  n_n535 ) ;
 assign n_n4451 = ( wire21  &  n_n455  &  n_n535 ) ;
 assign n_n4918 = ( n_n482  &  wire17  &  n_n520 ) ;
 assign n_n4919 = ( n_n482  &  n_n260  &  wire23 ) ;
 assign n_n4917 = ( n_n482  &  n_n260  &  wire20 ) ;
 assign n_n4985 = ( wire25  &  n_n509  &  n_n195 ) ;
 assign n_n4984 = ( n_n534  &  n_n509  &  wire18 ) ;
 assign n_n5031 = ( n_n491  &  n_n195  &  wire23 ) ;
 assign n_n5114 = ( n_n532  &  n_n509  &  wire12 ) ;
 assign n_n5116 = ( n_n509  &  wire12  &  n_n530 ) ;
 assign n_n5162 = ( n_n482  &  n_n532  &  wire12 ) ;
 assign n_n4582 = ( wire10  &  n_n535  &  n_n520 ) ;
 assign n_n4584 = ( n_n518  &  wire10  &  n_n534 ) ;
 assign n_n4586 = ( n_n518  &  wire10  &  n_n532 ) ;
 assign wire365 = ( i_9_  &  n_n518  &  n_n390  &  n_n530 ) | ( (~ i_9_)  &  n_n518  &  n_n390  &  n_n530 ) ;
 assign wire14091 = ( n_n4586 ) | ( n_n4591 ) | ( n_n4592 ) ;
 assign wire14092 = ( n_n4590 ) | ( n_n4587 ) | ( wire365 ) ;
 assign n_n3348 = ( n_n4582 ) | ( n_n4584 ) | ( wire14091 ) | ( wire14092 ) ;
 assign n_n4876 = ( wire17  &  n_n500  &  n_n530 ) ;
 assign n_n4870 = ( n_n509  &  wire17  &  n_n520 ) ;
 assign n_n4871 = ( n_n509  &  n_n260  &  wire23 ) ;
 assign n_n4872 = ( n_n534  &  wire17  &  n_n500 ) ;
 assign wire461 = ( n_n4870 ) | ( n_n4871 ) | ( n_n4872 ) ;
 assign wire13850 = ( n_n4881 ) | ( n_n4878 ) | ( n_n4880 ) | ( n_n4877 ) ;
 assign n_n3326 = ( n_n4879 ) | ( n_n4876 ) | ( wire461 ) | ( wire13850 ) ;
 assign n_n5327 = ( n_n65  &  n_n464  &  wire11 ) ;
 assign n_n2643 = ( n_n5326 ) | ( n_n5325 ) | ( n_n5327 ) ;
 assign n_n4577 = ( wire22  &  n_n390  &  n_n535 ) ;
 assign n_n4576 = ( n_n526  &  wire10  &  n_n535 ) ;
 assign n_n4569 = ( wire25  &  n_n390  &  n_n535 ) ;
 assign n_n4574 = ( wire10  &  n_n528  &  n_n535 ) ;
 assign n_n4581 = ( n_n390  &  n_n535  &  wire20 ) ;
 assign n_n4572 = ( wire10  &  n_n535  &  n_n530 ) ;
 assign n_n4573 = ( wire15  &  n_n390  &  n_n535 ) ;
 assign n_n4579 = ( wire21  &  n_n390  &  n_n535 ) ;
 assign wire14087 = ( n_n4597 ) | ( n_n4598 ) | ( n_n4595 ) | ( n_n4596 ) ;
 assign wire14088 = ( n_n4602 ) | ( n_n4593 ) | ( n_n4601 ) | ( wire108 ) ;
 assign wire14101 = ( n_n4579 ) | ( wire14094 ) | ( wire14097 ) | ( wire14099 ) ;
 assign n_n3282 = ( n_n3348 ) | ( wire14087 ) | ( wire14088 ) | ( wire14101 ) ;
 assign n_n4538 = ( n_n473  &  wire13  &  n_n532 ) ;
 assign n_n4525 = ( wire15  &  n_n482  &  n_n455 ) ;
 assign n_n4531 = ( n_n482  &  wire21  &  n_n455 ) ;
 assign n_n4551 = ( n_n473  &  n_n455  &  wire23 ) ;
 assign n_n4552 = ( n_n464  &  wire13  &  n_n534 ) ;
 assign n_n3871 = ( n_n4553 ) | ( n_n4551 ) | ( n_n4552 ) ;
 assign wire212 = ( i_9_  &  n_n473  &  n_n522  &  n_n455 ) | ( (~ i_9_)  &  n_n473  &  n_n522  &  n_n455 ) ;
 assign n_n4550 = ( n_n473  &  wire13  &  n_n520 ) ;
 assign n_n4543 = ( n_n473  &  n_n455  &  wire11 ) ;
 assign wire14107 = ( i_9_  &  n_n473  &  n_n524  &  n_n455 ) | ( (~ i_9_)  &  n_n473  &  n_n524  &  n_n455 ) ;
 assign wire202 = ( wire212 ) | ( n_n4550 ) | ( n_n4543 ) | ( wire14107 ) ;
 assign wire14115 = ( wire202 ) | ( n_n4542 ) | ( wire201 ) | ( wire14111 ) ;
 assign wire14116 = ( n_n3871 ) | ( wire14105 ) | ( wire14106 ) | ( wire14112 ) ;
 assign n_n3260 = ( n_n3281 ) | ( n_n3282 ) | ( wire14115 ) | ( wire14116 ) ;
 assign n_n4629 = ( n_n390  &  wire20  &  n_n500 ) ;
 assign n_n4583 = ( n_n390  &  n_n535  &  wire23 ) ;
 assign n_n4842 = ( n_n518  &  n_n532  &  wire17 ) ;
 assign n_n4844 = ( n_n518  &  wire17  &  n_n530 ) ;
 assign n_n5303 = ( n_n65  &  n_n482  &  wire23 ) ;
 assign n_n5182 = ( n_n473  &  n_n528  &  wire12 ) ;
 assign n_n5173 = ( n_n482  &  wire20  &  n_n130 ) ;
 assign n_n5165 = ( wire15  &  n_n482  &  n_n130 ) ;
 assign n_n5230 = ( wire19  &  n_n518  &  n_n528 ) ;
 assign n_n5166 = ( n_n482  &  n_n528  &  wire12 ) ;
 assign n_n5163 = ( n_n482  &  wire24  &  n_n130 ) ;
 assign n_n5214 = ( wire19  &  n_n528  &  n_n535 ) ;
 assign n_n5002 = ( n_n532  &  wire18  &  n_n500 ) ;
 assign n_n5053 = ( n_n473  &  wire15  &  n_n195 ) ;
 assign n_n5033 = ( wire25  &  n_n482  &  n_n195 ) ;
 assign n_n5051 = ( n_n473  &  wire24  &  n_n195 ) ;
 assign n_n5006 = ( n_n528  &  wire18  &  n_n500 ) ;
 assign n_n4454 = ( wire13  &  n_n535  &  n_n520 ) ;
 assign n_n4518 = ( n_n491  &  wire13  &  n_n520 ) ;
 assign n_n4517 = ( n_n491  &  n_n455  &  wire20 ) ;
 assign wire664 = ( n_n491  &  n_n455  &  wire23 ) ;
 assign n_n3152 = ( n_n4518 ) | ( n_n4517 ) | ( wire664 ) ;
 assign n_n4725 = ( n_n518  &  n_n325  &  wire20 ) ;
 assign n_n4726 = ( n_n518  &  wire14  &  n_n520 ) ;
 assign n_n4861 = ( wire15  &  n_n509  &  n_n260 ) ;
 assign n_n5103 = ( n_n518  &  wire11  &  n_n130 ) ;
 assign n_n5104 = ( n_n526  &  n_n518  &  wire12 ) ;
 assign n_n5102 = ( n_n518  &  n_n528  &  wire12 ) ;
 assign n_n4395 = ( n_n482  &  n_n536  &  wire24 ) ;
 assign n_n4357 = ( n_n536  &  n_n509  &  wire20 ) ;
 assign wire15032 = ( n_n4355 ) | ( n_n4356 ) | ( n_n4358 ) ;
 assign wire15033 = ( n_n4359 ) | ( n_n4364 ) | ( _27356 ) ;
 assign n_n2638 = ( n_n4366 ) | ( n_n4357 ) | ( wire15032 ) | ( wire15033 ) ;
 assign wire425 = ( i_9_  &  n_n491  &  n_n524  &  n_n536 ) | ( (~ i_9_)  &  n_n491  &  n_n524  &  n_n536 ) ;
 assign wire15028 = ( n_n4379 ) | ( n_n4367 ) | ( n_n4380 ) | ( n_n4368 ) ;
 assign wire15029 = ( n_n4378 ) | ( n_n4374 ) | ( n_n4384 ) | ( wire423 ) ;
 assign n_n2560 = ( n_n2638 ) | ( wire15038 ) | ( _27368 ) | ( _27369 ) ;
 assign n_n4426 = ( n_n464  &  wire16  &  n_n532 ) ;
 assign n_n4409 = ( wire25  &  n_n473  &  n_n536 ) ;
 assign wire15048 = ( n_n4408 ) | ( n_n4405 ) | ( n_n4406 ) ;
 assign wire15049 = ( n_n4397 ) | ( n_n4398 ) | ( wire15046 ) ;
 assign n_n2635 = ( n_n4404 ) | ( n_n4409 ) | ( wire15048 ) | ( wire15049 ) ;
 assign wire37 = ( i_9_  &  n_n464  &  n_n536  &  n_n534 ) | ( (~ i_9_)  &  n_n464  &  n_n536  &  n_n534 ) ;
 assign wire15044 = ( n_n4411 ) | ( n_n4412 ) | ( wire15042 ) ;
 assign n_n2559 = ( n_n2635 ) | ( _27388 ) | ( _27389 ) | ( _27390 ) ;
 assign n_n4315 = ( n_n536  &  wire24  &  n_n535 ) ;
 assign n_n4360 = ( wire16  &  n_n534  &  n_n500 ) ;
 assign n_n4487 = ( n_n455  &  n_n509  &  wire23 ) ;
 assign n_n4483 = ( wire21  &  n_n455  &  n_n509 ) ;
 assign n_n4837 = ( n_n535  &  n_n260  &  wire20 ) ;
 assign n_n4899 = ( n_n491  &  wire21  &  n_n260 ) ;
 assign n_n4986 = ( n_n532  &  n_n509  &  wire18 ) ;
 assign n_n5044 = ( n_n482  &  n_n522  &  wire18 ) ;
 assign n_n5115 = ( wire24  &  n_n509  &  n_n130 ) ;
 assign n_n5175 = ( n_n482  &  n_n130  &  wire23 ) ;
 assign n_n5177 = ( wire25  &  n_n473  &  n_n130 ) ;
 assign n_n5311 = ( n_n473  &  n_n65  &  wire11 ) ;
 assign n_n4798 = ( n_n473  &  wire14  &  n_n528 ) ;
 assign n_n4804 = ( n_n473  &  n_n522  &  wire14 ) ;
 assign n_n4794 = ( n_n473  &  n_n532  &  wire14 ) ;
 assign n_n4795 = ( n_n473  &  wire24  &  n_n325 ) ;
 assign n_n4793 = ( wire25  &  n_n473  &  n_n325 ) ;
 assign n_n4796 = ( n_n473  &  wire14  &  n_n530 ) ;
 assign n_n4797 = ( n_n473  &  wire15  &  n_n325 ) ;
 assign n_n4801 = ( n_n473  &  wire22  &  n_n325 ) ;
 assign n_n4933 = ( n_n473  &  n_n260  &  wire20 ) ;
 assign n_n4935 = ( n_n473  &  n_n260  &  wire23 ) ;
 assign wire249 = ( n_n4927 ) | ( n_n4924 ) | ( n_n4926 ) | ( n_n4925 ) ;
 assign wire289 = ( wire15  &  n_n518  &  n_n130 ) | ( wire22  &  n_n518  &  n_n130 ) ;
 assign n_n4497 = ( wire22  &  n_n455  &  n_n500 ) ;
 assign wire65 = ( i_9_  &  n_n524  &  n_n455  &  n_n500 ) | ( (~ i_9_)  &  n_n524  &  n_n455  &  n_n500 ) ;
 assign wire66 = ( i_9_  &  n_n455  &  n_n528  &  n_n500 ) | ( (~ i_9_)  &  n_n455  &  n_n528  &  n_n500 ) ;
 assign n_n4478 = ( wire13  &  n_n509  &  n_n528 ) ;
 assign n_n4477 = ( wire15  &  n_n455  &  n_n509 ) ;
 assign n_n4475 = ( n_n455  &  wire24  &  n_n509 ) ;
 assign n_n4476 = ( wire13  &  n_n509  &  n_n530 ) ;
 assign wire70 = ( wire21  &  n_n455  &  n_n509 ) | ( n_n455  &  n_n509  &  wire20 ) ;
 assign wire184 = ( n_n526  &  wire13  &  n_n509 ) | ( n_n524  &  wire13  &  n_n509 ) ;
 assign wire16576 = ( wire70 ) | ( wire184 ) ;
 assign wire693 = ( wire15  &  n_n535  &  n_n260 ) ;
 assign wire388 = ( n_n4830 ) | ( n_n4831 ) | ( n_n4828 ) | ( wire693 ) ;
 assign wire16351 = ( i_9_  &  n_n524  &  n_n535  &  n_n260 ) | ( (~ i_9_)  &  n_n524  &  n_n535  &  n_n260 ) ;
 assign wire16352 = ( n_n4832 ) | ( n_n4825 ) | ( n_n4826 ) ;
 assign wire176 = ( i_9_  &  n_n518  &  n_n260  &  n_n530 ) | ( (~ i_9_)  &  n_n518  &  n_n260  &  n_n530 ) ;
 assign wire16355 = ( n_n4842 ) | ( n_n4837 ) | ( n_n4841 ) ;
 assign wire16356 = ( n_n4839 ) | ( n_n4840 ) | ( wire176 ) ;
 assign n_n4822 = ( n_n464  &  wire14  &  n_n520 ) ;
 assign n_n4823 = ( n_n464  &  n_n325  &  wire23 ) ;
 assign n_n4806 = ( n_n473  &  wire14  &  n_n520 ) ;
 assign n_n4820 = ( n_n522  &  n_n464  &  wire14 ) ;
 assign n_n4818 = ( n_n524  &  n_n464  &  wire14 ) ;
 assign n_n4810 = ( n_n464  &  n_n532  &  wire14 ) ;
 assign wire186 = ( n_n464  &  wire21  &  n_n325 ) | ( n_n464  &  n_n325  &  wire20 ) ;
 assign n_n4415 = ( n_n473  &  n_n536  &  wire11 ) ;
 assign wire16520 = ( n_n4414 ) | ( n_n4411 ) | ( n_n4412 ) ;
 assign wire16521 = ( n_n4409 ) | ( n_n4410 ) | ( wire16518 ) ;
 assign n_n2263 = ( n_n4408 ) | ( n_n4415 ) | ( wire16520 ) | ( wire16521 ) ;
 assign wire16527 = ( wire98 ) | ( n_n4430 ) | ( n_n4439 ) | ( n_n4428 ) ;
 assign n_n4326 = ( wire16  &  n_n535  &  n_n520 ) ;
 assign n_n2446 = ( n_n4327 ) | ( n_n4324 ) | ( n_n4326 ) ;
 assign n_n4336 = ( n_n526  &  wire16  &  n_n518 ) ;
 assign wire14473 = ( wire22  &  n_n518  &  n_n536 ) | ( n_n518  &  wire21  &  n_n536 ) ;
 assign n_n2443 = ( wire14473 ) | ( n_n522  &  wire16  &  n_n518 ) ;
 assign n_n4328 = ( wire16  &  n_n518  &  n_n534 ) ;
 assign n_n4330 = ( wire16  &  n_n518  &  n_n532 ) ;
 assign n_n2445 = ( n_n4331 ) | ( n_n4328 ) | ( n_n4330 ) ;
 assign wire171 = ( wire22  &  n_n536  &  n_n535 ) | ( n_n536  &  wire11  &  n_n535 ) ;
 assign wire198 = ( i_9_  &  n_n518  &  n_n536  &  n_n530 ) | ( (~ i_9_)  &  n_n518  &  n_n536  &  n_n530 ) ;
 assign wire283 = ( i_9_  &  n_n536  &  n_n532  &  n_n535 ) | ( (~ i_9_)  &  n_n536  &  n_n532  &  n_n535 ) ;
 assign n_n2435 = ( n_n4388 ) | ( n_n4391 ) | ( n_n4390 ) ;
 assign n_n4386 = ( n_n491  &  n_n524  &  wire16 ) ;
 assign wire12447 = ( i_9_  &  n_n526  &  n_n491  &  n_n536 ) | ( (~ i_9_)  &  n_n526  &  n_n491  &  n_n536 ) ;
 assign wire14460 = ( wire15  &  n_n491  &  n_n536 ) | ( n_n491  &  n_n536  &  wire11 ) ;
 assign wire54 = ( n_n4386 ) | ( wire12447 ) | ( wire14460 ) ;
 assign n_n4370 = ( n_n524  &  wire16  &  n_n500 ) ;
 assign n_n4368 = ( n_n526  &  wire16  &  n_n500 ) ;
 assign wire282 = ( n_n4369 ) | ( n_n4370 ) | ( n_n4368 ) ;
 assign wire423 = ( i_9_  &  n_n491  &  n_n536  &  n_n534 ) | ( (~ i_9_)  &  n_n491  &  n_n536  &  n_n534 ) ;
 assign n_n4503 = ( n_n455  &  wire23  &  n_n500 ) ;
 assign n_n4502 = ( wire13  &  n_n520  &  n_n500 ) ;
 assign n_n4500 = ( n_n522  &  wire13  &  n_n500 ) ;
 assign n_n4546 = ( n_n473  &  n_n524  &  wire13 ) ;
 assign n_n4555 = ( n_n464  &  n_n455  &  wire24 ) ;
 assign wire213 = ( i_9_  &  n_n464  &  n_n455  &  n_n528 ) | ( (~ i_9_)  &  n_n464  &  n_n455  &  n_n528 ) ;
 assign n_n4656 = ( n_n482  &  n_n526  &  wire10 ) ;
 assign n_n4659 = ( n_n482  &  wire21  &  n_n390 ) ;
 assign n_n5106 = ( n_n524  &  n_n518  &  wire12 ) ;
 assign n_n4341 = ( n_n518  &  n_n536  &  wire20 ) ;
 assign n_n5117 = ( wire15  &  n_n509  &  n_n130 ) ;
 assign n_n5223 = ( n_n65  &  n_n535  &  wire23 ) ;
 assign n_n5328 = ( wire19  &  n_n526  &  n_n464 ) ;
 assign n_n5254 = ( wire19  &  n_n509  &  n_n520 ) ;
 assign n_n5249 = ( n_n65  &  wire22  &  n_n509 ) ;
 assign n_n5233 = ( n_n65  &  wire22  &  n_n518 ) ;
 assign n_n5236 = ( wire19  &  n_n522  &  n_n518 ) ;
 assign n_n5262 = ( wire19  &  n_n528  &  n_n500 ) ;
 assign n_n5278 = ( wire19  &  n_n491  &  n_n528 ) ;
 assign wire449 = ( i_9_  &  n_n65  &  n_n526  &  n_n535 ) | ( (~ i_9_)  &  n_n65  &  n_n526  &  n_n535 ) ;
 assign wire16774 = ( _64 ) | ( wire19  &  n_n522  &  n_n518 ) ;
 assign wire16775 = ( n_n5278 ) | ( n_n5290 ) | ( n_n5289 ) ;
 assign wire16776 = ( n_n5206 ) | ( n_n5223 ) | ( wire449 ) ;
 assign wire16777 = ( n_n5328 ) | ( n_n5254 ) | ( wire16773 ) ;
 assign n_n2083 = ( wire16774 ) | ( wire16775 ) | ( wire16776 ) | ( wire16777 ) ;
 assign n_n4375 = ( n_n536  &  wire23  &  n_n500 ) ;
 assign n_n4833 = ( wire22  &  n_n535  &  n_n260 ) ;
 assign n_n4875 = ( wire24  &  n_n260  &  n_n500 ) ;
 assign n_n4940 = ( n_n464  &  wire17  &  n_n530 ) ;
 assign n_n4939 = ( n_n464  &  wire24  &  n_n260 ) ;
 assign n_n4729 = ( wire25  &  n_n509  &  n_n325 ) ;
 assign n_n4728 = ( n_n534  &  n_n509  &  wire14 ) ;
 assign wire373 = ( i_9_  &  n_n509  &  n_n325  &  n_n520 ) | ( (~ i_9_)  &  n_n509  &  n_n325  &  n_n520 ) ;
 assign wire374 = ( i_9_  &  n_n522  &  n_n509  &  n_n325 ) | ( (~ i_9_)  &  n_n522  &  n_n509  &  n_n325 ) ;
 assign n_n5132 = ( wire12  &  n_n500  &  n_n530 ) ;
 assign n_n5128 = ( n_n534  &  wire12  &  n_n500 ) ;
 assign n_n5016 = ( n_n491  &  n_n534  &  wire18 ) ;
 assign wire732 = ( n_n473  &  wire12  &  n_n530 ) ;
 assign n_n4129 = ( n_n5181 ) | ( n_n5182 ) | ( wire732 ) ;
 assign n_n5306 = ( n_n473  &  wire19  &  n_n532 ) ;
 assign n_n5308 = ( n_n473  &  wire19  &  n_n530 ) ;
 assign n_n3019 = ( n_n5307 ) | ( n_n5306 ) | ( n_n5308 ) ;
 assign n_n5009 = ( wire22  &  n_n195  &  n_n500 ) ;
 assign n_n5335 = ( n_n65  &  n_n464  &  wire23 ) ;
 assign n_n4562 = ( n_n524  &  n_n464  &  wire13 ) ;
 assign n_n4506 = ( n_n491  &  wire13  &  n_n532 ) ;
 assign n_n4492 = ( wire13  &  n_n500  &  n_n530 ) ;
 assign n_n4580 = ( n_n522  &  wire10  &  n_n535 ) ;
 assign n_n4635 = ( n_n491  &  wire24  &  n_n390 ) ;
 assign wire12047 = ( n_n4591 ) | ( n_n4592 ) | ( wire745 ) ;
 assign wire12048 = ( n_n4617 ) | ( n_n4618 ) | ( n_n4576 ) | ( n_n4569 ) ;
 assign n_n1338 = ( n_n4580 ) | ( n_n4635 ) | ( wire12047 ) | ( wire12048 ) ;
 assign n_n4496 = ( n_n526  &  wire13  &  n_n500 ) ;
 assign n_n4535 = ( n_n482  &  n_n455  &  wire23 ) ;
 assign wire12054 = ( n_n4458 ) | ( n_n4436 ) | ( wire70 ) | ( n_n4474 ) ;
 assign n_n1326 = ( n_n1338 ) | ( wire12060 ) | ( wire12061 ) | ( _23853 ) ;
 assign n_n4743 = ( n_n509  &  n_n325  &  wire23 ) ;
 assign wire12067 = ( n_n4764 ) | ( n_n4763 ) | ( n_n4751 ) ;
 assign wire12068 = ( n_n4737 ) | ( n_n4756 ) | ( n_n4724 ) | ( n_n4759 ) ;
 assign n_n1336 = ( n_n4732 ) | ( n_n4743 ) | ( wire12067 ) | ( wire12068 ) ;
 assign n_n4788 = ( n_n482  &  n_n522  &  wire14 ) ;
 assign wire12074 = ( n_n4666 ) | ( n_n4649 ) | ( n_n4638 ) | ( n_n4655 ) ;
 assign wire12075 = ( n_n4658 ) | ( n_n4708 ) | ( n_n4706 ) | ( wire366 ) ;
 assign wire12083 = ( n_n4823 ) | ( n_n4806 ) | ( wire12080 ) | ( wire12081 ) ;
 assign n_n1325 = ( n_n1336 ) | ( wire12074 ) | ( wire12075 ) | ( wire12083 ) ;
 assign n_n4342 = ( wire16  &  n_n518  &  n_n520 ) ;
 assign n_n4608 = ( n_n526  &  wire10  &  n_n509 ) ;
 assign n_n4610 = ( n_n524  &  wire10  &  n_n509 ) ;
 assign n_n4606 = ( wire10  &  n_n509  &  n_n528 ) ;
 assign n_n4675 = ( n_n473  &  wire21  &  n_n390 ) ;
 assign n_n4676 = ( n_n473  &  n_n522  &  wire10 ) ;
 assign n_n4730 = ( n_n532  &  n_n509  &  wire14 ) ;
 assign n_n4802 = ( n_n473  &  n_n524  &  wire14 ) ;
 assign n_n4851 = ( n_n518  &  wire21  &  n_n260 ) ;
 assign n_n4852 = ( n_n522  &  n_n518  &  wire17 ) ;
 assign n_n4914 = ( n_n482  &  n_n524  &  wire17 ) ;
 assign n_n4962 = ( n_n524  &  n_n535  &  wire18 ) ;
 assign n_n4956 = ( n_n535  &  wire18  &  n_n530 ) ;
 assign n_n5020 = ( n_n491  &  wire18  &  n_n530 ) ;
 assign n_n5064 = ( n_n464  &  n_n534  &  wire18 ) ;
 assign n_n5189 = ( n_n473  &  wire20  &  n_n130 ) ;
 assign n_n5190 = ( n_n473  &  n_n520  &  wire12 ) ;
 assign n_n5188 = ( n_n473  &  n_n522  &  wire12 ) ;
 assign n_n4352 = ( n_n526  &  wire16  &  n_n509 ) ;
 assign n_n4351 = ( n_n536  &  wire11  &  n_n509 ) ;
 assign n_n4356 = ( n_n522  &  wire16  &  n_n509 ) ;
 assign wire67 = ( i_9_  &  n_n536  &  n_n532  &  n_n509 ) | ( (~ i_9_)  &  n_n536  &  n_n532  &  n_n509 ) ;
 assign wire11610 = ( n_n4357 ) | ( n_n4356 ) | ( n_n4358 ) ;
 assign wire11611 = ( wire67 ) | ( n_n4353 ) | ( n_n4354 ) ;
 assign n_n1120 = ( n_n4352 ) | ( n_n4351 ) | ( wire11610 ) | ( wire11611 ) ;
 assign n_n4507 = ( n_n491  &  n_n455  &  wire24 ) ;
 assign n_n4509 = ( wire15  &  n_n491  &  n_n455 ) ;
 assign n_n4508 = ( n_n491  &  wire13  &  n_n530 ) ;
 assign wire129 = ( i_9_  &  n_n526  &  n_n491  &  n_n455 ) | ( (~ i_9_)  &  n_n526  &  n_n491  &  n_n455 ) ;
 assign wire308 = ( i_9_  &  n_n491  &  n_n455  &  n_n528 ) | ( (~ i_9_)  &  n_n491  &  n_n455  &  n_n528 ) ;
 assign n_n4622 = ( wire10  &  n_n528  &  n_n500 ) ;
 assign n_n4621 = ( wire15  &  n_n390  &  n_n500 ) ;
 assign wire75 = ( n_n526  &  wire10  &  n_n500 ) ;
 assign n_n3861 = ( n_n4622 ) | ( n_n4621 ) | ( wire75 ) ;
 assign n_n5073 = ( wire22  &  n_n464  &  n_n195 ) ;
 assign n_n5074 = ( n_n524  &  n_n464  &  wire18 ) ;
 assign n_n5072 = ( n_n526  &  n_n464  &  wire18 ) ;
 assign n_n4152 = ( n_n5073 ) | ( n_n5074 ) | ( n_n5072 ) ;
 assign n_n4931 = ( n_n473  &  wire21  &  n_n260 ) ;
 assign wire180 = ( i_9_  &  n_n473  &  n_n260  &  n_n520 ) | ( (~ i_9_)  &  n_n473  &  n_n260  &  n_n520 ) ;
 assign wire382 = ( i_9_  &  n_n473  &  n_n522  &  n_n260 ) | ( (~ i_9_)  &  n_n473  &  n_n522  &  n_n260 ) ;
 assign n_n4978 = ( n_n524  &  n_n518  &  wire18 ) ;
 assign n_n4980 = ( n_n522  &  n_n518  &  wire18 ) ;
 assign n_n4897 = ( n_n491  &  wire22  &  n_n260 ) ;
 assign n_n1985 = ( n_n4885 ) | ( n_n4884 ) | ( n_n4883 ) ;
 assign n_n3815 = ( n_n4876 ) | ( n_n4875 ) | ( n_n4874 ) ;
 assign wire11818 = ( n_n526  &  wire17  &  n_n500 ) | ( n_n524  &  wire17  &  n_n500 ) ;
 assign n_n1077 = ( n_n4877 ) | ( n_n1985 ) | ( n_n3815 ) | ( wire11818 ) ;
 assign wire264 = ( n_n491  &  n_n528  &  wire17 ) | ( n_n491  &  wire17  &  n_n530 ) ;
 assign n_n4349 = ( wire15  &  n_n536  &  n_n509 ) ;
 assign n_n4348 = ( wire16  &  n_n509  &  n_n530 ) ;
 assign n_n1002 = ( n_n4350 ) | ( n_n4349 ) | ( n_n4348 ) ;
 assign n_n5172 = ( n_n482  &  n_n522  &  wire12 ) ;
 assign n_n4419 = ( n_n473  &  wire21  &  n_n536 ) ;
 assign n_n4605 = ( wire15  &  n_n390  &  n_n509 ) ;
 assign n_n4655 = ( n_n482  &  wire11  &  n_n390 ) ;
 assign n_n4683 = ( n_n464  &  wire24  &  n_n390 ) ;
 assign n_n4689 = ( wire22  &  n_n464  &  n_n390 ) ;
 assign n_n4697 = ( wire25  &  n_n325  &  n_n535 ) ;
 assign n_n4703 = ( wire11  &  n_n325  &  n_n535 ) ;
 assign n_n4712 = ( n_n518  &  n_n534  &  wire14 ) ;
 assign n_n4763 = ( n_n491  &  wire24  &  n_n325 ) ;
 assign n_n4915 = ( n_n482  &  wire21  &  n_n260 ) ;
 assign n_n4989 = ( wire15  &  n_n509  &  n_n195 ) ;
 assign n_n5011 = ( wire21  &  n_n195  &  n_n500 ) ;
 assign n_n5061 = ( n_n473  &  n_n195  &  wire20 ) ;
 assign n_n5070 = ( n_n464  &  n_n528  &  wire18 ) ;
 assign n_n5076 = ( n_n522  &  n_n464  &  wire18 ) ;
 assign n_n5135 = ( wire11  &  n_n130  &  n_n500 ) ;
 assign n_n5157 = ( n_n491  &  wire20  &  n_n130 ) ;
 assign n_n5201 = ( wire22  &  n_n464  &  n_n130 ) ;
 assign n_n5207 = ( n_n464  &  n_n130  &  wire23 ) ;
 assign n_n5237 = ( n_n65  &  n_n518  &  wire20 ) ;
 assign n_n5252 = ( wire19  &  n_n522  &  n_n509 ) ;
 assign n_n4353 = ( wire22  &  n_n536  &  n_n509 ) ;
 assign n_n4456 = ( n_n518  &  wire13  &  n_n534 ) ;
 assign n_n4671 = ( n_n473  &  wire11  &  n_n390 ) ;
 assign n_n4747 = ( wire24  &  n_n325  &  n_n500 ) ;
 assign n_n4772 = ( n_n522  &  n_n491  &  wire14 ) ;
 assign n_n4773 = ( n_n491  &  n_n325  &  wire20 ) ;
 assign n_n4771 = ( n_n491  &  wire21  &  n_n325 ) ;
 assign wire12393 = ( i_9_  &  n_n522  &  n_n491  &  n_n325 ) | ( (~ i_9_)  &  n_n522  &  n_n491  &  n_n325 ) ;
 assign n_n5023 = ( n_n491  &  wire11  &  n_n195 ) ;
 assign n_n5024 = ( n_n526  &  n_n491  &  wire18 ) ;
 assign n_n5082 = ( n_n532  &  n_n535  &  wire12 ) ;
 assign n_n5084 = ( n_n535  &  wire12  &  n_n530 ) ;
 assign n_n5275 = ( n_n65  &  n_n491  &  wire24 ) ;
 assign n_n5276 = ( wire19  &  n_n491  &  n_n530 ) ;
 assign n_n4600 = ( wire10  &  n_n534  &  n_n509 ) ;
 assign wire45 = ( i_9_  &  n_n518  &  n_n390  &  n_n520 ) | ( (~ i_9_)  &  n_n518  &  n_n390  &  n_n520 ) ;
 assign n_n4775 = ( n_n491  &  n_n325  &  wire23 ) ;
 assign n_n4204 = ( n_n4776 ) | ( n_n4774 ) | ( n_n4775 ) ;
 assign n_n4065 = ( n_n4827 ) | ( n_n4824 ) | ( wire388 ) | ( wire13156 ) ;
 assign wire13162 = ( n_n4816 ) | ( n_n4806 ) | ( n_n4805 ) | ( n_n4815 ) ;
 assign wire13163 = ( n_n4817 ) | ( n_n4800 ) | ( n_n4803 ) | ( n_n4804 ) ;
 assign wire13166 = ( n_n4801 ) | ( n_n4818 ) | ( n_n4197 ) | ( wire390 ) ;
 assign wire13177 = ( n_n4839 ) | ( n_n4840 ) | ( n_n4838 ) ;
 assign wire13178 = ( n_n4834 ) | ( n_n4835 ) | ( n_n4832 ) | ( n_n4833 ) ;
 assign wire13181 = ( wire13171 ) | ( wire13174 ) | ( _25555 ) ;
 assign wire13228 = ( wire13215 ) | ( wire13216 ) | ( _25613 ) | ( _25616 ) ;
 assign wire13229 = ( n_n814 ) | ( wire13222 ) | ( wire13223 ) | ( wire13224 ) ;
 assign wire13233 = ( wire295 ) | ( wire174 ) | ( wire461 ) | ( _25630 ) ;
 assign wire13236 = ( n_n4058 ) | ( n_n4056 ) | ( wire13213 ) | ( wire13234 ) ;
 assign n_n3990 = ( wire13228 ) | ( wire13229 ) | ( wire13233 ) | ( wire13236 ) ;
 assign n_n4753 = ( wire22  &  n_n325  &  n_n500 ) ;
 assign n_n4752 = ( n_n526  &  wire14  &  n_n500 ) ;
 assign n_n4075 = ( n_n4694 ) | ( n_n4700 ) | ( n_n4219 ) | ( wire13244 ) ;
 assign wire13249 = ( n_n4710 ) | ( n_n4709 ) | ( n_n4705 ) | ( n_n4706 ) ;
 assign wire13250 = ( n_n4722 ) | ( n_n4721 ) | ( wire173 ) ;
 assign wire13254 = ( n_n4717 ) | ( wire13251 ) | ( _25663 ) | ( _25671 ) ;
 assign n_n4013 = ( n_n4075 ) | ( wire13249 ) | ( wire13250 ) | ( wire13254 ) ;
 assign wire47 = ( n_n532  &  wire14  &  n_n500 ) | ( n_n534  &  wire14  &  n_n500 ) ;
 assign wire13270 = ( wire13259 ) | ( wire13260 ) | ( wire13263 ) | ( wire13264 ) ;
 assign n_n3992 = ( n_n4013 ) | ( wire13277 ) | ( _25724 ) | ( _25725 ) ;
 assign n_n4457 = ( wire25  &  n_n518  &  n_n455 ) ;
 assign n_n5075 = ( n_n464  &  wire21  &  n_n195 ) ;
 assign n_n5079 = ( n_n464  &  n_n195  &  wire23 ) ;
 assign n_n5088 = ( n_n526  &  n_n535  &  wire12 ) ;
 assign n_n5078 = ( n_n464  &  n_n520  &  wire18 ) ;
 assign n_n5083 = ( wire24  &  n_n535  &  n_n130 ) ;
 assign wire123 = ( i_9_  &  n_n535  &  n_n130  &  n_n530 ) | ( (~ i_9_)  &  n_n535  &  n_n130  &  n_n530 ) ;
 assign wire122 = ( wire15  &  n_n518  &  n_n130 ) | ( n_n518  &  wire24  &  n_n130 ) ;
 assign wire232 = ( i_9_  &  n_n524  &  n_n535  &  n_n130 ) | ( (~ i_9_)  &  n_n524  &  n_n535  &  n_n130 ) ;
 assign n_n5063 = ( n_n473  &  n_n195  &  wire23 ) ;
 assign n_n5058 = ( n_n473  &  n_n524  &  wire18 ) ;
 assign wire160 = ( n_n464  &  n_n532  &  wire18 ) | ( n_n464  &  wire18  &  n_n530 ) ;
 assign n_n4891 = ( n_n491  &  wire24  &  n_n260 ) ;
 assign n_n4836 = ( n_n522  &  wire17  &  n_n535 ) ;
 assign wire14260 = ( n_n4883 ) | ( n_n4869 ) | ( n_n4870 ) ;
 assign wire14261 = ( n_n4895 ) | ( n_n4825 ) | ( n_n4879 ) | ( n_n4841 ) ;
 assign n_n3558 = ( n_n4891 ) | ( n_n4836 ) | ( wire14260 ) | ( wire14261 ) ;
 assign wire14267 = ( n_n4958 ) | ( n_n4921 ) | ( n_n4963 ) | ( n_n4916 ) ;
 assign wire14268 = ( wire352 ) | ( n_n4933 ) | ( n_n4948 ) | ( n_n4973 ) ;
 assign n_n3557 = ( wire14267 ) | ( wire14268 ) ;
 assign n_n3560 = ( n_n4708 ) | ( n_n4695 ) | ( wire14316 ) | ( wire14317 ) ;
 assign n_n3561 = ( n_n4660 ) | ( n_n4665 ) | ( wire14322 ) | ( wire14323 ) ;
 assign wire14332 = ( n_n4747 ) | ( n_n4752 ) | ( wire14329 ) | ( wire14330 ) ;
 assign n_n3548 = ( n_n3560 ) | ( n_n3561 ) | ( wire14332 ) ;
 assign n_n4505 = ( wire25  &  n_n491  &  n_n455 ) ;
 assign n_n5095 = ( n_n535  &  n_n130  &  wire23 ) ;
 assign n_n5158 = ( n_n491  &  n_n520  &  wire12 ) ;
 assign n_n5154 = ( n_n491  &  n_n524  &  wire12 ) ;
 assign n_n3469 = ( n_n4770 ) | ( n_n4773 ) | ( n_n4771 ) ;
 assign n_n5013 = ( n_n195  &  wire20  &  n_n500 ) ;
 assign n_n5150 = ( n_n491  &  n_n528  &  wire12 ) ;
 assign n_n5147 = ( n_n491  &  wire24  &  n_n130 ) ;
 assign wire76 = ( i_9_  &  n_n491  &  n_n130  &  n_n530 ) | ( (~ i_9_)  &  n_n491  &  n_n130  &  n_n530 ) ;
 assign wire196 = ( i_9_  &  n_n526  &  n_n491  &  n_n130 ) | ( (~ i_9_)  &  n_n526  &  n_n491  &  n_n130 ) ;
 assign wire57 = ( i_9_  &  n_n524  &  n_n518  &  n_n195 ) | ( (~ i_9_)  &  n_n524  &  n_n518  &  n_n195 ) ;
 assign wire251 = ( i_9_  &  n_n518  &  n_n520  &  n_n195 ) | ( (~ i_9_)  &  n_n518  &  n_n520  &  n_n195 ) ;
 assign n_n4948 = ( n_n522  &  n_n464  &  wire17 ) ;
 assign n_n4957 = ( wire15  &  n_n535  &  n_n195 ) ;
 assign n_n4971 = ( n_n518  &  wire24  &  n_n195 ) ;
 assign wire342 = ( i_9_  &  n_n524  &  n_n535  &  n_n195 ) | ( (~ i_9_)  &  n_n524  &  n_n535  &  n_n195 ) ;
 assign n_n4471 = ( n_n518  &  n_n455  &  wire23 ) ;
 assign n_n4490 = ( wire13  &  n_n532  &  n_n500 ) ;
 assign n_n4479 = ( n_n455  &  wire11  &  n_n509 ) ;
 assign n_n901 = ( n_n4478 ) | ( n_n4477 ) | ( n_n4479 ) ;
 assign wire14120 = ( n_n4463 ) | ( n_n4466 ) | ( n_n4465 ) ;
 assign n_n3358 = ( wire14120 ) | ( wire128 ) | ( wire291 ) | ( _26304 ) ;
 assign wire14126 = ( _26306 ) | ( _26307 ) ;
 assign wire14127 = ( n_n4467 ) | ( n_n4470 ) | ( n_n4489 ) | ( n_n4469 ) ;
 assign wire14131 = ( wire184 ) | ( n_n901 ) | ( wire787 ) | ( wire14128 ) ;
 assign n_n3285 = ( n_n3358 ) | ( wire14126 ) | ( wire14127 ) | ( wire14131 ) ;
 assign n_n4423 = ( n_n473  &  n_n536  &  wire23 ) ;
 assign n_n4421 = ( n_n473  &  n_n536  &  wire20 ) ;
 assign wire84 = ( i_9_  &  n_n464  &  n_n536  &  n_n532 ) | ( (~ i_9_)  &  n_n464  &  n_n536  &  n_n532 ) ;
 assign n_n4446 = ( wire13  &  n_n528  &  n_n535 ) ;
 assign wire470 = ( n_n4445 ) | ( n_n4444 ) | ( n_n4446 ) ;
 assign n_n4630 = ( wire10  &  n_n520  &  n_n500 ) ;
 assign n_n5065 = ( wire25  &  n_n464  &  n_n195 ) ;
 assign n_n5287 = ( n_n65  &  n_n491  &  wire23 ) ;
 assign n_n5281 = ( n_n65  &  n_n491  &  wire22 ) ;
 assign n_n5268 = ( wire19  &  n_n522  &  n_n500 ) ;
 assign n_n5261 = ( n_n65  &  wire15  &  n_n500 ) ;
 assign wire13709 = ( n_n5293 ) | ( n_n5240 ) | ( n_n5261 ) ;
 assign wire13710 = ( n_n5274 ) | ( n_n5300 ) | ( n_n5254 ) | ( n_n5287 ) ;
 assign n_n4332 = ( wire16  &  n_n518  &  n_n530 ) ;
 assign n_n4329 = ( wire25  &  n_n518  &  n_n536 ) ;
 assign n_n4448 = ( n_n526  &  wire13  &  n_n535 ) ;
 assign n_n4449 = ( wire22  &  n_n455  &  n_n535 ) ;
 assign n_n4447 = ( n_n455  &  wire11  &  n_n535 ) ;
 assign n_n5029 = ( n_n491  &  n_n195  &  wire20 ) ;
 assign n_n4468 = ( n_n522  &  n_n518  &  wire13 ) ;
 assign n_n3162 = ( n_n4467 ) | ( n_n4466 ) | ( n_n4468 ) ;
 assign n_n4472 = ( wire13  &  n_n534  &  n_n509 ) ;
 assign n_n4469 = ( n_n518  &  n_n455  &  wire20 ) ;
 assign n_n4474 = ( wire13  &  n_n532  &  n_n509 ) ;
 assign wire15423 = ( n_n4472 ) | ( n_n4469 ) | ( wire15421 ) ;
 assign n_n3001 = ( n_n4479 ) | ( n_n3162 ) | ( n_n4474 ) | ( wire15423 ) ;
 assign wire465 = ( i_9_  &  n_n390  &  n_n509  &  n_n520 ) | ( (~ i_9_)  &  n_n390  &  n_n509  &  n_n520 ) ;
 assign n_n4620 = ( wire10  &  n_n500  &  n_n530 ) ;
 assign n_n5001 = ( wire25  &  n_n195  &  n_n500 ) ;
 assign n_n2601 = ( n_n4837 ) | ( n_n4841 ) | ( n_n3461 ) | ( wire14894 ) ;
 assign n_n2602 = ( n_n4824 ) | ( n_n4823 ) | ( wire14898 ) | ( wire14899 ) ;
 assign wire14904 = ( n_n4856 ) | ( n_n4853 ) | ( n_n4858 ) | ( n_n4845 ) ;
 assign wire14905 = ( n_n4852 ) | ( wire11768 ) | ( wire14903 ) ;
 assign n_n4867 = ( wire21  &  n_n509  &  n_n260 ) ;
 assign n_n4866 = ( n_n524  &  n_n509  &  wire17 ) ;
 assign n_n4889 = ( wire25  &  n_n491  &  n_n260 ) ;
 assign wire12179 = ( i_9_  &  n_n491  &  n_n532  &  n_n260 ) | ( (~ i_9_)  &  n_n491  &  n_n532  &  n_n260 ) ;
 assign n_n2597 = ( n_n3450 ) | ( wire49 ) | ( _388 ) | ( _27584 ) ;
 assign n_n4863 = ( wire11  &  n_n509  &  n_n260 ) ;
 assign n_n2727 = ( n_n4859 ) | ( n_n4860 ) | ( n_n4861 ) ;
 assign wire14927 = ( wire85 ) | ( n_n4197 ) | ( wire12225 ) | ( wire14924 ) ;
 assign n_n4965 = ( n_n535  &  n_n195  &  wire20 ) ;
 assign wire228 = ( i_9_  &  n_n526  &  n_n518  &  n_n195 ) | ( (~ i_9_)  &  n_n526  &  n_n518  &  n_n195 ) ;
 assign n_n2611 = ( n_n4710 ) | ( n_n4709 ) | ( n_n4219 ) | ( wire15008 ) ;
 assign wire15011 = ( n_n4737 ) | ( n_n4738 ) | ( n_n4723 ) ;
 assign wire15012 = ( n_n4712 ) | ( n_n4736 ) | ( n_n4722 ) | ( n_n4721 ) ;
 assign wire15016 = ( wire13246 ) | ( n_n856 ) | ( _364 ) | ( _27671 ) ;
 assign wire315 = ( i_9_  &  n_n482  &  n_n534  &  n_n325 ) | ( (~ i_9_)  &  n_n482  &  n_n534  &  n_n325 ) ;
 assign n_n4321 = ( wire22  &  n_n536  &  n_n535 ) ;
 assign n_n4972 = ( n_n518  &  wire18  &  n_n530 ) ;
 assign n_n5118 = ( n_n509  &  n_n528  &  wire12 ) ;
 assign n_n5119 = ( wire11  &  n_n509  &  n_n130 ) ;
 assign n_n5229 = ( n_n65  &  wire15  &  n_n518 ) ;
 assign n_n5228 = ( wire19  &  n_n518  &  n_n530 ) ;
 assign n_n5295 = ( n_n65  &  n_n482  &  wire11 ) ;
 assign n_n4540 = ( n_n473  &  wire13  &  n_n530 ) ;
 assign n_n4536 = ( n_n473  &  wire13  &  n_n534 ) ;
 assign n_n4532 = ( n_n482  &  n_n522  &  wire13 ) ;
 assign n_n4541 = ( n_n473  &  wire15  &  n_n455 ) ;
 assign wire416 = ( i_9_  &  n_n473  &  n_n455  &  n_n528 ) | ( (~ i_9_)  &  n_n473  &  n_n455  &  n_n528 ) ;
 assign n_n4681 = ( wire25  &  n_n464  &  n_n390 ) ;
 assign n_n4679 = ( n_n473  &  n_n390  &  wire23 ) ;
 assign n_n4677 = ( n_n473  &  n_n390  &  wire20 ) ;
 assign n_n4678 = ( n_n473  &  wire10  &  n_n520 ) ;
 assign wire81 = ( n_n464  &  wire10  &  n_n532 ) ;
 assign wire16404 = ( n_n4669 ) | ( n_n4670 ) | ( wire81 ) ;
 assign wire16405 = ( n_n4673 ) | ( n_n4676 ) | ( n_n4681 ) | ( n_n4679 ) ;
 assign wire414 = ( i_9_  &  n_n509  &  n_n528  &  n_n130 ) | ( (~ i_9_)  &  n_n509  &  n_n528  &  n_n130 ) ;
 assign wire345 = ( wire16  &  n_n532  &  n_n500 ) | ( wire16  &  n_n534  &  n_n500 ) ;
 assign wire164 = ( i_9_  &  n_n526  &  n_n491  &  n_n325 ) | ( (~ i_9_)  &  n_n526  &  n_n491  &  n_n325 ) ;
 assign n_n4465 = ( wire22  &  n_n518  &  n_n455 ) ;
 assign n_n4443 = ( n_n455  &  wire24  &  n_n535 ) ;
 assign n_n5121 = ( wire22  &  n_n509  &  n_n130 ) ;
 assign n_n5122 = ( n_n524  &  n_n509  &  wire12 ) ;
 assign n_n4486 = ( wire13  &  n_n509  &  n_n520 ) ;
 assign n_n4484 = ( n_n522  &  wire13  &  n_n509 ) ;
 assign wire199 = ( wire22  &  n_n455  &  n_n509 ) | ( n_n455  &  wire11  &  n_n509 ) ;
 assign n_n4893 = ( wire15  &  n_n491  &  n_n260 ) ;
 assign wire154 = ( i_9_  &  n_n482  &  n_n532  &  n_n260 ) | ( (~ i_9_)  &  n_n482  &  n_n532  &  n_n260 ) ;
 assign wire16784 = ( n_n4902 ) | ( n_n4856 ) | ( n_n4894 ) | ( n_n4854 ) ;
 assign wire16785 = ( n_n4865 ) | ( n_n4905 ) | ( n_n4893 ) | ( wire154 ) ;
 assign n_n2095 = ( wire16784 ) | ( wire16785 ) ;
 assign n_n5168 = ( n_n482  &  n_n526  &  wire12 ) ;
 assign wire16795 = ( n_n5142 ) | ( n_n5168 ) | ( wire679 ) ;
 assign wire16796 = ( n_n5123 ) | ( n_n5131 ) | ( n_n5137 ) | ( n_n5146 ) ;
 assign n_n2091 = ( n_n5193 ) | ( n_n5182 ) | ( wire16795 ) | ( wire16796 ) ;
 assign n_n4973 = ( wire15  &  n_n518  &  n_n195 ) ;
 assign wire16790 = ( n_n5034 ) | ( n_n5099 ) | ( n_n5097 ) | ( n_n5019 ) ;
 assign n_n2084 = ( n_n2091 ) | ( wire16804 ) | ( _29050 ) | ( _29051 ) ;
 assign n_n4377 = ( wire25  &  n_n491  &  n_n536 ) ;
 assign n_n4710 = ( wire14  &  n_n535  &  n_n520 ) ;
 assign n_n4709 = ( n_n325  &  n_n535  &  wire20 ) ;
 assign n_n4765 = ( wire15  &  n_n491  &  n_n325 ) ;
 assign n_n4603 = ( wire24  &  n_n390  &  n_n509 ) ;
 assign n_n4604 = ( wire10  &  n_n509  &  n_n530 ) ;
 assign n_n2037 = ( n_n4600 ) | ( n_n4603 ) | ( n_n4604 ) ;
 assign n_n4588 = ( n_n518  &  wire10  &  n_n530 ) ;
 assign n_n4595 = ( n_n518  &  wire21  &  n_n390 ) ;
 assign wire16038 = ( wire45 ) | ( n_n4591 ) | ( n_n4592 ) ;
 assign n_n1877 = ( n_n2037 ) | ( n_n4588 ) | ( n_n4595 ) | ( wire16038 ) ;
 assign wire12309 = ( n_n5064 ) | ( n_n5058 ) | ( wire755 ) ;
 assign wire12310 = ( n_n5060 ) | ( n_n5055 ) | ( n_n5059 ) | ( n_n5056 ) ;
 assign n_n1450 = ( n_n5067 ) | ( n_n5061 ) | ( wire12309 ) | ( wire12310 ) ;
 assign n_n5152 = ( n_n526  &  n_n491  &  wire12 ) ;
 assign n_n5149 = ( wire15  &  n_n491  &  n_n130 ) ;
 assign wire195 = ( i_9_  &  n_n491  &  n_n520  &  n_n130 ) | ( (~ i_9_)  &  n_n491  &  n_n520  &  n_n130 ) ;
 assign wire358 = ( i_9_  &  n_n491  &  n_n524  &  n_n130 ) | ( (~ i_9_)  &  n_n491  &  n_n524  &  n_n130 ) ;
 assign wire406 = ( i_9_  &  n_n491  &  n_n528  &  n_n130 ) | ( (~ i_9_)  &  n_n491  &  n_n528  &  n_n130 ) ;
 assign n_n5288 = ( n_n482  &  wire19  &  n_n534 ) ;
 assign n_n4751 = ( wire11  &  n_n325  &  n_n500 ) ;
 assign wire12122 = ( n_n4954 ) | ( wire771 ) | ( wire772 ) ;
 assign wire12123 = ( n_n4987 ) | ( n_n5005 ) | ( wire12120 ) ;
 assign n_n1333 = ( n_n4971 ) | ( n_n4972 ) | ( wire12122 ) | ( wire12123 ) ;
 assign n_n4435 = ( n_n464  &  wire21  &  n_n536 ) ;
 assign n_n4626 = ( n_n524  &  wire10  &  n_n500 ) ;
 assign n_n4627 = ( wire21  &  n_n390  &  n_n500 ) ;
 assign n_n4625 = ( wire22  &  n_n390  &  n_n500 ) ;
 assign n_n4660 = ( n_n482  &  n_n522  &  wire10 ) ;
 assign n_n4719 = ( n_n518  &  wire11  &  n_n325 ) ;
 assign n_n4954 = ( n_n532  &  n_n535  &  wire18 ) ;
 assign n_n4955 = ( wire24  &  n_n535  &  n_n195 ) ;
 assign n_n5133 = ( wire15  &  n_n130  &  n_n500 ) ;
 assign n_n5138 = ( n_n524  &  wire12  &  n_n500 ) ;
 assign n_n5139 = ( wire21  &  n_n130  &  n_n500 ) ;
 assign n_n5309 = ( n_n473  &  n_n65  &  wire15 ) ;
 assign n_n4387 = ( n_n491  &  wire21  &  n_n536 ) ;
 assign wire420 = ( n_n491  &  wire22  &  n_n536 ) | ( n_n491  &  n_n536  &  wire11 ) ;
 assign n_n4619 = ( wire24  &  n_n390  &  n_n500 ) ;
 assign wire179 = ( i_9_  &  n_n473  &  n_n532  &  n_n325 ) | ( (~ i_9_)  &  n_n473  &  n_n532  &  n_n325 ) ;
 assign n_n4750 = ( wire14  &  n_n528  &  n_n500 ) ;
 assign n_n4745 = ( wire25  &  n_n325  &  n_n500 ) ;
 assign n_n4736 = ( n_n526  &  n_n509  &  wire14 ) ;
 assign wire293 = ( wire21  &  n_n509  &  n_n325 ) | ( n_n509  &  n_n325  &  wire20 ) ;
 assign n_n4722 = ( n_n524  &  n_n518  &  wire14 ) ;
 assign n_n4721 = ( wire22  &  n_n518  &  n_n325 ) ;
 assign wire457 = ( _22059 ) | ( wire22  &  n_n518  &  n_n325 ) ;
 assign n_n5159 = ( n_n491  &  n_n130  &  wire23 ) ;
 assign n_n5160 = ( n_n482  &  n_n534  &  wire12 ) ;
 assign wire287 = ( i_9_  &  n_n522  &  n_n491  &  n_n130 ) | ( (~ i_9_)  &  n_n522  &  n_n491  &  n_n130 ) ;
 assign n_n5169 = ( n_n482  &  wire22  &  n_n130 ) ;
 assign wire33 = ( i_9_  &  n_n482  &  n_n130  &  n_n530 ) | ( (~ i_9_)  &  n_n482  &  n_n130  &  n_n530 ) ;
 assign wire107 = ( i_9_  &  n_n482  &  n_n524  &  n_n130 ) | ( (~ i_9_)  &  n_n482  &  n_n524  &  n_n130 ) ;
 assign wire113 = ( i_9_  &  n_n473  &  n_n526  &  n_n130 ) | ( (~ i_9_)  &  n_n473  &  n_n526  &  n_n130 ) ;
 assign wire254 = ( i_9_  &  n_n482  &  n_n528  &  n_n130 ) | ( (~ i_9_)  &  n_n482  &  n_n528  &  n_n130 ) ;
 assign n_n4658 = ( n_n482  &  n_n524  &  wire10 ) ;
 assign n_n5108 = ( n_n522  &  n_n518  &  wire12 ) ;
 assign n_n4510 = ( n_n491  &  wire13  &  n_n528 ) ;
 assign n_n4424 = ( n_n464  &  wire16  &  n_n534 ) ;
 assign n_n4498 = ( n_n524  &  wire13  &  n_n500 ) ;
 assign n_n4591 = ( n_n518  &  wire11  &  n_n390 ) ;
 assign n_n4663 = ( n_n482  &  n_n390  &  wire23 ) ;
 assign n_n4698 = ( n_n532  &  wire14  &  n_n535 ) ;
 assign n_n4705 = ( wire22  &  n_n325  &  n_n535 ) ;
 assign n_n4805 = ( n_n473  &  n_n325  &  wire20 ) ;
 assign n_n4841 = ( wire25  &  n_n518  &  n_n260 ) ;
 assign n_n4944 = ( n_n526  &  n_n464  &  wire17 ) ;
 assign n_n5068 = ( n_n464  &  wire18  &  n_n530 ) ;
 assign n_n5187 = ( n_n473  &  wire21  &  n_n130 ) ;
 assign n_n5199 = ( n_n464  &  wire11  &  n_n130 ) ;
 assign n_n5260 = ( wire19  &  n_n500  &  n_n530 ) ;
 assign n_n5272 = ( wire19  &  n_n491  &  n_n534 ) ;
 assign n_n4405 = ( n_n482  &  n_n536  &  wire20 ) ;
 assign n_n4406 = ( n_n482  &  wire16  &  n_n520 ) ;
 assign n_n4462 = ( n_n518  &  wire13  &  n_n528 ) ;
 assign n_n4501 = ( n_n455  &  wire20  &  n_n500 ) ;
 assign n_n4684 = ( n_n464  &  wire10  &  n_n530 ) ;
 assign n_n4222 = ( n_n4683 ) | ( wire81 ) | ( n_n4684 ) ;
 assign n_n4741 = ( n_n509  &  n_n325  &  wire20 ) ;
 assign n_n4740 = ( n_n522  &  n_n509  &  wire14 ) ;
 assign n_n4819 = ( n_n464  &  wire21  &  n_n325 ) ;
 assign n_n5077 = ( n_n464  &  n_n195  &  wire20 ) ;
 assign n_n5221 = ( n_n65  &  n_n535  &  wire20 ) ;
 assign n_n5220 = ( wire19  &  n_n522  &  n_n535 ) ;
 assign n_n834 = ( n_n4849 ) | ( n_n4850 ) | ( n_n4848 ) ;
 assign n_n5134 = ( n_n528  &  wire12  &  n_n500 ) ;
 assign n_n5125 = ( n_n509  &  wire20  &  n_n130 ) ;
 assign wire336 = ( n_n522  &  n_n509  &  wire12 ) | ( n_n509  &  n_n520  &  wire12 ) ;
 assign wire13322 = ( n_n5130 ) | ( n_n5127 ) | ( wire336 ) ;
 assign wire13323 = ( n_n5121 ) | ( n_n5122 ) | ( n_n5125 ) | ( wire13320 ) ;
 assign wire13325 = ( wire13283 ) | ( wire13284 ) | ( wire13287 ) | ( wire13288 ) ;
 assign wire13327 = ( wire13303 ) | ( wire13304 ) | ( wire13317 ) | ( wire13318 ) ;
 assign n_n3988 = ( wire13322 ) | ( wire13323 ) | ( wire13325 ) | ( wire13327 ) ;
 assign n_n5290 = ( n_n482  &  wire19  &  n_n532 ) ;
 assign n_n5291 = ( n_n65  &  n_n482  &  wire24 ) ;
 assign n_n5292 = ( n_n482  &  wire19  &  n_n530 ) ;
 assign n_n5304 = ( n_n473  &  wire19  &  n_n534 ) ;
 assign wire13329 = ( n_n5305 ) | ( n_n5306 ) | ( wire63 ) ;
 assign wire13347 = ( n_n5266 ) | ( n_n5271 ) | ( n_n5270 ) | ( wire77 ) ;
 assign wire441 = ( i_9_  &  n_n65  &  n_n522  &  n_n491 ) | ( (~ i_9_)  &  n_n65  &  n_n522  &  n_n491 ) ;
 assign wire13365 = ( wire13354 ) | ( wire13355 ) | ( wire13359 ) | ( wire13360 ) ;
 assign wire13374 = ( wire13329 ) | ( wire13372 ) | ( _25847 ) | ( _25860 ) ;
 assign n_n3987 = ( wire13374 ) | ( _25825 ) | ( _25826 ) | ( _25862 ) ;
 assign n_n4410 = ( n_n473  &  wire16  &  n_n532 ) ;
 assign n_n4652 = ( n_n482  &  wire10  &  n_n530 ) ;
 assign n_n4650 = ( n_n482  &  wire10  &  n_n532 ) ;
 assign wire14658 = ( n_n5055 ) | ( n_n5056 ) | ( n_n5051 ) ;
 assign wire14659 = ( n_n5048 ) | ( n_n5047 ) | ( wire14656 ) ;
 assign n_n3681 = ( n_n5045 ) | ( n_n5053 ) | ( wire14658 ) | ( wire14659 ) ;
 assign wire14661 = ( n_n5027 ) | ( n_n5028 ) | ( n_n5031 ) ;
 assign wire14662 = ( n_n5024 ) | ( wire253 ) | ( wire13400 ) ;
 assign wire14667 = ( n_n1570 ) | ( n_n5044 ) | ( wire14665 ) | ( _26834 ) ;
 assign wire159 = ( n_n464  &  wire11  &  n_n195 ) | ( n_n464  &  wire24  &  n_n195 ) ;
 assign n_n5226 = ( wire19  &  n_n518  &  n_n532 ) ;
 assign n_n5218 = ( wire19  &  n_n524  &  n_n535 ) ;
 assign wire435 = ( wire19  &  n_n522  &  n_n509 ) | ( wire19  &  n_n524  &  n_n509 ) ;
 assign n_n5153 = ( n_n491  &  wire22  &  n_n130 ) ;
 assign n_n5021 = ( wire15  &  n_n491  &  n_n195 ) ;
 assign n_n4654 = ( n_n482  &  wire10  &  n_n528 ) ;
 assign wire140 = ( i_9_  &  n_n482  &  n_n532  &  n_n390 ) | ( (~ i_9_)  &  n_n482  &  n_n532  &  n_n390 ) ;
 assign wire391 = ( i_9_  &  n_n482  &  n_n526  &  n_n390 ) | ( (~ i_9_)  &  n_n482  &  n_n526  &  n_n390 ) ;
 assign n_n4665 = ( wire25  &  n_n473  &  n_n390 ) ;
 assign wire72 = ( n_n482  &  wire21  &  n_n390 ) | ( n_n482  &  n_n390  &  wire20 ) ;
 assign wire418 = ( i_9_  &  n_n464  &  n_n390  &  n_n534 ) | ( (~ i_9_)  &  n_n464  &  n_n390  &  n_n534 ) ;
 assign wire248 = ( wire21  &  n_n509  &  n_n195 ) | ( n_n509  &  n_n195  &  wire20 ) ;
 assign n_n4394 = ( n_n482  &  wire16  &  n_n532 ) ;
 assign wire14168 = ( n_n4398 ) | ( n_n4405 ) | ( n_n4406 ) ;
 assign n_n3363 = ( wire14168 ) | ( _26246 ) | ( _26247 ) | ( _26248 ) ;
 assign wire14173 = ( n_n4414 ) | ( n_n4411 ) | ( n_n4412 ) ;
 assign n_n3362 = ( wire14173 ) | ( wire79 ) | ( wire14171 ) | ( _26253 ) ;
 assign wire14178 = ( n_n4392 ) | ( n_n4384 ) | ( wire425 ) ;
 assign wire14179 = ( n_n4388 ) | ( n_n4391 ) | ( n_n4390 ) | ( wire14177 ) ;
 assign n_n3287 = ( n_n3363 ) | ( n_n3362 ) | ( wire14178 ) | ( wire14179 ) ;
 assign n_n4279 = ( _25342 ) | ( wire25  &  n_n518  &  n_n536 ) ;
 assign wire14183 = ( wire198 ) | ( wire106 ) ;
 assign wire363 = ( n_n4318 ) | ( n_n4321 ) | ( wire13512 ) ;
 assign n_n3370 = ( wire363 ) | ( wire364 ) | ( _708 ) | ( _26294 ) ;
 assign wire156 = ( i_9_  &  n_n518  &  n_n536  &  n_n520 ) | ( (~ i_9_)  &  n_n518  &  n_n536  &  n_n520 ) ;
 assign wire14163 = ( wire11607 ) | ( wire423 ) | ( wire14160 ) | ( _26270 ) ;
 assign wire14164 = ( wire14153 ) | ( wire14154 ) | ( wire14158 ) | ( wire14159 ) ;
 assign wire14195 = ( wire14183 ) | ( n_n3370 ) | ( _26291 ) | ( _26299 ) ;
 assign n_n3262 = ( n_n3287 ) | ( wire14163 ) | ( wire14164 ) | ( wire14195 ) ;
 assign n_n4896 = ( n_n526  &  n_n491  &  wire17 ) ;
 assign n_n4428 = ( n_n464  &  wire16  &  n_n530 ) ;
 assign wire403 = ( n_n518  &  wire13  &  n_n532 ) | ( n_n518  &  wire13  &  n_n534 ) ;
 assign n_n4499 = ( wire21  &  n_n455  &  n_n500 ) ;
 assign n_n4545 = ( n_n473  &  wire22  &  n_n455 ) ;
 assign wire471 = ( i_9_  &  n_n522  &  n_n464  &  n_n455 ) | ( (~ i_9_)  &  n_n522  &  n_n464  &  n_n455 ) ;
 assign n_n4376 = ( n_n491  &  wire16  &  n_n534 ) ;
 assign n_n3176 = ( wire423 ) | ( n_n491  &  wire16  &  n_n532 ) ;
 assign n_n4585 = ( wire25  &  n_n518  &  n_n390 ) ;
 assign n_n4873 = ( wire25  &  n_n260  &  n_n500 ) ;
 assign n_n4932 = ( n_n473  &  n_n522  &  wire17 ) ;
 assign n_n4592 = ( n_n526  &  n_n518  &  wire10 ) ;
 assign n_n5052 = ( n_n473  &  wire18  &  n_n530 ) ;
 assign wire15601 = ( n_n5055 ) | ( n_n5056 ) | ( n_n5052 ) ;
 assign wire15602 = ( n_n5049 ) | ( n_n5046 ) | ( wire15598 ) ;
 assign n_n2956 = ( n_n5047 ) | ( n_n5051 ) | ( wire15601 ) | ( wire15602 ) ;
 assign n_n5235 = ( n_n65  &  n_n518  &  wire21 ) ;
 assign n_n5234 = ( wire19  &  n_n524  &  n_n518 ) ;
 assign n_n5286 = ( wire19  &  n_n491  &  n_n520 ) ;
 assign n_n5285 = ( n_n65  &  n_n491  &  wire20 ) ;
 assign n_n1764 = ( n_n4667 ) | ( n_n4664 ) | ( n_n4663 ) ;
 assign n_n3810 = ( n_n4898 ) | ( n_n4897 ) | ( n_n4896 ) ;
 assign n_n2304 = ( n_n5130 ) | ( n_n5133 ) | ( n_n5134 ) ;
 assign n_n5256 = ( wire19  &  n_n534  &  n_n500 ) ;
 assign n_n5253 = ( n_n65  &  n_n509  &  wire20 ) ;
 assign n_n1139 = ( n_n5255 ) | ( n_n5256 ) | ( n_n5253 ) ;
 assign n_n4414 = ( n_n473  &  wire16  &  n_n528 ) ;
 assign wire215 = ( i_9_  &  n_n473  &  n_n536  &  n_n520 ) | ( (~ i_9_)  &  n_n473  &  n_n536  &  n_n520 ) ;
 assign wire16691 = ( wire62 ) | ( wire181 ) ;
 assign wire16692 = ( n_n5232 ) | ( n_n5237 ) | ( wire183 ) ;
 assign wire16696 = ( n_n5251 ) | ( wire435 ) | ( n_n1139 ) | ( wire16693 ) ;
 assign n_n5170 = ( n_n482  &  n_n524  &  wire12 ) ;
 assign wire168 = ( i_9_  &  n_n482  &  n_n534  &  n_n130 ) | ( (~ i_9_)  &  n_n482  &  n_n534  &  n_n130 ) ;
 assign wire16682 = ( n_n5215 ) | ( n_n2291 ) | ( wire13350 ) | ( wire16679 ) ;
 assign wire16683 = ( wire16673 ) | ( wire16674 ) | ( wire16677 ) | ( wire16678 ) ;
 assign n_n2214 = ( wire166 ) | ( n_n5061 ) | ( wire669 ) | ( _28888 ) ;
 assign wire16753 = ( wire203 ) | ( wire205 ) ;
 assign wire16754 = ( n_n5270 ) | ( n_n5269 ) | ( wire438 ) ;
 assign wire16758 = ( n_n5280 ) | ( wire16755 ) | ( _27476 ) | ( _28931 ) ;
 assign n_n5333 = ( n_n65  &  n_n464  &  wire20 ) ;
 assign n_n4429 = ( wire15  &  n_n464  &  n_n536 ) ;
 assign n_n4813 = ( wire15  &  n_n464  &  n_n325 ) ;
 assign n_n4815 = ( n_n464  &  wire11  &  n_n325 ) ;
 assign wire85 = ( n_n464  &  wire14  &  n_n528 ) ;
 assign wire16811 = ( n_n4847 ) | ( n_n4817 ) | ( wire85 ) ;
 assign wire16812 = ( n_n4827 ) | ( n_n4816 ) | ( n_n4833 ) | ( n_n4813 ) ;
 assign n_n2096 = ( n_n4838 ) | ( n_n4815 ) | ( wire16811 ) | ( wire16812 ) ;
 assign n_n4715 = ( n_n518  &  wire24  &  n_n325 ) ;
 assign n_n4714 = ( n_n518  &  n_n532  &  wire14 ) ;
 assign n_n5225 = ( wire25  &  n_n65  &  n_n518 ) ;
 assign n_n5224 = ( wire19  &  n_n518  &  n_n534 ) ;
 assign n_n1530 = ( n_n5226 ) | ( n_n5225 ) | ( n_n5224 ) ;
 assign wire437 = ( i_9_  &  n_n482  &  n_n526  &  n_n130 ) | ( (~ i_9_)  &  n_n482  &  n_n526  &  n_n130 ) ;
 assign n_n5279 = ( n_n65  &  n_n491  &  wire11 ) ;
 assign n_n5277 = ( n_n65  &  wire15  &  n_n491 ) ;
 assign n_n4708 = ( n_n522  &  wire14  &  n_n535 ) ;
 assign n_n4706 = ( n_n524  &  wire14  &  n_n535 ) ;
 assign wire366 = ( n_n518  &  n_n532  &  wire14 ) | ( n_n518  &  n_n534  &  wire14 ) ;
 assign n_n4427 = ( n_n464  &  n_n536  &  wire24 ) ;
 assign n_n4716 = ( n_n518  &  wire14  &  n_n530 ) ;
 assign n_n4807 = ( n_n473  &  n_n325  &  wire23 ) ;
 assign n_n1162 = ( n_n5136 ) | ( n_n5135 ) | ( n_n5134 ) ;
 assign n_n5312 = ( n_n473  &  wire19  &  n_n526 ) ;
 assign n_n5313 = ( n_n473  &  n_n65  &  wire22 ) ;
 assign n_n4596 = ( n_n522  &  n_n518  &  wire10 ) ;
 assign wire256 = ( wire10  &  n_n532  &  n_n509 ) | ( wire10  &  n_n509  &  n_n530 ) ;
 assign wire11912 = ( n_n5131 ) | ( n_n5132 ) | ( wire336 ) ;
 assign n_n1059 = ( n_n5128 ) | ( n_n5133 ) | ( n_n1162 ) | ( wire11912 ) ;
 assign wire11914 = ( i_9_  &  n_n518  &  n_n520  &  n_n130 ) | ( (~ i_9_)  &  n_n518  &  n_n520  &  n_n130 ) ;
 assign wire28 = ( wire335 ) | ( n_n5115 ) | ( wire11914 ) ;
 assign n_n4672 = ( n_n473  &  n_n526  &  wire10 ) ;
 assign n_n4418 = ( n_n473  &  n_n524  &  wire16 ) ;
 assign n_n4688 = ( n_n526  &  n_n464  &  wire10 ) ;
 assign n_n4961 = ( wire22  &  n_n535  &  n_n195 ) ;
 assign n_n5140 = ( n_n522  &  wire12  &  n_n500 ) ;
 assign n_n5194 = ( n_n464  &  n_n532  &  wire12 ) ;
 assign n_n5259 = ( n_n65  &  wire24  &  n_n500 ) ;
 assign n_n5271 = ( n_n65  &  wire23  &  n_n500 ) ;
 assign n_n4537 = ( wire25  &  n_n473  &  n_n455 ) ;
 assign n_n4614 = ( wire10  &  n_n509  &  n_n520 ) ;
 assign wire13202 = ( n_n4911 ) | ( n_n4912 ) | ( n_n4915 ) ;
 assign wire13203 = ( n_n4909 ) | ( n_n4916 ) | ( wire154 ) ;
 assign n_n4058 = ( n_n4917 ) | ( n_n4914 ) | ( wire13202 ) | ( wire13203 ) ;
 assign n_n4016 = ( n_n4083 ) | ( wire13445 ) | ( wire13446 ) | ( wire13452 ) ;
 assign wire13468 = ( wire13457 ) | ( wire13458 ) | ( wire13462 ) | ( wire13463 ) ;
 assign n_n3993 = ( n_n4016 ) | ( wire13481 ) | ( _25314 ) | ( _25315 ) ;
 assign n_n4021 = ( n_n4099 ) | ( wire13538 ) | ( _25336 ) | ( _25337 ) ;
 assign wire13520 = ( wire363 ) | ( wire13509 ) | ( wire13510 ) | ( wire13515 ) ;
 assign n_n3995 = ( n_n4021 ) | ( wire13546 ) | ( _25381 ) | ( _25382 ) ;
 assign wire12471 = ( i_9_  &  n_n518  &  n_n455  &  n_n530 ) | ( (~ i_9_)  &  n_n518  &  n_n455  &  n_n530 ) ;
 assign wire55 = ( wire12471 ) | ( n_n518  &  wire13  &  n_n528 ) ;
 assign wire13553 = ( n_n4455 ) | ( wire403 ) | ( wire13550 ) | ( wire13552 ) ;
 assign wire13554 = ( wire13438 ) | ( wire13439 ) | ( wire13501 ) | ( wire13502 ) ;
 assign n_n4707 = ( wire21  &  n_n325  &  n_n535 ) ;
 assign n_n4701 = ( wire15  &  n_n325  &  n_n535 ) ;
 assign n_n4643 = ( n_n491  &  wire21  &  n_n390 ) ;
 assign n_n4642 = ( n_n491  &  n_n524  &  wire10 ) ;
 assign wire14393 = ( n_n4615 ) | ( n_n4618 ) | ( n_n4629 ) | ( n_n4630 ) ;
 assign n_n3716 = ( n_n3861 ) | ( n_n4620 ) | ( n_n4625 ) | ( wire14393 ) ;
 assign wire14398 = ( n_n4648 ) | ( n_n4647 ) | ( n_n4645 ) | ( wire14396 ) ;
 assign n_n3650 = ( n_n3716 ) | ( wire14403 ) | ( wire14404 ) | ( _26648 ) ;
 assign n_n4556 = ( n_n464  &  wire13  &  n_n530 ) ;
 assign wire455 = ( i_9_  &  n_n524  &  n_n464  &  n_n455 ) | ( (~ i_9_)  &  n_n524  &  n_n464  &  n_n455 ) ;
 assign wire91 = ( n_n464  &  wire13  &  n_n520 ) ;
 assign wire430 = ( i_9_  &  n_n464  &  n_n455  &  n_n532 ) | ( (~ i_9_)  &  n_n464  &  n_n455  &  n_n532 ) ;
 assign n_n4609 = ( wire22  &  n_n390  &  n_n509 ) ;
 assign wire14422 = ( n_n4591 ) | ( n_n4592 ) | ( n_n4596 ) ;
 assign wire14423 = ( n_n4593 ) | ( n_n4594 ) | ( wire45 ) ;
 assign n_n3718 = ( n_n4597 ) | ( n_n4588 ) | ( wire14422 ) | ( wire14423 ) ;
 assign wire14419 = ( n_n3871 ) | ( wire455 ) | ( wire671 ) | ( wire14416 ) ;
 assign wire14420 = ( wire14409 ) | ( wire14410 ) | ( wire14414 ) | ( wire14415 ) ;
 assign wire14436 = ( n_n3718 ) | ( wire14428 ) | ( wire14429 ) | ( wire14434 ) ;
 assign n_n4358 = ( wire16  &  n_n509  &  n_n520 ) ;
 assign n_n4493 = ( wire15  &  n_n455  &  n_n500 ) ;
 assign n_n5148 = ( n_n491  &  wire12  &  n_n530 ) ;
 assign n_n3461 = ( n_n4831 ) | ( n_n4832 ) | ( n_n4833 ) ;
 assign wire11769 = ( wire21  &  n_n535  &  n_n260 ) | ( n_n535  &  n_n260  &  wire20 ) ;
 assign n_n3329 = ( n_n3461 ) | ( wire13807 ) | ( _660 ) | ( _26486 ) ;
 assign n_n5126 = ( n_n509  &  n_n520  &  wire12 ) ;
 assign wire13923 = ( n_n5121 ) | ( n_n5122 ) | ( n_n5126 ) ;
 assign wire13924 = ( n_n5131 ) | ( n_n5124 ) | ( n_n5127 ) | ( n_n5132 ) ;
 assign n_n3307 = ( n_n5128 ) | ( n_n5125 ) | ( wire13923 ) | ( wire13924 ) ;
 assign wire13796 = ( n_n2130 ) | ( n_n4204 ) | ( n_n3469 ) | ( wire13790 ) ;
 assign wire13797 = ( wire13788 ) | ( wire13789 ) | ( wire13791 ) | ( wire13792 ) ;
 assign n_n4808 = ( n_n464  &  n_n534  &  wire14 ) ;
 assign wire13803 = ( n_n4825 ) | ( n_n4815 ) | ( n_n4826 ) ;
 assign wire13804 = ( n_n4830 ) | ( wire693 ) | ( wire186 ) ;
 assign n_n3330 = ( n_n4827 ) | ( n_n4822 ) | ( wire13803 ) | ( wire13804 ) ;
 assign wire13813 = ( n_n4857 ) | ( n_n4860 ) | ( n_n4866 ) | ( wire13810 ) ;
 assign n_n3275 = ( n_n3329 ) | ( _26498 ) | ( _26499 ) | ( _26500 ) ;
 assign n_n2710 = ( n_n4942 ) | ( wire59 ) | ( n_n4940 ) ;
 assign wire13855 = ( n_n4898 ) | ( n_n4901 ) | ( n_n4904 ) | ( n_n4897 ) ;
 assign wire13856 = ( n_n4902 ) | ( n_n4907 ) | ( wire49 ) ;
 assign wire13860 = ( n_n3450 ) | ( n_n4883 ) | ( wire13857 ) | ( _26367 ) ;
 assign n_n3274 = ( n_n3326 ) | ( wire13855 ) | ( wire13856 ) | ( wire13860 ) ;
 assign wire13867 = ( wire22  &  n_n464  &  n_n260 ) | ( n_n464  &  wire11  &  n_n260 ) ;
 assign wire58 = ( wire13867 ) | ( n_n526  &  n_n464  &  wire17 ) ;
 assign wire13844 = ( n_n3803 ) | ( wire13833 ) | ( wire13834 ) | ( wire13840 ) ;
 assign n_n3257 = ( n_n3274 ) | ( wire13877 ) | ( _26416 ) | ( _26417 ) ;
 assign wire12778 = ( wire21  &  n_n509  &  n_n325 ) | ( n_n509  &  n_n325  &  wire20 ) ;
 assign wire456 = ( n_n4737 ) | ( n_n4738 ) | ( wire373 ) | ( wire12778 ) ;
 assign n_n4799 = ( n_n473  &  wire11  &  n_n325 ) ;
 assign wire13746 = ( n_n4724 ) | ( n_n4799 ) | ( n_n4723 ) ;
 assign wire13747 = ( n_n4779 ) | ( n_n4786 ) | ( n_n4755 ) | ( n_n4781 ) ;
 assign wire13753 = ( n_n4571 ) | ( n_n4578 ) | ( n_n4570 ) | ( n_n4594 ) ;
 assign n_n4685 = ( wire15  &  n_n464  &  n_n390 ) ;
 assign n_n4520 = ( n_n482  &  wire13  &  n_n534 ) ;
 assign n_n5008 = ( n_n526  &  wire18  &  n_n500 ) ;
 assign n_n4623 = ( wire11  &  n_n390  &  n_n500 ) ;
 assign wire304 = ( n_n522  &  wire17  &  n_n535 ) | ( n_n524  &  wire17  &  n_n535 ) ;
 assign wire14894 = ( n_n4839 ) | ( n_n4840 ) | ( wire304 ) ;
 assign wire14898 = ( n_n4830 ) | ( wire693 ) | ( n_n4818 ) ;
 assign wire14899 = ( n_n4821 ) | ( n_n4822 ) | ( wire14896 ) ;
 assign wire433 = ( i_9_  &  n_n65  &  n_n534  &  n_n500 ) | ( (~ i_9_)  &  n_n65  &  n_n534  &  n_n500 ) ;
 assign n_n5242 = ( wire19  &  n_n532  &  n_n509 ) ;
 assign wire320 = ( n_n65  &  n_n518  &  wire20 ) | ( n_n65  &  n_n518  &  wire23 ) ;
 assign n_n5264 = ( wire19  &  n_n526  &  n_n500 ) ;
 assign n_n5270 = ( wire19  &  n_n520  &  n_n500 ) ;
 assign wire77 = ( i_9_  &  n_n65  &  n_n522  &  n_n500 ) | ( (~ i_9_)  &  n_n65  &  n_n522  &  n_n500 ) ;
 assign wire334 = ( i_9_  &  n_n65  &  n_n524  &  n_n500 ) | ( (~ i_9_)  &  n_n65  &  n_n524  &  n_n500 ) ;
 assign wire149 = ( wire19  &  n_n522  &  n_n464 ) | ( wire19  &  n_n464  &  n_n520 ) ;
 assign n_n5315 = ( n_n473  &  n_n65  &  wire21 ) ;
 assign wire13557 = ( n_n473  &  wire19  &  n_n524 ) | ( n_n473  &  wire19  &  n_n520 ) ;
 assign wire267 = ( wire115 ) | ( n_n5315 ) | ( wire13557 ) ;
 assign wire15195 = ( n_n5303 ) | ( n_n5304 ) | ( wire63 ) ;
 assign wire15198 = ( wire203 ) | ( wire438 ) ;
 assign wire218 = ( i_9_  &  n_n65  &  n_n491  &  n_n524 ) | ( (~ i_9_)  &  n_n65  &  n_n491  &  n_n524 ) ;
 assign wire385 = ( i_9_  &  n_n65  &  n_n518  &  n_n532 ) | ( (~ i_9_)  &  n_n65  &  n_n518  &  n_n532 ) ;
 assign wire399 = ( i_9_  &  n_n536  &  n_n509  &  n_n528 ) | ( (~ i_9_)  &  n_n536  &  n_n509  &  n_n528 ) ;
 assign wire125 = ( wire25  &  n_n491  &  n_n130 ) | ( n_n491  &  wire24  &  n_n130 ) ;
 assign wire16749 = ( n_n5293 ) | ( n_n5296 ) | ( n_n5297 ) | ( n_n5298 ) ;
 assign wire44 = ( i_9_  &  n_n482  &  n_n520  &  n_n130 ) | ( (~ i_9_)  &  n_n482  &  n_n520  &  n_n130 ) ;
 assign wire332 = ( i_9_  &  n_n482  &  n_n522  &  n_n130 ) | ( (~ i_9_)  &  n_n482  &  n_n522  &  n_n130 ) ;
 assign n_n5080 = ( n_n534  &  n_n535  &  wire12 ) ;
 assign wire209 = ( i_9_  &  n_n522  &  n_n464  &  n_n195 ) | ( (~ i_9_)  &  n_n522  &  n_n464  &  n_n195 ) ;
 assign wire90 = ( n_n5075 ) | ( n_n5078 ) | ( n_n5080 ) | ( wire209 ) ;
 assign n_n5090 = ( n_n524  &  n_n535  &  wire12 ) ;
 assign wire13305 = ( i_9_  &  n_n522  &  n_n535  &  n_n130 ) | ( (~ i_9_)  &  n_n522  &  n_n535  &  n_n130 ) ;
 assign wire13306 = ( i_9_  &  n_n526  &  n_n535  &  n_n130 ) | ( (~ i_9_)  &  n_n526  &  n_n535  &  n_n130 ) ;
 assign wire144 = ( n_n5091 ) | ( n_n5090 ) | ( wire13305 ) | ( wire13306 ) ;
 assign wire239 = ( wire10  &  n_n528  &  n_n535 ) | ( wire10  &  n_n535  &  n_n530 ) ;
 assign n_n4411 = ( n_n473  &  n_n536  &  wire24 ) ;
 assign n_n5219 = ( n_n65  &  wire21  &  n_n535 ) ;
 assign wire12156 = ( n_n4982 ) | ( wire134 ) | ( n_n4985 ) | ( n_n4986 ) ;
 assign n_n1521 = ( n_n5272 ) | ( n_n5271 ) | ( n_n5270 ) ;
 assign n_n4528 = ( n_n482  &  n_n526  &  wire13 ) ;
 assign n_n4529 = ( n_n482  &  wire22  &  n_n455 ) ;
 assign n_n5319 = ( n_n473  &  n_n65  &  wire23 ) ;
 assign wire328 = ( i_9_  &  n_n473  &  n_n536  &  n_n530 ) | ( (~ i_9_)  &  n_n473  &  n_n536  &  n_n530 ) ;
 assign n_n4542 = ( n_n473  &  wire13  &  n_n528 ) ;
 assign wire201 = ( i_9_  &  n_n473  &  n_n455  &  n_n530 ) | ( (~ i_9_)  &  n_n473  &  n_n455  &  n_n530 ) ;
 assign n_n4549 = ( n_n473  &  n_n455  &  wire20 ) ;
 assign n_n4691 = ( n_n464  &  wire21  &  n_n390 ) ;
 assign n_n3849 = ( n_n4690 ) | ( n_n4689 ) | ( n_n4691 ) ;
 assign n_n4692 = ( n_n522  &  n_n464  &  wire10 ) ;
 assign wire11862 = ( n_n4685 ) | ( n_n4686 ) | ( n_n4695 ) | ( n_n4696 ) ;
 assign n_n1093 = ( n_n4683 ) | ( n_n3849 ) | ( n_n4692 ) | ( wire11862 ) ;
 assign wire299 = ( i_9_  &  n_n195  &  n_n500  &  n_n530 ) | ( (~ i_9_)  &  n_n195  &  n_n500  &  n_n530 ) ;
 assign n_n1050 = ( wire318 ) | ( wire435 ) | ( n_n1139 ) | ( _22433 ) ;
 assign n_n5269 = ( n_n65  &  wire20  &  n_n500 ) ;
 assign n_n5257 = ( wire25  &  n_n65  &  n_n500 ) ;
 assign wire62 = ( i_9_  &  n_n65  &  n_n532  &  n_n500 ) | ( (~ i_9_)  &  n_n65  &  n_n532  &  n_n500 ) ;
 assign wire92 = ( n_n65  &  wire11  &  n_n500 ) ;
 assign wire409 = ( i_9_  &  n_n65  &  n_n500  &  n_n530 ) | ( (~ i_9_)  &  n_n65  &  n_n500  &  n_n530 ) ;
 assign wire11923 = ( wire19  &  n_n526  &  n_n500 ) | ( wire19  &  n_n524  &  n_n500 ) ;
 assign wire11927 = ( wire62 ) | ( wire92 ) | ( wire11924 ) ;
 assign n_n1048 = ( n_n1521 ) | ( wire438 ) | ( wire333 ) | ( _22464 ) ;
 assign wire63 = ( i_9_  &  n_n65  &  n_n482  &  n_n522 ) | ( (~ i_9_)  &  n_n65  &  n_n482  &  n_n522 ) ;
 assign wire200 = ( n_n482  &  wire19  &  n_n526 ) | ( n_n482  &  wire19  &  n_n524 ) ;
 assign wire11929 = ( n_n5288 ) | ( wire441 ) | ( n_n5286 ) ;
 assign n_n1017 = ( n_n1048 ) | ( wire11939 ) | ( _22494 ) | ( _22495 ) ;
 assign wire11944 = ( n_n5305 ) | ( wire459 ) | ( n_n5306 ) ;
 assign wire11946 = ( wire25  &  n_n65  &  n_n464 ) | ( n_n65  &  n_n464  &  wire24 ) ;
 assign wire175 = ( i_9_  &  n_n65  &  n_n464  &  n_n530 ) | ( (~ i_9_)  &  n_n65  &  n_n464  &  n_n530 ) ;
 assign n_n4686 = ( n_n464  &  wire10  &  n_n528 ) ;
 assign n_n4354 = ( n_n524  &  wire16  &  n_n509 ) ;
 assign n_n5196 = ( n_n464  &  wire12  &  n_n530 ) ;
 assign n_n5203 = ( n_n464  &  wire21  &  n_n130 ) ;
 assign n_n5210 = ( wire19  &  n_n532  &  n_n535 ) ;
 assign n_n5217 = ( n_n65  &  wire22  &  n_n535 ) ;
 assign wire13566 = ( n_n5321 ) | ( n_n5313 ) | ( n_n5319 ) | ( wire13562 ) ;
 assign wire13567 = ( wire175 ) | ( wire13559 ) | ( wire13560 ) | ( wire13561 ) ;
 assign n_n3996 = ( wire267 ) | ( wire13566 ) | ( wire13567 ) ;
 assign n_n4929 = ( n_n473  &  wire22  &  n_n260 ) ;
 assign n_n4766 = ( n_n491  &  wire14  &  n_n528 ) ;
 assign wire447 = ( n_n4770 ) | ( n_n4771 ) | ( wire12393 ) | ( wire164 ) ;
 assign n_n1592 = ( n_n4921 ) | ( n_n4918 ) | ( n_n4919 ) ;
 assign n_n4742 = ( n_n509  &  wire14  &  n_n520 ) ;
 assign n_n4527 = ( n_n482  &  n_n455  &  wire11 ) ;
 assign n_n4713 = ( wire25  &  n_n518  &  n_n325 ) ;
 assign wire14347 = ( n_n4720 ) | ( n_n4719 ) | ( wire14344 ) ;
 assign wire14350 = ( wire221 ) | ( wire442 ) ;
 assign wire14351 = ( n_n4693 ) | ( wire12422 ) | ( wire14349 ) ;
 assign n_n4657 = ( n_n482  &  wire22  &  n_n390 ) ;
 assign wire14363 = ( n_n4688 ) | ( n_n4685 ) | ( n_n4686 ) ;
 assign n_n3711 = ( n_n4222 ) | ( n_n3849 ) | ( wire14363 ) ;
 assign wire14362 = ( n_n4676 ) | ( n_n4679 ) | ( wire418 ) | ( n_n4672 ) ;
 assign n_n3649 = ( n_n3711 ) | ( _27223 ) | ( _27224 ) | ( _27225 ) ;
 assign n_n3724 = ( n_n4524 ) | ( n_n4517 ) | ( n_n3879 ) | ( wire14448 ) ;
 assign wire14453 = ( wire129 ) | ( wire378 ) ;
 assign wire14454 = ( n_n4504 ) | ( n_n4503 ) | ( wire379 ) ;
 assign wire14458 = ( n_n4534 ) | ( wire11543 ) | ( wire14452 ) | ( wire14455 ) ;
 assign n_n3653 = ( n_n3724 ) | ( wire14453 ) | ( wire14454 ) | ( wire14458 ) ;
 assign n_n3729 = ( n_n4461 ) | ( wire14517 ) | ( _600 ) | ( _26776 ) ;
 assign wire14522 = ( n_n4427 ) | ( wire14519 ) | ( wire14520 ) ;
 assign n_n3655 = ( n_n3729 ) | ( _26794 ) | ( _26795 ) | ( _26796 ) ;
 assign n_n5144 = ( n_n491  &  n_n534  &  wire12 ) ;
 assign n_n5143 = ( n_n130  &  wire23  &  n_n500 ) ;
 assign n_n2685 = ( n_n5120 ) | ( n_n5117 ) | ( n_n5119 ) ;
 assign wire13929 = ( n_n5111 ) | ( n_n5112 ) | ( wire335 ) ;
 assign n_n3308 = ( n_n5109 ) | ( n_n5113 ) | ( n_n2685 ) | ( wire13929 ) ;
 assign n_n5007 = ( wire11  &  n_n195  &  n_n500 ) ;
 assign wire211 = ( i_9_  &  n_n522  &  n_n130  &  n_n500 ) | ( (~ i_9_)  &  n_n522  &  n_n130  &  n_n500 ) ;
 assign wire14065 = ( n_n3307 ) | ( n_n3308 ) | ( wire14061 ) | ( wire14062 ) ;
 assign wire14066 = ( wire14042 ) | ( wire14058 ) | ( _26043 ) ;
 assign wire14068 = ( wire13977 ) | ( wire14025 ) | ( _26177 ) ;
 assign n_n4953 = ( wire25  &  n_n535  &  n_n195 ) ;
 assign wire13772 = ( n_n4803 ) | ( n_n4804 ) | ( n_n4818 ) ;
 assign wire13773 = ( n_n4816 ) | ( n_n4811 ) | ( n_n4828 ) | ( n_n4842 ) ;
 assign n_n4334 = ( wire16  &  n_n518  &  n_n528 ) ;
 assign wire158 = ( i_9_  &  n_n473  &  n_n534  &  n_n325 ) | ( (~ i_9_)  &  n_n473  &  n_n534  &  n_n325 ) ;
 assign wire380 = ( n_n473  &  wire14  &  n_n528 ) | ( n_n473  &  wire14  &  n_n530 ) ;
 assign n_n4874 = ( n_n532  &  wire17  &  n_n500 ) ;
 assign wire49 = ( i_9_  &  n_n491  &  n_n260  &  n_n530 ) | ( (~ i_9_)  &  n_n491  &  n_n260  &  n_n530 ) ;
 assign wire87 = ( n_n65  &  n_n518  &  wire11 ) ;
 assign wire182 = ( i_9_  &  n_n65  &  n_n526  &  n_n518 ) | ( (~ i_9_)  &  n_n65  &  n_n526  &  n_n518 ) ;
 assign n_n5215 = ( n_n65  &  wire11  &  n_n535 ) ;
 assign wire220 = ( i_9_  &  n_n522  &  n_n464  &  n_n130 ) | ( (~ i_9_)  &  n_n522  &  n_n464  &  n_n130 ) ;
 assign wire384 = ( n_n65  &  n_n535  &  wire20 ) | ( n_n65  &  n_n535  &  wire23 ) ;
 assign wire454 = ( n_n65  &  wire15  &  n_n535 ) | ( n_n65  &  wire24  &  n_n535 ) ;
 assign n_n4534 = ( n_n482  &  wire13  &  n_n520 ) ;
 assign n_n2630 = ( n_n3162 ) | ( n_n4465 ) | ( n_n4462 ) | ( wire15069 ) ;
 assign wire15065 = ( wire128 ) | ( wire291 ) ;
 assign wire15066 = ( wire368 ) | ( n_n4446 ) | ( wire15063 ) ;
 assign wire15075 = ( wire236 ) | ( n_n910 ) | ( wire15071 ) | ( _27260 ) ;
 assign n_n2558 = ( n_n2630 ) | ( wire15065 ) | ( wire15066 ) | ( wire15075 ) ;
 assign wire15079 = ( n_n4515 ) | ( wire791 ) | ( n_n4518 ) ;
 assign wire15080 = ( n_n4520 ) | ( wire789 ) | ( wire15077 ) ;
 assign n_n2626 = ( n_n4521 ) | ( n_n4511 ) | ( wire15079 ) | ( wire15080 ) ;
 assign wire15094 = ( n_n4510 ) | ( n_n1677 ) | ( wire14200 ) | ( wire15091 ) ;
 assign wire15095 = ( wire15084 ) | ( wire15085 ) | ( wire15089 ) | ( wire15090 ) ;
 assign wire15103 = ( n_n2626 ) | ( wire15061 ) | ( wire15062 ) | ( wire15101 ) ;
 assign wire82 = ( n_n4553 ) | ( n_n4554 ) | ( n_n4552 ) ;
 assign wire783 = ( n_n464  &  n_n455  &  wire23 ) ;
 assign wire11564 = ( n_n524  &  n_n464  &  wire13 ) | ( n_n464  &  wire13  &  n_n520 ) ;
 assign wire224 = ( n_n4568 ) | ( wire471 ) | ( wire783 ) | ( wire11564 ) ;
 assign n_n5248 = ( wire19  &  n_n526  &  n_n509 ) ;
 assign n_n4412 = ( n_n473  &  wire16  &  n_n530 ) ;
 assign n_n5280 = ( wire19  &  n_n526  &  n_n491 ) ;
 assign n_n5195 = ( n_n464  &  wire24  &  n_n130 ) ;
 assign n_n5197 = ( wire15  &  n_n464  &  n_n130 ) ;
 assign n_n5209 = ( wire25  &  n_n65  &  n_n535 ) ;
 assign n_n5208 = ( wire19  &  n_n534  &  n_n535 ) ;
 assign n_n2291 = ( n_n5210 ) | ( n_n5209 ) | ( n_n5208 ) ;
 assign wire451 = ( n_n464  &  n_n532  &  wire12 ) | ( n_n464  &  wire12  &  n_n530 ) ;
 assign n_n4723 = ( n_n518  &  wire21  &  n_n325 ) ;
 assign n_n4892 = ( n_n491  &  wire17  &  n_n530 ) ;
 assign n_n5213 = ( n_n65  &  wire15  &  n_n535 ) ;
 assign n_n1532 = ( n_n5210 ) | ( n_n5209 ) | ( n_n5213 ) ;
 assign wire288 = ( i_9_  &  n_n520  &  n_n130  &  n_n500 ) | ( (~ i_9_)  &  n_n520  &  n_n130  &  n_n500 ) ;
 assign n_n5247 = ( n_n65  &  wire11  &  n_n509 ) ;
 assign wire446 = ( i_9_  &  n_n65  &  n_n526  &  n_n509 ) | ( (~ i_9_)  &  n_n65  &  n_n526  &  n_n509 ) ;
 assign wire12349 = ( n_n5251 ) | ( wire435 ) | ( n_n5257 ) | ( n_n5247 ) ;
 assign n_n1435 = ( n_n5254 ) | ( n_n5259 ) | ( wire446 ) | ( wire12349 ) ;
 assign n_n1103 = ( wire213 ) | ( wire82 ) | ( wire11539 ) | ( _22987 ) ;
 assign wire181 = ( i_9_  &  n_n65  &  n_n518  &  n_n530 ) | ( (~ i_9_)  &  n_n65  &  n_n518  &  n_n530 ) ;
 assign wire452 = ( n_n464  &  n_n528  &  wire12 ) | ( n_n464  &  wire12  &  n_n530 ) ;
 assign n_n5211 = ( n_n65  &  wire24  &  n_n535 ) ;
 assign n_n1111 = ( wire403 ) | ( wire291 ) | ( wire11507 ) | ( _22846 ) ;
 assign wire11511 = ( wire70 ) | ( n_n522  &  wire13  &  n_n509 ) ;
 assign wire11512 = ( n_n4489 ) | ( wire184 ) | ( n_n4486 ) | ( wire787 ) ;
 assign wire11518 = ( n_n4465 ) | ( wire11505 ) | ( wire11515 ) | ( wire11516 ) ;
 assign wire79 = ( i_9_  &  n_n473  &  n_n524  &  n_n536 ) | ( (~ i_9_)  &  n_n473  &  n_n524  &  n_n536 ) ;
 assign wire11543 = ( n_n482  &  n_n455  &  wire20 ) | ( n_n482  &  n_n455  &  wire23 ) ;
 assign n_n3875 = ( wire11543 ) | ( n_n482  &  wire13  &  n_n520 ) ;
 assign wire11602 = ( n_n4399 ) | ( n_n4396 ) | ( wire11599 ) ;
 assign wire11605 = ( wire11591 ) | ( wire11592 ) | ( wire11597 ) | ( wire11598 ) ;
 assign n_n1040 = ( wire11602 ) | ( wire11605 ) | ( _23360 ) ;
 assign n_n4322 = ( n_n524  &  wire16  &  n_n535 ) ;
 assign wire11614 = ( n_n4372 ) | ( n_n4371 ) | ( n_n4361 ) | ( n_n4359 ) ;
 assign wire11618 = ( n_n3533 ) | ( n_n1308 ) | ( wire282 ) | ( wire11613 ) ;
 assign n_n1041 = ( n_n1120 ) | ( n_n3176 ) | ( wire11614 ) | ( wire11618 ) ;
 assign n_n4695 = ( n_n464  &  n_n390  &  wire23 ) ;
 assign n_n4826 = ( n_n532  &  wire17  &  n_n535 ) ;
 assign n_n5151 = ( n_n491  &  wire11  &  n_n130 ) ;
 assign wire773 = ( wire25  &  n_n464  &  n_n325 ) ;
 assign n_n4197 = ( n_n4811 ) | ( n_n4810 ) | ( wire773 ) ;
 assign wire330 = ( i_9_  &  n_n528  &  n_n260  &  n_n500 ) | ( (~ i_9_)  &  n_n528  &  n_n260  &  n_n500 ) ;
 assign n_n5071 = ( n_n464  &  wire11  &  n_n195 ) ;
 assign n_n1167 = ( n_n5100 ) | ( n_n5103 ) | ( n_n5102 ) ;
 assign wire14211 = ( n_n3285 ) | ( wire14208 ) | ( _26353 ) | ( _26354 ) ;
 assign n_n2997 = ( wire170 ) | ( n_n3152 ) | ( wire129 ) | ( _28000 ) ;
 assign n_n5198 = ( n_n464  &  n_n528  &  wire12 ) ;
 assign wire14615 = ( wire19  &  n_n526  &  n_n535 ) | ( wire19  &  n_n528  &  n_n535 ) ;
 assign n_n3037 = ( wire14615 ) | ( n_n65  &  wire11  &  n_n535 ) ;
 assign wire183 = ( n_n65  &  wire21  &  n_n535 ) | ( n_n65  &  n_n535  &  wire20 ) ;
 assign wire453 = ( wire25  &  n_n464  &  n_n130 ) | ( n_n464  &  wire24  &  n_n130 ) ;
 assign n_n5246 = ( wire19  &  n_n509  &  n_n528 ) ;
 assign n_n5176 = ( n_n473  &  n_n534  &  wire12 ) ;
 assign wire80 = ( n_n473  &  wire21  &  n_n390 ) | ( n_n473  &  n_n390  &  wire20 ) ;
 assign wire157 = ( i_9_  &  n_n473  &  n_n390  &  n_n530 ) | ( (~ i_9_)  &  n_n473  &  n_n390  &  n_n530 ) ;
 assign wire15239 = ( n_n5129 ) | ( n_n5124 ) | ( n_n5128 ) | ( n_n5122 ) ;
 assign n_n2579 = ( n_n5125 ) | ( n_n5126 ) | ( n_n2685 ) | ( wire15239 ) ;
 assign wire88 = ( n_n535  &  n_n520  &  wire12 ) ;
 assign wire15245 = ( n_n5096 ) | ( n_n5099 ) | ( wire15241 ) ;
 assign n_n2541 = ( n_n2579 ) | ( wire15247 ) | ( _27424 ) | ( _27425 ) ;
 assign wire297 = ( wire25  &  n_n491  &  n_n195 ) | ( wire15  &  n_n491  &  n_n195 ) ;
 assign wire394 = ( i_9_  &  n_n526  &  n_n195  &  n_n500 ) | ( (~ i_9_)  &  n_n526  &  n_n195  &  n_n500 ) ;
 assign wire15235 = ( wire15226 ) | ( wire15227 ) | ( wire15230 ) | ( wire15231 ) ;
 assign wire14838 = ( n_n4475 ) | ( n_n4476 ) | ( n_n4457 ) ;
 assign wire14839 = ( n_n4463 ) | ( n_n4494 ) | ( wire14836 ) ;
 assign wire14854 = ( n_n4673 ) | ( n_n4690 ) | ( n_n4692 ) ;
 assign wire14855 = ( n_n4656 ) | ( n_n4697 ) | ( n_n4681 ) | ( n_n4660 ) ;
 assign wire361 = ( i_9_  &  n_n482  &  n_n455  &  n_n530 ) | ( (~ i_9_)  &  n_n482  &  n_n455  &  n_n530 ) ;
 assign wire378 = ( i_9_  &  n_n482  &  n_n455  &  n_n528 ) | ( (~ i_9_)  &  n_n482  &  n_n455  &  n_n528 ) ;
 assign wire341 = ( i_9_  &  n_n518  &  n_n534  &  n_n195 ) | ( (~ i_9_)  &  n_n518  &  n_n534  &  n_n195 ) ;
 assign wire362 = ( n_n535  &  n_n195  &  wire20 ) | ( n_n535  &  n_n195  &  wire23 ) ;
 assign wire203 = ( i_9_  &  n_n65  &  n_n491  &  n_n534 ) | ( (~ i_9_)  &  n_n65  &  n_n491  &  n_n534 ) ;
 assign wire205 = ( i_9_  &  n_n65  &  n_n526  &  n_n500 ) | ( (~ i_9_)  &  n_n65  &  n_n526  &  n_n500 ) ;
 assign wire438 = ( i_9_  &  n_n65  &  n_n491  &  n_n530 ) | ( (~ i_9_)  &  n_n65  &  n_n491  &  n_n530 ) ;
 assign n_n4699 = ( wire24  &  n_n325  &  n_n535 ) ;
 assign n_n4687 = ( n_n464  &  wire11  &  n_n390 ) ;
 assign wire340 = ( n_n482  &  n_n526  &  wire17 ) | ( n_n482  &  n_n528  &  wire17 ) ;
 assign n_n5250 = ( wire19  &  n_n524  &  n_n509 ) ;
 assign n_n5205 = ( n_n464  &  wire20  &  n_n130 ) ;
 assign n_n801 = ( n_n5004 ) | ( n_n5003 ) | ( n_n5006 ) ;
 assign wire12255 = ( n_n522  &  wire18  &  n_n500 ) | ( n_n524  &  wire18  &  n_n500 ) ;
 assign wire12256 = ( wire21  &  n_n195  &  n_n500 ) | ( n_n195  &  wire20  &  n_n500 ) ;
 assign n_n1454 = ( n_n5008 ) | ( n_n801 ) | ( _1244 ) | ( _24270 ) ;
 assign wire12352 = ( n_n5241 ) | ( n_n5242 ) | ( n_n5246 ) ;
 assign wire12353 = ( n_n5240 ) | ( n_n5245 ) | ( wire320 ) ;
 assign n_n1436 = ( n_n5243 ) | ( n_n5235 ) | ( wire12352 ) | ( wire12353 ) ;
 assign n_n5330 = ( wire19  &  n_n524  &  n_n464 ) ;
 assign n_n5331 = ( n_n65  &  n_n464  &  wire21 ) ;
 assign wire421 = ( i_9_  &  n_n455  &  n_n532  &  n_n535 ) | ( (~ i_9_)  &  n_n455  &  n_n532  &  n_n535 ) ;
 assign wire225 = ( i_9_  &  n_n473  &  n_n390  &  n_n534 ) | ( (~ i_9_)  &  n_n473  &  n_n390  &  n_n534 ) ;
 assign wire11856 = ( i_9_  &  n_n482  &  n_n522  &  n_n390 ) | ( (~ i_9_)  &  n_n482  &  n_n522  &  n_n390 ) ;
 assign wire253 = ( i_9_  &  n_n482  &  n_n534  &  n_n195 ) | ( (~ i_9_)  &  n_n482  &  n_n534  &  n_n195 ) ;
 assign wire12009 = ( n_n5096 ) | ( n_n5099 ) | ( wire12007 ) ;
 assign n_n1061 = ( n_n5098 ) | ( n_n5105 ) | ( n_n1167 ) | ( wire12009 ) ;
 assign wire12014 = ( _22574 ) | ( _22575 ) ;
 assign wire12015 = ( n_n5078 ) | ( n_n5083 ) | ( wire232 ) | ( n_n5095 ) ;
 assign wire12020 = ( n_n5069 ) | ( n_n5066 ) | ( n_n4152 ) | ( wire12018 ) ;
 assign n_n1022 = ( n_n1061 ) | ( wire12014 ) | ( wire12015 ) | ( wire12020 ) ;
 assign wire104 = ( i_9_  &  n_n526  &  n_n509  &  n_n195 ) | ( (~ i_9_)  &  n_n526  &  n_n509  &  n_n195 ) ;
 assign wire12004 = ( wire11992 ) | ( wire11993 ) | ( wire11995 ) | ( wire11996 ) ;
 assign n_n4323 = ( wire21  &  n_n536  &  n_n535 ) ;
 assign wire128 = ( i_9_  &  n_n455  &  n_n535  &  n_n520 ) | ( (~ i_9_)  &  n_n455  &  n_n535  &  n_n520 ) ;
 assign n_n910 = ( n_n4434 ) | ( n_n4433 ) | ( n_n4435 ) ;
 assign n_n4631 = ( n_n390  &  wire23  &  n_n500 ) ;
 assign wire12595 = ( n_n4597 ) | ( n_n4601 ) | ( n_n4631 ) ;
 assign wire12596 = ( n_n4578 ) | ( n_n4611 ) | ( n_n4633 ) | ( n_n4581 ) ;
 assign n_n4761 = ( wire25  &  n_n491  &  n_n325 ) ;
 assign n_n4680 = ( n_n464  &  wire10  &  n_n534 ) ;
 assign wire343 = ( n_n522  &  wire18  &  n_n500 ) | ( n_n524  &  wire18  &  n_n500 ) ;
 assign wire379 = ( n_n482  &  n_n522  &  wire13 ) | ( n_n482  &  n_n524  &  wire13 ) ;
 assign wire15444 = ( n_n4535 ) | ( n_n4536 ) | ( n_n4529 ) ;
 assign wire15445 = ( n_n4526 ) | ( n_n4533 ) | ( wire379 ) ;
 assign n_n2996 = ( n_n4524 ) | ( n_n4537 ) | ( wire15444 ) | ( wire15445 ) ;
 assign wire431 = ( i_9_  &  n_n482  &  n_n390  &  n_n528 ) | ( (~ i_9_)  &  n_n482  &  n_n390  &  n_n528 ) ;
 assign n_n2670 = ( n_n5200 ) | ( n_n5199 ) | ( n_n5198 ) ;
 assign n_n4402 = ( n_n482  &  n_n524  &  wire16 ) ;
 assign wire238 = ( wire15  &  n_n390  &  n_n535 ) | ( wire11  &  n_n390  &  n_n535 ) ;
 assign wire276 = ( i_9_  &  n_n524  &  n_n390  &  n_n535 ) | ( (~ i_9_)  &  n_n524  &  n_n390  &  n_n535 ) ;
 assign n_n4702 = ( wire14  &  n_n528  &  n_n535 ) ;
 assign wire12159 = ( n_n4998 ) | ( wire104 ) | ( wire743 ) ;
 assign n_n4599 = ( n_n518  &  n_n390  &  wire23 ) ;
 assign wire364 = ( i_9_  &  n_n536  &  n_n535  &  n_n530 ) | ( (~ i_9_)  &  n_n536  &  n_n535  &  n_n530 ) ;
 assign n_n5283 = ( n_n65  &  n_n491  &  wire21 ) ;
 assign wire333 = ( i_9_  &  n_n65  &  n_n491  &  n_n532 ) | ( (~ i_9_)  &  n_n65  &  n_n491  &  n_n532 ) ;
 assign n_n4632 = ( n_n491  &  wire10  &  n_n534 ) ;
 assign wire139 = ( i_9_  &  n_n491  &  n_n390  &  n_n520 ) | ( (~ i_9_)  &  n_n491  &  n_n390  &  n_n520 ) ;
 assign wire11646 = ( n_n4671 ) | ( n_n4672 ) | ( n_n4723 ) ;
 assign wire11647 = ( n_n4667 ) | ( n_n4703 ) | ( n_n4658 ) | ( wire775 ) ;
 assign n_n953 = ( n_n4684 ) | ( n_n4708 ) | ( wire11646 ) | ( wire11647 ) ;
 assign wire99 = ( i_9_  &  n_n526  &  n_n390  &  n_n535 ) | ( (~ i_9_)  &  n_n526  &  n_n390  &  n_n535 ) ;
 assign wire11642 = ( n_n4633 ) | ( n_n4605 ) | ( n_n4632 ) | ( wire139 ) ;
 assign wire787 = ( wire22  &  n_n455  &  n_n509 ) ;
 assign wire13020 = ( n_n4470 ) | ( n_n4476 ) | ( n_n4472 ) ;
 assign n_n725 = ( wire184 ) | ( n_n901 ) | ( wire787 ) | ( wire13020 ) ;
 assign wire52 = ( i_9_  &  n_n518  &  n_n528  &  n_n260 ) | ( (~ i_9_)  &  n_n518  &  n_n528  &  n_n260 ) ;
 assign wire150 = ( wire22  &  n_n464  &  n_n325 ) | ( n_n464  &  n_n325  &  wire23 ) ;
 assign n_n4645 = ( n_n491  &  n_n390  &  wire20 ) ;
 assign wire310 = ( n_n491  &  wire22  &  n_n390 ) | ( n_n491  &  wire21  &  n_n390 ) ;
 assign n_n4696 = ( n_n534  &  wire14  &  n_n535 ) ;
 assign n_n4762 = ( n_n491  &  n_n532  &  wire14 ) ;
 assign n_n1952 = ( n_n5069 ) | ( n_n5070 ) | ( n_n5071 ) ;
 assign wire13512 = ( i_9_  &  n_n524  &  n_n536  &  n_n535 ) | ( (~ i_9_)  &  n_n524  &  n_n536  &  n_n535 ) ;
 assign wire407 = ( i_9_  &  n_n491  &  n_n532  &  n_n130 ) | ( (~ i_9_)  &  n_n491  &  n_n532  &  n_n130 ) ;
 assign wire13209 = ( n_n4930 ) | ( n_n4939 ) | ( wire180 ) | ( n_n4944 ) ;
 assign n_n4056 = ( wire13209 ) | ( _25638 ) | ( _25639 ) ;
 assign wire42 = ( i_9_  &  n_n473  &  n_n532  &  n_n260 ) | ( (~ i_9_)  &  n_n473  &  n_n532  &  n_n260 ) ;
 assign n_n814 = ( n_n4945 ) | ( n_n4946 ) | ( n_n4947 ) ;
 assign wire141 = ( n_n532  &  n_n535  &  wire18 ) | ( n_n534  &  n_n535  &  wire18 ) ;
 assign wire317 = ( n_n464  &  n_n260  &  wire20 ) | ( n_n464  &  n_n260  &  wire23 ) ;
 assign n_n5192 = ( n_n464  &  n_n534  &  wire12 ) ;
 assign wire106 = ( n_n536  &  n_n535  &  wire20 ) | ( n_n536  &  n_n535  &  wire23 ) ;
 assign wire375 = ( i_9_  &  n_n524  &  n_n518  &  n_n260 ) | ( (~ i_9_)  &  n_n524  &  n_n518  &  n_n260 ) ;
 assign n_n4558 = ( n_n464  &  wire13  &  n_n528 ) ;
 assign wire417 = ( i_9_  &  n_n473  &  n_n390  &  n_n520 ) | ( (~ i_9_)  &  n_n473  &  n_n390  &  n_n520 ) ;
 assign wire12449 = ( n_n491  &  wire16  &  n_n528 ) | ( n_n491  &  wire16  &  n_n530 ) ;
 assign wire27 = ( wire12449 ) | ( wire15  &  n_n491  &  n_n536 ) ;
 assign wire12207 = ( n_n4779 ) | ( n_n4780 ) | ( n_n4775 ) ;
 assign wire12208 = ( n_n4782 ) | ( n_n4781 ) | ( wire315 ) ;
 assign n_n1472 = ( n_n4778 ) | ( n_n4783 ) | ( wire12207 ) | ( wire12208 ) ;
 assign n_n763 = ( n_n5218 ) | ( n_n5217 ) | ( n_n5215 ) ;
 assign wire286 = ( wire21  &  n_n509  &  n_n130 ) | ( n_n509  &  wire20  &  n_n130 ) ;
 assign wire12871 = ( n_n5241 ) | ( n_n5234 ) | ( n_n5242 ) ;
 assign wire12872 = ( n_n5240 ) | ( n_n5238 ) | ( wire318 ) ;
 assign n_n667 = ( n_n5244 ) | ( n_n5243 ) | ( wire12871 ) | ( wire12872 ) ;
 assign wire12874 = ( i_9_  &  n_n65  &  n_n535  &  n_n520 ) | ( (~ i_9_)  &  n_n65  &  n_n535  &  n_n520 ) ;
 assign n_n761 = ( wire12874 ) | ( wire19  &  n_n518  &  n_n534 ) ;
 assign wire12876 = ( wire182 ) | ( wire19  &  n_n518  &  n_n532 ) ;
 assign wire12877 = ( n_n5228 ) | ( n_n5225 ) | ( wire183 ) ;
 assign wire12881 = ( n_n2291 ) | ( n_n763 ) | ( n_n761 ) | ( wire12875 ) ;
 assign n_n635 = ( n_n667 ) | ( wire12876 ) | ( wire12877 ) | ( wire12881 ) ;
 assign wire12884 = ( i_9_  &  n_n524  &  n_n130  &  n_n500 ) | ( (~ i_9_)  &  n_n524  &  n_n130  &  n_n500 ) ;
 assign n_n777 = ( wire12884 ) | ( n_n522  &  wire12  &  n_n500 ) ;
 assign n_n3772 = ( n_n5130 ) | ( n_n5131 ) | ( n_n5132 ) ;
 assign wire12894 = ( n_n5133 ) | ( n_n5153 ) | ( n_n5148 ) | ( wire12883 ) ;
 assign wire12898 = ( wire12888 ) | ( wire12889 ) | ( wire12892 ) | ( wire12893 ) ;
 assign n_n637 = ( n_n777 ) | ( n_n3772 ) | ( wire12894 ) | ( wire12898 ) ;
 assign n_n4559 = ( n_n464  &  n_n455  &  wire11 ) ;
 assign n_n5227 = ( n_n65  &  n_n518  &  wire24 ) ;
 assign n_n4694 = ( n_n464  &  wire10  &  n_n520 ) ;
 assign n_n4700 = ( wire14  &  n_n535  &  n_n530 ) ;
 assign n_n4219 = ( n_n4704 ) | ( n_n4703 ) | ( n_n4702 ) ;
 assign wire221 = ( i_9_  &  n_n532  &  n_n325  &  n_n535 ) | ( (~ i_9_)  &  n_n532  &  n_n325  &  n_n535 ) ;
 assign wire13244 = ( n_n4697 ) | ( n_n4695 ) | ( wire221 ) ;
 assign wire173 = ( i_9_  &  n_n518  &  n_n532  &  n_n325 ) | ( (~ i_9_)  &  n_n518  &  n_n532  &  n_n325 ) ;
 assign wire13246 = ( i_9_  &  n_n518  &  n_n325  &  n_n520 ) | ( (~ i_9_)  &  n_n518  &  n_n325  &  n_n520 ) ;
 assign wire13156 = ( n_n4821 ) | ( n_n4822 ) | ( n_n4823 ) ;
 assign wire12225 = ( i_9_  &  n_n464  &  n_n325  &  n_n530 ) | ( (~ i_9_)  &  n_n464  &  n_n325  &  n_n530 ) ;
 assign wire390 = ( n_n4820 ) | ( n_n4819 ) | ( wire85 ) | ( wire12225 ) ;
 assign wire13576 = ( n_n526  &  n_n518  &  wire12 ) | ( n_n526  &  wire12  &  n_n500 ) ;
 assign n_n3926 = ( n_n5144 ) | ( wire422 ) | ( wire13577 ) | ( _25931 ) ;
 assign wire13585 = ( n_n5240 ) | ( n_n5222 ) | ( n_n5227 ) ;
 assign wire13586 = ( n_n5236 ) | ( n_n5278 ) | ( n_n5260 ) | ( n_n5286 ) ;
 assign n_n3924 = ( n_n5219 ) | ( n_n5250 ) | ( wire13585 ) | ( wire13586 ) ;
 assign wire13592 = ( n_n5293 ) | ( n_n5296 ) | ( n_n5323 ) | ( n_n5311 ) ;
 assign n_n3923 = ( wire13592 ) | ( _25945 ) ;
 assign wire13598 = ( n_n4927 ) | ( n_n4958 ) | ( n_n4961 ) ;
 assign wire13599 = ( n_n4920 ) | ( n_n4987 ) | ( n_n4963 ) | ( n_n4974 ) ;
 assign n_n3928 = ( n_n4994 ) | ( n_n5009 ) | ( wire13598 ) | ( wire13599 ) ;
 assign wire13897 = ( n_n522  &  wire14  &  n_n535 ) | ( n_n524  &  wire14  &  n_n535 ) ;
 assign n_n2378 = ( n_n4704 ) | ( n_n4703 ) | ( n_n4705 ) ;
 assign n_n4693 = ( n_n464  &  n_n390  &  wire20 ) ;
 assign n_n3051 = ( n_n5129 ) | ( n_n5127 ) | ( n_n5126 ) ;
 assign wire15507 = ( n_n4389 ) | ( n_n4390 ) | ( wire420 ) ;
 assign wire15426 = ( n_n4448 ) | ( n_n4447 ) | ( wire421 ) ;
 assign n_n3003 = ( n_n4440 ) | ( wire470 ) | ( n_n4449 ) | ( wire15426 ) ;
 assign wire14917 = ( n_n4807 ) | ( n_n4808 ) | ( n_n4799 ) ;
 assign wire14918 = ( wire14914 ) | ( wire14915 ) ;
 assign n_n4910 = ( n_n482  &  n_n528  &  wire17 ) ;
 assign wire190 = ( wire22  &  n_n390  &  n_n500 ) | ( wire21  &  n_n390  &  n_n500 ) ;
 assign wire12458 = ( n_n4408 ) | ( n_n4405 ) | ( n_n4406 ) ;
 assign wire12459 = ( n_n4411 ) | ( n_n4412 ) | ( wire79 ) ;
 assign n_n1501 = ( n_n4403 ) | ( n_n4415 ) | ( wire12458 ) | ( wire12459 ) ;
 assign wire12465 = ( n_n4401 ) | ( n_n4396 ) | ( n_n4395 ) | ( n_n4402 ) ;
 assign n_n1426 = ( n_n1501 ) | ( wire12467 ) | ( _23478 ) | ( _23479 ) ;
 assign wire12316 = ( n_n5039 ) | ( wire356 ) | ( n_n5049 ) | ( n_n5052 ) ;
 assign n_n1409 = ( n_n1450 ) | ( wire12323 ) | ( _24226 ) | ( _24227 ) ;
 assign wire12332 = ( n_n5087 ) | ( n_n5088 ) | ( n_n5077 ) ;
 assign wire12333 = ( n_n5085 ) | ( n_n5082 ) | ( n_n5084 ) | ( n_n5079 ) ;
 assign n_n1448 = ( n_n5078 ) | ( n_n5083 ) | ( wire12332 ) | ( wire12333 ) ;
 assign wire12327 = ( n_n5112 ) | ( n_n5110 ) | ( wire414 ) ;
 assign wire12328 = ( n_n5108 ) | ( wire12326 ) | ( _24250 ) ;
 assign wire12340 = ( wire289 ) | ( wire12335 ) | ( wire12337 ) | ( _24258 ) ;
 assign n_n1408 = ( n_n1448 ) | ( wire12327 ) | ( wire12328 ) | ( wire12340 ) ;
 assign wire347 = ( wire15  &  n_n455  &  n_n500 ) | ( n_n455  &  wire11  &  n_n500 ) ;
 assign n_n789 = ( n_n5064 ) | ( n_n5063 ) | ( n_n5065 ) ;
 assign wire12902 = ( n_n5059 ) | ( n_n5073 ) | ( wire160 ) ;
 assign n_n680 = ( n_n5061 ) | ( n_n5058 ) | ( n_n789 ) | ( wire12902 ) ;
 assign wire12908 = ( n_n5057 ) | ( wire166 ) | ( n_n5047 ) | ( n_n5051 ) ;
 assign n_n639 = ( n_n680 ) | ( wire12914 ) | ( _24749 ) | ( _24750 ) ;
 assign wire12930 = ( wire12921 ) | ( wire12922 ) | ( wire12925 ) | ( wire12926 ) ;
 assign n_n625 = ( n_n639 ) | ( wire12946 ) | ( _24805 ) | ( _24806 ) ;
 assign n_n4548 = ( n_n473  &  n_n522  &  wire13 ) ;
 assign wire13531 = ( n_n4393 ) | ( n_n4390 ) | ( n_n4394 ) ;
 assign n_n4099 = ( wire425 ) | ( wire420 ) | ( wire13531 ) | ( _25322 ) ;
 assign wire13529 = ( n_n4416 ) | ( n_n4415 ) | ( n_n4414 ) | ( wire13526 ) ;
 assign wire445 = ( n_n464  &  wire21  &  n_n390 ) | ( n_n464  &  n_n390  &  wire20 ) ;
 assign wire422 = ( wire22  &  n_n130  &  n_n500 ) | ( wire21  &  n_n130  &  n_n500 ) ;
 assign wire442 = ( i_9_  &  n_n325  &  n_n535  &  n_n530 ) | ( (~ i_9_)  &  n_n325  &  n_n535  &  n_n530 ) ;
 assign wire386 = ( i_9_  &  n_n65  &  n_n522  &  n_n518 ) | ( (~ i_9_)  &  n_n65  &  n_n522  &  n_n518 ) ;
 assign wire789 = ( n_n491  &  n_n455  &  wire23 ) ;
 assign n_n3879 = ( n_n4518 ) | ( n_n4520 ) | ( wire789 ) ;
 assign n_n2058 = ( n_n4459 ) | ( n_n4456 ) | ( n_n4457 ) ;
 assign wire324 = ( i_9_  &  n_n534  &  n_n260  &  n_n500 ) | ( (~ i_9_)  &  n_n534  &  n_n260  &  n_n500 ) ;
 assign wire305 = ( i_9_  &  n_n482  &  n_n260  &  n_n530 ) | ( (~ i_9_)  &  n_n482  &  n_n260  &  n_n530 ) ;
 assign wire291 = ( wire15  &  n_n518  &  n_n455 ) | ( n_n518  &  n_n455  &  wire24 ) ;
 assign wire11507 = ( n_n4464 ) | ( n_n4463 ) | ( n_n4462 ) ;
 assign wire12682 = ( n_n4806 ) | ( n_n4805 ) | ( n_n4815 ) ;
 assign wire12683 = ( n_n4830 ) | ( n_n4800 ) | ( _25094 ) ;
 assign n_n554 = ( n_n4870 ) | ( n_n4819 ) | ( wire12682 ) | ( wire12683 ) ;
 assign wire279 = ( i_9_  &  n_n518  &  n_n534  &  n_n130 ) | ( (~ i_9_)  &  n_n518  &  n_n534  &  n_n130 ) ;
 assign wire13445 = ( n_n4612 ) | ( wire45 ) | ( n_n4609 ) ;
 assign wire13446 = ( wire108 ) | ( n_n4600 ) | ( wire13443 ) ;
 assign wire13452 = ( n_n4573 ) | ( wire239 ) | ( wire13448 ) | ( wire13450 ) ;
 assign wire401 = ( i_9_  &  n_n390  &  n_n528  &  n_n500 ) | ( (~ i_9_)  &  n_n390  &  n_n528  &  n_n500 ) ;
 assign wire14316 = ( n_n4744 ) | ( n_n4697 ) | ( n_n4721 ) ;
 assign wire14317 = ( n_n4717 ) | ( n_n4703 ) | ( n_n4736 ) | ( n_n4741 ) ;
 assign wire434 = ( n_n65  &  wire21  &  n_n509 ) | ( n_n65  &  n_n509  &  wire20 ) ;
 assign wire15511 = ( n_n4353 ) | ( n_n4358 ) | ( n_n4354 ) ;
 assign wire15512 = ( n_n4367 ) | ( n_n4368 ) | ( wire15509 ) ;
 assign n_n3009 = ( n_n4365 ) | ( n_n4356 ) | ( wire15511 ) | ( wire15512 ) ;
 assign wire11520 = ( i_9_  &  n_n522  &  n_n455  &  n_n535 ) | ( (~ i_9_)  &  n_n522  &  n_n455  &  n_n535 ) ;
 assign n_n3889 = ( wire11520 ) | ( wire13  &  n_n535  &  n_n520 ) ;
 assign wire16388 = ( n_n4725 ) | ( n_n4726 ) | ( n_n4729 ) ;
 assign wire16389 = ( wire244 ) | ( n_n4722 ) | ( n_n4721 ) ;
 assign n_n1677 = ( n_n4488 ) | ( n_n4487 ) | ( n_n4486 ) ;
 assign wire12493 = ( n_n4470 ) | ( n_n4469 ) | ( wire199 ) ;
 assign wire12234 = ( n_n4842 ) | ( n_n4851 ) | ( n_n4841 ) ;
 assign n_n1467 = ( wire52 ) | ( wire12234 ) | ( wire12232 ) | ( _24115 ) ;
 assign wire12231 = ( n_n4838 ) | ( n_n4833 ) | ( wire304 ) | ( wire735 ) ;
 assign wire11866 = ( n_n4718 ) | ( n_n4717 ) | ( n_n4716 ) ;
 assign wire11867 = ( n_n4711 ) | ( n_n4712 ) | ( wire173 ) ;
 assign n_n1091 = ( n_n4710 ) | ( n_n4719 ) | ( wire11866 ) | ( wire11867 ) ;
 assign wire13338 = ( n_n5258 ) | ( n_n5254 ) | ( wire434 ) ;
 assign wire124 = ( i_9_  &  n_n522  &  n_n518  &  n_n536 ) | ( (~ i_9_)  &  n_n522  &  n_n518  &  n_n536 ) ;
 assign wire12363 = ( wire149 ) | ( wire175 ) ;
 assign wire12364 = ( n_n5333 ) | ( n_n5330 ) | ( wire12361 ) ;
 assign wire12368 = ( n_n5314 ) | ( n_n5322 ) | ( wire115 ) ;
 assign wire12369 = ( n_n5318 ) | ( n_n5320 ) | ( n_n5312 ) | ( wire12366 ) ;
 assign n_n1402 = ( wire12363 ) | ( wire12364 ) | ( wire12368 ) | ( wire12369 ) ;
 assign wire12371 = ( i_9_  &  n_n65  &  n_n491  &  n_n528 ) | ( (~ i_9_)  &  n_n65  &  n_n491  &  n_n528 ) ;
 assign wire12372 = ( wire25  &  n_n65  &  n_n491 ) | ( n_n65  &  n_n491  &  wire24 ) ;
 assign wire204 = ( n_n5276 ) | ( n_n5277 ) | ( wire12371 ) | ( wire12372 ) ;
 assign wire11666 = ( n_n4518 ) | ( n_n4476 ) | ( n_n4500 ) ;
 assign wire11667 = ( n_n4477 ) | ( n_n4496 ) | ( n_n4505 ) | ( n_n4490 ) ;
 assign n_n956 = ( n_n4479 ) | ( n_n4468 ) | ( wire11666 ) | ( wire11667 ) ;
 assign n_n951 = ( n_n4832 ) | ( n_n4850 ) | ( wire11680 ) | ( wire11681 ) ;
 assign wire11675 = ( n_n4778 ) | ( n_n4801 ) | ( wire11671 ) ;
 assign wire11676 = ( n_n4773 ) | ( n_n4813 ) | ( n_n4742 ) | ( wire150 ) ;
 assign wire11690 = ( n_n4967 ) | ( n_n4986 ) | ( wire11687 ) | ( wire11688 ) ;
 assign n_n948 = ( n_n5075 ) | ( n_n5063 ) | ( wire11718 ) | ( wire11719 ) ;
 assign n_n949 = ( n_n5044 ) | ( n_n5011 ) | ( wire11725 ) | ( wire11726 ) ;
 assign wire11734 = ( wire11698 ) | ( wire11699 ) | ( wire11731 ) | ( wire11732 ) ;
 assign wire11735 = ( wire11705 ) | ( wire11706 ) | ( wire11712 ) | ( wire11713 ) ;
 assign wire13342 = ( n_n5244 ) | ( wire318 ) | ( n_n5243 ) ;
 assign wire600 = ( (~ i_9_)  &  (~ i_7_)  &  i_8_  &  (~ i_6_) ) | ( (~ i_9_)  &  i_7_  &  (~ i_8_)  &  (~ i_6_) ) ;
 assign n_n1478 = ( wire221 ) | ( wire12403 ) | ( wire12401 ) | ( _23753 ) ;
 assign n_n1476 = ( n_n4730 ) | ( n_n4722 ) | ( wire12408 ) | ( wire12409 ) ;
 assign wire12416 = ( n_n4715 ) | ( n_n4716 ) | ( wire12413 ) | ( wire12414 ) ;
 assign n_n5289 = ( wire25  &  n_n65  &  n_n482 ) ;
 assign wire255 = ( i_9_  &  n_n522  &  n_n518  &  n_n390 ) | ( (~ i_9_)  &  n_n522  &  n_n518  &  n_n390 ) ;
 assign n_n1727 = ( n_n4572 ) | ( n_n4518 ) | ( wire15822 ) | ( wire15823 ) ;
 assign wire15829 = ( n_n4641 ) | ( n_n4648 ) | ( n_n4651 ) | ( n_n4622 ) ;
 assign wire15830 = ( n_n4620 ) | ( n_n4627 ) | ( n_n4631 ) | ( wire255 ) ;
 assign n_n1712 = ( n_n1727 ) | ( wire15836 ) | ( wire15837 ) | ( _28538 ) ;
 assign wire15908 = ( n_n4420 ) | ( n_n4407 ) | ( n_n4412 ) ;
 assign wire15909 = ( n_n4373 ) | ( n_n4392 ) | ( n_n4426 ) | ( n_n4419 ) ;
 assign n_n1730 = ( n_n4394 ) | ( n_n4376 ) | ( wire15908 ) | ( wire15909 ) ;
 assign wire15914 = ( n_n4432 ) | ( n_n4468 ) | ( n_n4435 ) ;
 assign wire15915 = ( n_n4464 ) | ( n_n4455 ) | ( n_n4433 ) | ( n_n4441 ) ;
 assign n_n1729 = ( n_n4458 ) | ( n_n4451 ) | ( wire15914 ) | ( wire15915 ) ;
 assign n_n1725 = ( n_n4678 ) | ( n_n1764 ) | ( n_n4687 ) | ( wire15920 ) ;
 assign n_n1724 = ( n_n1760 ) | ( wire444 ) | ( wire15922 ) | ( _28546 ) ;
 assign wire15930 = ( n_n4784 ) | ( n_n4754 ) | ( wire15927 ) ;
 assign wire15931 = ( n_n4748 ) | ( n_n4772 ) | ( wire164 ) | ( n_n4766 ) ;
 assign n_n1711 = ( n_n1725 ) | ( n_n1724 ) | ( wire15930 ) | ( wire15931 ) ;
 assign n_n5282 = ( wire19  &  n_n491  &  n_n524 ) ;
 assign n_n5298 = ( n_n482  &  wire19  &  n_n524 ) ;
 assign wire13629 = ( n_n4724 ) | ( n_n4679 ) | ( n_n4686 ) ;
 assign wire13630 = ( n_n4663 ) | ( n_n4665 ) | ( n_n4672 ) | ( n_n4707 ) ;
 assign wire13635 = ( n_n4842 ) | ( n_n4867 ) | ( n_n4841 ) ;
 assign wire13636 = ( n_n4913 ) | ( n_n4903 ) | ( n_n4905 ) | ( n_n4846 ) ;
 assign wire261 = ( i_9_  &  n_n491  &  n_n534  &  n_n260 ) | ( (~ i_9_)  &  n_n491  &  n_n534  &  n_n260 ) ;
 assign n_n3694 = ( wire264 ) | ( n_n3810 ) | ( wire261 ) | ( _26964 ) ;
 assign n_n2761 = ( n_n4648 ) | ( n_n4647 ) | ( n_n4645 ) ;
 assign wire15750 = ( wire173 ) | ( wire15748 ) ;
 assign wire466 = ( n_n5155 ) | ( wire195 ) | ( n_n5160 ) | ( wire287 ) ;
 assign wire15605 = ( n_n5089 ) | ( n_n5098 ) | ( n_n5095 ) ;
 assign wire15606 = ( n_n5087 ) | ( n_n5088 ) | ( wire122 ) ;
 assign n_n2953 = ( n_n5091 ) | ( n_n5100 ) | ( wire15605 ) | ( wire15606 ) ;
 assign wire15609 = ( n_n5057 ) | ( n_n5058 ) | ( n_n5065 ) ;
 assign wire15610 = ( n_n5066 ) | ( n_n5063 ) | ( wire159 ) ;
 assign n_n2955 = ( n_n5072 ) | ( n_n5061 ) | ( wire15609 ) | ( wire15610 ) ;
 assign wire15616 = ( n_n5086 ) | ( n_n5073 ) | ( wire15612 ) ;
 assign wire15617 = ( n_n5079 ) | ( wire209 ) | ( wire15614 ) ;
 assign n_n2915 = ( n_n2953 ) | ( n_n2955 ) | ( wire15616 ) | ( wire15617 ) ;
 assign wire265 = ( i_9_  &  n_n526  &  n_n491  &  n_n195 ) | ( (~ i_9_)  &  n_n526  &  n_n491  &  n_n195 ) ;
 assign wire15633 = ( n_n3772 ) | ( n_n3051 ) | ( wire15626 ) | ( wire15627 ) ;
 assign wire15634 = ( wire15623 ) | ( wire15624 ) | ( wire15628 ) | ( wire15629 ) ;
 assign wire15642 = ( n_n2956 ) | ( wire15639 ) | ( _28238 ) | ( _28239 ) ;
 assign n_n2902 = ( n_n2915 ) | ( wire15633 ) | ( wire15634 ) | ( wire15642 ) ;
 assign wire15405 = ( n_n4757 ) | ( n_n4760 ) | ( n_n4815 ) ;
 assign wire15406 = ( n_n4769 ) | ( n_n4794 ) | ( n_n4797 ) | ( n_n4788 ) ;
 assign wire15069 = ( n_n4464 ) | ( n_n4471 ) | ( n_n4472 ) | ( n_n4469 ) ;
 assign n_n1840 = ( wire123 ) | ( wire209 ) | ( n_n1952 ) | ( _28607 ) ;
 assign wire15950 = ( wire279 ) | ( wire15947 ) ;
 assign wire15951 = ( n_n5089 ) | ( n_n5086 ) | ( n_n5088 ) | ( wire232 ) ;
 assign wire15957 = ( wire160 ) | ( wire15952 ) | ( wire15954 ) | ( _28618 ) ;
 assign n_n1801 = ( n_n1840 ) | ( wire15950 ) | ( wire15951 ) | ( wire15957 ) ;
 assign wire15961 = ( n_n5118 ) | ( n_n5121 ) | ( n_n5122 ) ;
 assign wire15962 = ( n_n5123 ) | ( n_n5114 ) | ( wire336 ) ;
 assign n_n1837 = ( n_n5115 ) | ( n_n5128 ) | ( wire15961 ) | ( wire15962 ) ;
 assign wire15968 = ( n_n5113 ) | ( n_n5104 ) | ( n_n5106 ) | ( wire122 ) ;
 assign n_n1800 = ( n_n1837 ) | ( wire15972 ) | ( _28636 ) | ( _28637 ) ;
 assign wire15977 = ( n_n5048 ) | ( n_n5047 ) | ( n_n5044 ) ;
 assign n_n1842 = ( wire97 ) | ( wire15977 ) | ( wire15975 ) | ( _28642 ) ;
 assign wire15920 = ( n_n4676 ) | ( n_n4655 ) | ( wire391 ) ;
 assign wire12783 = ( n_n4705 ) | ( n_n4706 ) | ( n_n4713 ) ;
 assign wire12784 = ( n_n4711 ) | ( n_n4712 ) | ( n_n4710 ) | ( n_n4709 ) ;
 assign n_n707 = ( n_n4708 ) | ( n_n4707 ) | ( wire12783 ) | ( wire12784 ) ;
 assign n_n691 = ( wire249 ) | ( wire42 ) | ( _1152 ) | ( _24602 ) ;
 assign wire12966 = ( n_n5327 ) | ( n_n5328 ) | ( wire149 ) | ( wire12963 ) ;
 assign wire12967 = ( wire148 ) | ( n_n5322 ) | ( wire11946 ) | ( wire175 ) ;
 assign n_n632 = ( wire12966 ) | ( wire12967 ) ;
 assign n_n700 = ( n_n4808 ) | ( n_n4799 ) | ( wire12756 ) | ( wire12757 ) ;
 assign wire12762 = ( n_n4782 ) | ( n_n4781 ) | ( wire12759 ) ;
 assign n_n646 = ( n_n700 ) | ( wire12766 ) | ( _24485 ) | ( _24486 ) ;
 assign wire12753 = ( wire12742 ) | ( wire12743 ) | ( wire12747 ) | ( wire12748 ) ;
 assign n_n627 = ( n_n646 ) | ( wire12774 ) | ( _24526 ) | ( _24527 ) ;
 assign wire683 = ( wire24  &  n_n509  &  n_n325 ) ;
 assign n_n856 = ( n_n4734 ) | ( n_n4729 ) | ( wire683 ) ;
 assign wire12790 = ( n_n4720 ) | ( n_n4728 ) | ( wire12787 ) ;
 assign wire12791 = ( n_n4725 ) | ( n_n4726 ) | ( n_n4721 ) | ( wire12788 ) ;
 assign wire12796 = ( n_n3849 ) | ( n_n4702 ) | ( n_n4694 ) | ( wire12794 ) ;
 assign n_n648 = ( n_n707 ) | ( wire12790 ) | ( wire12791 ) | ( wire12796 ) ;
 assign wire12814 = ( wire12799 ) | ( wire12800 ) | ( wire12804 ) | ( wire12805 ) ;
 assign n_n628 = ( n_n648 ) | ( wire12826 ) | ( _24594 ) | ( _24595 ) ;
 assign wire12865 = ( n_n691 ) | ( wire12862 ) | ( _24620 ) | ( _24621 ) ;
 assign wire12866 = ( wire12843 ) | ( wire12844 ) | ( wire12857 ) | ( wire12858 ) ;
 assign n_n1760 = ( n_n4738 ) | ( n_n4733 ) | ( n_n4736 ) ;
 assign wire15333 = ( n_n4634 ) | ( n_n4687 ) | ( n_n4631 ) ;
 assign wire15334 = ( n_n4659 ) | ( wire75 ) | ( n_n4689 ) | ( n_n4698 ) ;
 assign wire53 = ( i_9_  &  n_n524  &  n_n518  &  n_n536 ) | ( (~ i_9_)  &  n_n524  &  n_n518  &  n_n536 ) ;
 assign wire16159 = ( n_n473  &  n_n526  &  wire17 ) | ( n_n473  &  n_n534  &  wire17 ) ;
 assign n_n1852 = ( wire249 ) | ( n_n4932 ) | ( wire42 ) | ( wire16159 ) ;
 assign wire16164 = ( n_n4940 ) | ( n_n4939 ) | ( wire180 ) ;
 assign wire16165 = ( n_n4937 ) | ( n_n4938 ) | ( wire305 ) ;
 assign wire16168 = ( n_n4919 ) | ( n_n4910 ) | ( wire13870 ) | ( wire16166 ) ;
 assign n_n1805 = ( n_n1852 ) | ( wire16164 ) | ( wire16165 ) | ( wire16168 ) ;
 assign wire16158 = ( wire16148 ) | ( wire16149 ) | ( wire16152 ) | ( wire16153 ) ;
 assign wire444 = ( n_n526  &  n_n464  &  wire10 ) | ( n_n524  &  n_n464  &  wire10 ) ;
 assign wire12403 = ( n_n4695 ) | ( n_n4696 ) | ( n_n4700 ) ;
 assign wire12969 = ( n_n5303 ) | ( n_n5304 ) | ( wire63 ) ;
 assign wire12970 = ( n_n5307 ) | ( n_n5308 ) | ( n_n5309 ) ;
 assign n_n662 = ( n_n5302 ) | ( n_n5306 ) | ( wire12969 ) | ( wire12970 ) ;
 assign wire12971 = ( n_n473  &  wire19  &  n_n526 ) | ( n_n473  &  wire19  &  n_n522 ) ;
 assign wire12975 = ( n_n5318 ) | ( n_n5320 ) | ( n_n5315 ) | ( wire12972 ) ;
 assign n_n661 = ( wire269 ) | ( wire12971 ) | ( wire12975 ) ;
 assign wire13001 = ( wire12984 ) | ( wire12998 ) | ( _24885 ) | ( _24886 ) ;
 assign wire14470 = ( n_n4372 ) | ( n_n4371 ) | ( n_n4376 ) ;
 assign wire14471 = ( n_n4367 ) | ( n_n4368 ) | ( wire14468 ) ;
 assign n_n3736 = ( n_n4366 ) | ( n_n4375 ) | ( wire14470 ) | ( wire14471 ) ;
 assign wire15348 = ( n_n4898 ) | ( n_n4877 ) | ( n_n4876 ) | ( n_n4899 ) ;
 assign wire15349 = ( n_n4886 ) | ( n_n4915 ) | ( wire154 ) | ( n_n4874 ) ;
 assign wire15008 = ( n_n4705 ) | ( n_n4706 ) | ( wire15007 ) ;
 assign wire13055 = ( wire16  &  n_n528  &  n_n500 ) | ( wire16  &  n_n500  &  n_n530 ) ;
 assign wire16188 = ( n_n4803 ) | ( n_n4804 ) | ( n_n4799 ) ;
 assign wire16189 = ( n_n4807 ) | ( n_n4808 ) | ( wire16186 ) ;
 assign n_n1862 = ( n_n4802 ) | ( n_n4805 ) | ( wire16188 ) | ( wire16189 ) ;
 assign wire16193 = ( _28370 ) | ( n_n464  &  wire11  &  n_n325 ) ;
 assign wire16194 = ( n_n4834 ) | ( n_n4833 ) | ( wire150 ) ;
 assign wire16198 = ( wire388 ) | ( n_n4197 ) | ( wire16195 ) ;
 assign n_n1808 = ( n_n1862 ) | ( wire16193 ) | ( wire16194 ) | ( wire16198 ) ;
 assign wire16217 = ( n_n4882 ) | ( n_n4881 ) | ( wire16215 ) ;
 assign n_n1856 = ( n_n4876 ) | ( wire461 ) | ( n_n4875 ) | ( wire16217 ) ;
 assign wire16213 = ( wire176 ) | ( n_n4841 ) | ( wire16211 ) | ( _28382 ) ;
 assign wire16214 = ( wire16203 ) | ( wire16204 ) | ( wire16206 ) | ( wire16207 ) ;
 assign wire16224 = ( n_n1856 ) | ( wire16184 ) | ( wire16185 ) | ( wire16222 ) ;
 assign wire15822 = ( n_n4593 ) | ( n_n4594 ) | ( n_n4552 ) ;
 assign wire15823 = ( n_n4511 ) | ( n_n4590 ) | ( wire15819 ) ;
 assign wire15851 = ( n_n4849 ) | ( n_n4790 ) | ( n_n4813 ) ;
 assign wire15852 = ( n_n4821 ) | ( n_n4842 ) | ( wire15848 ) ;
 assign n_n1722 = ( n_n4801 ) | ( n_n4820 ) | ( wire15851 ) | ( wire15852 ) ;
 assign wire15858 = ( n_n4887 ) | ( n_n4930 ) | ( n_n4929 ) ;
 assign wire15859 = ( n_n4912 ) | ( n_n4968 ) | ( n_n4967 ) | ( n_n4899 ) ;
 assign n_n1721 = ( n_n4915 ) | ( n_n4961 ) | ( wire15858 ) | ( wire15859 ) ;
 assign wire13028 = ( wire15  &  n_n491  &  n_n455 ) | ( n_n491  &  n_n455  &  wire24 ) ;
 assign n_n722 = ( n_n4247 ) | ( wire308 ) | ( _1050 ) | ( _24893 ) ;
 assign wire13034 = ( n_n4502 ) | ( n_n4501 ) | ( wire378 ) ;
 assign wire13035 = ( n_n4521 ) | ( n_n4504 ) | ( n_n4524 ) | ( n_n4503 ) ;
 assign wire13039 = ( n_n4498 ) | ( n_n3879 ) | ( wire13027 ) | ( wire13036 ) ;
 assign n_n653 = ( n_n722 ) | ( wire13034 ) | ( wire13035 ) | ( wire13039 ) ;
 assign wire13016 = ( n_n4421 ) | ( wire215 ) | ( n_n910 ) | ( wire13013 ) ;
 assign wire13017 = ( wire13005 ) | ( wire13006 ) | ( wire13015 ) ;
 assign wire13046 = ( n_n725 ) | ( wire13025 ) | ( wire13026 ) | ( wire13044 ) ;
 assign n_n630 = ( n_n653 ) | ( wire13016 ) | ( wire13017 ) | ( wire13046 ) ;
 assign wire14544 = ( n_n5279 ) | ( n_n5270 ) | ( n_n5280 ) ;
 assign n_n3664 = ( wire203 ) | ( wire438 ) | ( wire14544 ) | ( _27142 ) ;
 assign wire15521 = ( n_n4325 ) | ( n_n4314 ) | ( n_n4328 ) ;
 assign n_n3012 = ( n_n4317 ) | ( n_n4326 ) | ( wire363 ) | ( wire15521 ) ;
 assign wire15517 = ( n_n4344 ) | ( n_n4342 ) | ( wire124 ) ;
 assign wire15769 = ( n_n4683 ) | ( n_n4678 ) | ( n_n4684 ) ;
 assign wire15770 = ( n_n4671 ) | ( n_n4672 ) | ( wire80 ) ;
 assign n_n2985 = ( n_n4674 ) | ( n_n4681 ) | ( wire15769 ) | ( wire15770 ) ;
 assign wire15774 = ( wire444 ) | ( n_n464  &  n_n390  &  wire20 ) ;
 assign wire15775 = ( n_n4712 ) | ( n_n4685 ) | ( wire15773 ) ;
 assign wire15778 = ( n_n4710 ) | ( n_n4709 ) | ( n_n4219 ) | ( wire15776 ) ;
 assign n_n2925 = ( n_n2985 ) | ( wire15774 ) | ( wire15775 ) | ( wire15778 ) ;
 assign n_n2832 = ( n_n5140 ) | ( n_n5144 ) | ( wire15354 ) | ( wire15355 ) ;
 assign n_n2834 = ( n_n5033 ) | ( n_n4989 ) | ( wire15360 ) | ( wire15361 ) ;
 assign wire15367 = ( n_n5092 ) | ( n_n5069 ) | ( n_n5084 ) | ( n_n5078 ) ;
 assign wire15368 = ( n_n5068 ) | ( n_n5080 ) | ( n_n5090 ) | ( wire279 ) ;
 assign wire15389 = ( n_n4959 ) | ( n_n4960 ) | ( n_n4961 ) ;
 assign wire15390 = ( n_n4963 ) | ( n_n4964 ) | ( n_n4974 ) | ( n_n4967 ) ;
 assign wire16099 = ( n_n4389 ) | ( n_n4388 ) | ( n_n4393 ) | ( n_n4390 ) ;
 assign wire16094 = ( n_n4430 ) | ( n_n4416 ) | ( wire37 ) ;
 assign wire16105 = ( n_n4403 ) | ( n_n4400 ) | ( wire16102 ) | ( wire16103 ) ;
 assign wire16233 = ( n_n4760 ) | ( n_n4767 ) | ( _28413 ) ;
 assign wire12408 = ( n_n4725 ) | ( n_n4726 ) | ( n_n4721 ) ;
 assign wire12409 = ( n_n4720 ) | ( n_n4727 ) | ( n_n4729 ) | ( n_n4719 ) ;
 assign wire13073 = ( n_n4389 ) | ( n_n4390 ) | ( n_n4394 ) ;
 assign wire13074 = ( n_n4383 ) | ( n_n4388 ) | ( n_n4396 ) | ( n_n4395 ) ;
 assign n_n732 = ( n_n4393 ) | ( n_n4386 ) | ( wire13073 ) | ( wire13074 ) ;
 assign wire13070 = ( n_n4416 ) | ( n_n4415 ) | ( n_n4414 ) | ( wire13067 ) ;
 assign n_n656 = ( n_n732 ) | ( wire13078 ) | ( _24973 ) | ( _24974 ) ;
 assign wire13066 = ( wire27 ) | ( wire13059 ) | ( wire13060 ) | ( wire13062 ) ;
 assign n_n631 = ( n_n656 ) | ( wire13087 ) | ( _25017 ) | ( _25018 ) ;
 assign n_n715 = ( n_n4603 ) | ( n_n4591 ) | ( wire13100 ) | ( wire13101 ) ;
 assign wire13106 = ( n_n4584 ) | ( n_n4583 ) | ( wire238 ) ;
 assign wire13107 = ( n_n4568 ) | ( wire783 ) | ( wire99 ) ;
 assign wire13111 = ( n_n881 ) | ( wire13105 ) | ( wire13108 ) ;
 assign n_n651 = ( n_n715 ) | ( wire13106 ) | ( wire13107 ) | ( wire13111 ) ;
 assign wire13124 = ( wire13113 ) | ( wire13114 ) | ( wire13118 ) | ( wire13119 ) ;
 assign n_n629 = ( n_n651 ) | ( wire13132 ) | ( _25084 ) | ( _25085 ) ;
 assign wire14322 = ( n_n4658 ) | ( n_n4687 ) | ( wire775 ) ;
 assign wire14323 = ( n_n4646 ) | ( n_n4668 ) | ( wire14320 ) ;
 assign wire15653 = ( n_n5279 ) | ( n_n5280 ) | ( n_n5283 ) ;
 assign n_n2939 = ( wire333 ) | ( wire15653 ) | ( wire15651 ) | ( _28305 ) ;
 assign wire15354 = ( n_n5111 ) | ( n_n5113 ) | ( n_n5143 ) ;
 assign wire15355 = ( n_n5161 ) | ( n_n5120 ) | ( n_n5135 ) | ( n_n5147 ) ;
 assign wire15360 = ( n_n5064 ) | ( n_n5001 ) | ( wire755 ) ;
 assign wire15361 = ( n_n4990 ) | ( n_n5027 ) | ( n_n5048 ) | ( n_n5053 ) ;
 assign wire11873 = ( n_n4704 ) | ( n_n4697 ) | ( wire11870 ) ;
 assign wire11874 = ( n_n4707 ) | ( n_n4702 ) | ( n_n4700 ) | ( wire221 ) ;
 assign n_n1032 = ( n_n1093 ) | ( n_n1091 ) | ( wire11873 ) | ( wire11874 ) ;
 assign wire11718 = ( n_n5093 ) | ( n_n5054 ) | ( n_n5068 ) ;
 assign wire11719 = ( n_n5106 ) | ( n_n5070 ) | ( wire11715 ) ;
 assign wire12756 = ( n_n4803 ) | ( n_n4804 ) | ( wire686 ) ;
 assign wire12757 = ( n_n4811 ) | ( n_n4801 ) | ( n_n4802 ) | ( n_n4807 ) ;
 assign wire14752 = ( i_9_  &  n_n532  &  n_n535  &  n_n195 ) | ( (~ i_9_)  &  n_n532  &  n_n535  &  n_n195 ) ;
 assign wire14754 = ( n_n4959 ) | ( n_n4962 ) | ( n_n4961 ) ;
 assign n_n3689 = ( n_n3803 ) | ( n_n4953 ) | ( wire14752 ) | ( wire14754 ) ;
 assign wire14448 = ( n_n4515 ) | ( wire791 ) | ( wire14446 ) ;
 assign wire11725 = ( n_n5040 ) | ( n_n4999 ) | ( n_n5024 ) ;
 assign wire11726 = ( n_n5025 ) | ( n_n5049 ) | ( n_n5047 ) | ( n_n5051 ) ;
 assign wire13100 = ( n_n4595 ) | ( n_n4596 ) | ( n_n4599 ) ;
 assign wire13101 = ( n_n4598 ) | ( n_n4593 ) | ( n_n4594 ) | ( n_n4600 ) ;
 assign wire14618 = ( n_n5201 ) | ( n_n5192 ) | ( wire761 ) ;
 assign wire14619 = ( n_n5200 ) | ( n_n5193 ) | ( wire452 ) ;
 assign n_n3670 = ( n_n5199 ) | ( n_n5194 ) | ( wire14618 ) | ( wire14619 ) ;
 assign wire15663 = ( n_n5300 ) | ( n_n5299 ) | ( wire15660 ) ;
 assign n_n2937 = ( n_n5303 ) | ( n_n3019 ) | ( n_n5313 ) | ( wire15663 ) ;
 assign wire15451 = ( n_n4547 ) | ( n_n4544 ) | ( wire15448 ) ;
 assign wire15452 = ( n_n4550 ) | ( n_n4545 ) | ( wire201 ) | ( n_n4549 ) ;
 assign wire15870 = ( n_n5111 ) | ( n_n5081 ) | ( n_n5080 ) ;
 assign wire15871 = ( n_n5098 ) | ( n_n5087 ) | ( n_n5116 ) | ( n_n5102 ) ;
 assign n_n1718 = ( n_n5078 ) | ( n_n5108 ) | ( wire15870 ) | ( wire15871 ) ;
 assign wire15875 = ( n_n473  &  n_n522  &  wire12 ) | ( n_n473  &  n_n520  &  wire12 ) ;
 assign n_n1717 = ( n_n5138 ) | ( wire15873 ) | ( wire15876 ) | ( _28496 ) ;
 assign wire11680 = ( n_n4834 ) | ( n_n4844 ) | ( n_n4833 ) ;
 assign wire11681 = ( n_n4857 ) | ( n_n4847 ) | ( wire11677 ) ;
 assign wire16300 = ( _28574 ) | ( _28575 ) ;
 assign wire16305 = ( n_n5275 ) | ( n_n5271 ) | ( n_n5264 ) | ( wire77 ) ;
 assign wire15995 = ( n_n4488 ) | ( n_n4489 ) | ( n_n4490 ) | ( wire15993 ) ;
 assign wire14438 = ( wire21  &  n_n455  &  n_n509 ) | ( n_n455  &  n_n509  &  wire23 ) ;
 assign wire16034 = ( n_n4570 ) | ( n_n4569 ) | ( wire266 ) ;
 assign n_n1879 = ( wire99 ) | ( wire16034 ) | ( wire16032 ) | ( _28741 ) ;
 assign wire16040 = ( _28709 ) | ( wire22  &  n_n390  &  n_n509 ) ;
 assign wire16041 = ( wire465 ) | ( wire12519 ) | ( _28710 ) ;
 assign wire16048 = ( n_n4626 ) | ( n_n4625 ) | ( wire16045 ) | ( wire16046 ) ;
 assign n_n1872 = ( n_n4674 ) | ( n_n4661 ) | ( wire16052 ) | ( wire16053 ) ;
 assign wire16059 = ( n_n4646 ) | ( n_n4659 ) | ( wire16056 ) ;
 assign wire11852 = ( wire11841 ) | ( wire11842 ) | ( wire11846 ) | ( wire11847 ) ;
 assign wire14517 = ( n_n4455 ) | ( n_n4456 ) | ( n_n4457 ) | ( n_n4462 ) ;
 assign n_n3699 = ( n_n3820 ) | ( _26878 ) | ( _26879 ) | ( _26880 ) ;
 assign wire14701 = ( n_n4806 ) | ( n_n4805 ) | ( n_n4808 ) ;
 assign wire14702 = ( n_n4804 ) | ( n_n4815 ) | ( _26883 ) ;
 assign n_n3701 = ( n_n4810 ) | ( n_n4813 ) | ( wire14701 ) | ( wire14702 ) ;
 assign wire14708 = ( n_n4817 ) | ( n_n4828 ) | ( n_n4823 ) | ( n_n4820 ) ;
 assign wire14709 = ( n_n4821 ) | ( n_n4822 ) | ( n_n4826 ) | ( wire14706 ) ;
 assign n_n3645 = ( n_n3699 ) | ( n_n3701 ) | ( wire14708 ) | ( wire14709 ) ;
 assign wire16052 = ( n_n4669 ) | ( n_n4670 ) | ( n_n4665 ) ;
 assign wire16053 = ( n_n4666 ) | ( n_n4662 ) | ( n_n4671 ) | ( n_n4672 ) ;
 assign wire16266 = ( n_n5239 ) | ( n_n5240 ) | ( n_n5246 ) ;
 assign wire16267 = ( n_n5244 ) | ( n_n5241 ) | ( wire386 ) ;
 assign n_n1828 = ( n_n5234 ) | ( n_n5242 ) | ( wire16266 ) | ( wire16267 ) ;
 assign wire16272 = ( n_n5228 ) | ( n_n5220 ) | ( wire182 ) ;
 assign wire14723 = ( wire14714 ) | ( wire14715 ) | ( wire14718 ) | ( wire14719 ) ;
 assign wire14624 = ( n_n5189 ) | ( n_n5190 ) | ( n_n5203 ) ;
 assign wire14625 = ( wire14621 ) | ( wire14622 ) ;
 assign wire14629 = ( n_n4129 ) | ( n_n1532 ) | ( n_n3037 ) | ( wire14623 ) ;
 assign wire14760 = ( n_n4983 ) | ( n_n4984 ) | ( n_n4972 ) ;
 assign wire14761 = ( n_n4981 ) | ( n_n4987 ) | ( wire14756 ) ;
 assign wire14764 = ( n_n4965 ) | ( wire13215 ) | ( wire13836 ) | ( wire14762 ) ;
 assign wire15766 = ( n_n4771 ) | ( wire11748 ) | ( _27835 ) ;
 assign wire15767 = ( wire15756 ) | ( wire15757 ) | ( wire15760 ) | ( wire15761 ) ;
 assign wire15786 = ( wire15750 ) | ( wire15784 ) | ( _27854 ) | ( _27861 ) ;
 assign wire266 = ( n_n464  &  n_n455  &  wire23 ) ;
 assign wire606 = ( n_n522  &  n_n491  &  wire13 ) ;
 assign wire617 = ( n_n455  &  n_n509  &  wire20 ) ;
 assign wire636 = ( n_n524  &  n_n464  &  wire12 ) ;
 assign wire656 = ( n_n65  &  n_n482  &  wire20 ) ;
 assign wire669 = ( n_n473  &  n_n520  &  wire18 ) ;
 assign wire671 = ( n_n522  &  n_n464  &  wire13 ) ;
 assign wire675 = ( wire16  &  n_n532  &  n_n509 ) ;
 assign wire677 = ( wire15  &  n_n518  &  n_n536 ) ;
 assign wire679 = ( wire20  &  n_n130  &  n_n500 ) ;
 assign wire686 = ( wire25  &  n_n464  &  n_n325 ) ;
 assign wire695 = ( n_n491  &  n_n520  &  wire18 ) ;
 assign wire706 = ( n_n518  &  n_n532  &  wire18 ) ;
 assign wire724 = ( n_n482  &  n_n524  &  wire13 ) ;
 assign wire735 = ( wire15  &  n_n535  &  n_n260 ) ;
 assign wire743 = ( n_n509  &  n_n195  &  wire20 ) ;
 assign wire745 = ( n_n491  &  wire10  &  n_n530 ) ;
 assign wire755 = ( n_n473  &  n_n520  &  wire18 ) ;
 assign wire761 = ( n_n524  &  n_n464  &  wire12 ) ;
 assign wire765 = ( n_n473  &  wire12  &  n_n530 ) ;
 assign wire767 = ( wire24  &  n_n509  &  n_n325 ) ;
 assign wire771 = ( wire25  &  n_n518  &  n_n195 ) ;
 assign wire772 = ( n_n518  &  n_n532  &  wire18 ) ;
 assign wire775 = ( wire15  &  n_n482  &  n_n390 ) ;
 assign wire11482 = ( n_n4432 ) | ( n_n4435 ) | ( wire421 ) ;
 assign wire11483 = ( n_n4440 ) | ( n_n4434 ) | ( wire236 ) | ( n_n4438 ) ;
 assign wire11488 = ( n_n491  &  n_n524  &  wire13 ) | ( n_n491  &  wire13  &  n_n532 ) ;
 assign wire11489 = ( wire15  &  n_n491  &  n_n455 ) | ( n_n491  &  n_n455  &  wire24 ) ;
 assign wire11491 = ( wire308 ) | ( wire11488 ) ;
 assign wire11492 = ( n_n4508 ) | ( wire129 ) | ( wire11489 ) ;
 assign wire11495 = ( n_n4515 ) | ( wire791 ) | ( n_n4492 ) ;
 assign wire11496 = ( wire65 ) | ( n_n4520 ) | ( wire789 ) ;
 assign wire11497 = ( n_n4502 ) | ( n_n4501 ) | ( wire347 ) ;
 assign wire11498 = ( n_n4521 ) | ( n_n4504 ) | ( n_n4517 ) | ( n_n4497 ) ;
 assign wire11505 = ( i_9_  &  n_n524  &  n_n518  &  n_n455 ) | ( (~ i_9_)  &  n_n524  &  n_n518  &  n_n455 ) ;
 assign wire11513 = ( wire25  &  n_n455  &  n_n509 ) | ( n_n455  &  n_n509  &  wire23 ) ;
 assign wire11515 = ( n_n4470 ) | ( n_n4475 ) | ( n_n4469 ) ;
 assign wire11516 = ( n_n4471 ) | ( n_n4472 ) | ( wire11513 ) ;
 assign wire11521 = ( n_n526  &  wire13  &  n_n535 ) | ( n_n524  &  wire13  &  n_n535 ) ;
 assign wire11522 = ( n_n4445 ) | ( wire368 ) | ( n_n4446 ) ;
 assign wire11523 = ( n_n4454 ) | ( wire11520 ) | ( wire11521 ) ;
 assign wire11524 = ( n_n473  &  n_n536  &  wire20 ) | ( n_n473  &  n_n536  &  wire23 ) ;
 assign wire11527 = ( wire37 ) | ( n_n4428 ) | ( wire11524 ) ;
 assign wire11529 = ( wire11482 ) | ( wire11483 ) | ( wire11522 ) | ( wire11523 ) ;
 assign wire11532 = ( i_9_  &  n_n473  &  n_n455  &  n_n532 ) | ( (~ i_9_)  &  n_n473  &  n_n455  &  n_n532 ) ;
 assign wire11534 = ( n_n473  &  wire22  &  n_n455 ) | ( n_n473  &  n_n455  &  wire11 ) ;
 assign wire11535 = ( n_n473  &  n_n455  &  wire20 ) | ( n_n473  &  n_n455  &  wire23 ) ;
 assign wire11536 = ( n_n4547 ) | ( n_n4544 ) | ( wire11534 ) ;
 assign wire11539 = ( wire15  &  n_n464  &  n_n455 ) | ( wire22  &  n_n464  &  n_n455 ) ;
 assign wire11547 = ( i_9_  &  n_n532  &  n_n390  &  n_n500 ) | ( (~ i_9_)  &  n_n532  &  n_n390  &  n_n500 ) ;
 assign wire11548 = ( n_n4617 ) | ( n_n4613 ) | ( n_n4612 ) | ( n_n4611 ) ;
 assign wire11549 = ( n_n4616 ) | ( wire465 ) | ( wire11547 ) ;
 assign wire11553 = ( n_n4634 ) | ( n_n4639 ) | ( n_n4642 ) | ( n_n4631 ) ;
 assign wire11554 = ( n_n4629 ) | ( n_n4630 ) | ( wire190 ) ;
 assign wire11555 = ( n_n4637 ) | ( n_n4648 ) | ( n_n4628 ) | ( n_n4635 ) ;
 assign wire11558 = ( wire309 ) | ( n_n3861 ) | ( n_n4626 ) | ( wire11555 ) ;
 assign wire11559 = ( wire11548 ) | ( wire11549 ) | ( wire11553 ) | ( wire11554 ) ;
 assign wire11560 = ( n_n524  &  wire10  &  n_n509 ) | ( wire10  &  n_n534  &  n_n509 ) ;
 assign wire11562 = ( wire45 ) | ( wire256 ) ;
 assign wire11563 = ( wire396 ) | ( n_n4596 ) | ( wire11560 ) ;
 assign wire11566 = ( n_n524  &  wire10  &  n_n535 ) | ( wire10  &  n_n535  &  n_n520 ) ;
 assign wire11567 = ( wire25  &  n_n390  &  n_n535 ) | ( wire15  &  n_n390  &  n_n535 ) ;
 assign wire11568 = ( wire21  &  n_n390  &  n_n535 ) | ( n_n390  &  n_n535  &  wire23 ) ;
 assign wire11570 = ( n_n4593 ) | ( n_n4594 ) | ( wire365 ) ;
 assign wire11571 = ( wire11566 ) | ( wire11567 ) ;
 assign wire11574 = ( n_n4591 ) | ( n_n4592 ) | ( wire224 ) | ( wire11568 ) ;
 assign wire11575 = ( wire11562 ) | ( wire11563 ) | ( wire11570 ) | ( wire11571 ) ;
 assign wire11578 = ( n_n4537 ) | ( n_n4534 ) | ( wire11543 ) | ( wire11532 ) ;
 assign wire11581 = ( n_n1103 ) | ( wire11578 ) | ( _23016 ) | ( _23017 ) ;
 assign wire11582 = ( wire11558 ) | ( wire11559 ) | ( wire11574 ) | ( wire11575 ) ;
 assign wire11583 = ( wire16  &  n_n532  &  n_n535 ) | ( wire16  &  n_n534  &  n_n535 ) ;
 assign wire11584 = ( n_n526  &  wire16  &  n_n535 ) | ( wire16  &  n_n528  &  n_n535 ) ;
 assign wire11585 = ( wire22  &  n_n536  &  n_n535 ) | ( n_n536  &  wire24  &  n_n535 ) ;
 assign wire11586 = ( wire364 ) | ( wire11584 ) ;
 assign wire11587 = ( n_n4313 ) | ( wire11583 ) | ( wire11585 ) ;
 assign wire11588 = ( wire15  &  n_n491  &  n_n536 ) | ( n_n491  &  n_n536  &  wire20 ) ;
 assign wire11589 = ( n_n522  &  n_n491  &  wire16 ) | ( n_n491  &  n_n524  &  wire16 ) ;
 assign wire11591 = ( wire420 ) | ( wire11588 ) ;
 assign wire11592 = ( n_n4379 ) | ( n_n4380 ) | ( n_n4387 ) | ( wire11589 ) ;
 assign wire11593 = ( n_n482  &  wire21  &  n_n536 ) | ( n_n482  &  n_n536  &  wire23 ) ;
 assign wire11597 = ( n_n4404 ) | ( n_n4415 ) | ( wire11593 ) ;
 assign wire11598 = ( n_n4408 ) | ( n_n4406 ) | ( n_n4411 ) | ( wire328 ) ;
 assign wire11599 = ( n_n482  &  n_n526  &  wire16 ) | ( n_n482  &  wire16  &  n_n534 ) ;
 assign wire11613 = ( _1490 ) | ( wire16  &  n_n534  &  n_n500 ) ;
 assign wire11620 = ( i_9_  &  n_n524  &  n_n518  &  n_n536 ) | ( (~ i_9_)  &  n_n524  &  n_n518  &  n_n536 ) ;
 assign wire11625 = ( n_n4337 ) | ( n_n4344 ) | ( n_n4345 ) | ( n_n4343 ) ;
 assign wire11626 = ( n_n4342 ) | ( wire11620 ) | ( _23446 ) ;
 assign wire11628 = ( wire16  &  n_n518  &  n_n534 ) | ( wire16  &  n_n518  &  n_n528 ) ;
 assign wire11630 = ( n_n4331 ) | ( n_n4327 ) | ( n_n4330 ) | ( n_n4329 ) ;
 assign wire11631 = ( wire198 ) | ( n_n4322 ) | ( wire11628 ) ;
 assign wire11633 = ( wire11586 ) | ( wire11587 ) | ( wire11625 ) | ( wire11626 ) ;
 assign wire11634 = ( wire11630 ) | ( wire11631 ) | ( wire11633 ) ;
 assign wire11638 = ( n_n522  &  n_n491  &  wire10 ) | ( n_n491  &  wire10  &  n_n528 ) ;
 assign wire11653 = ( n_n4601 ) | ( n_n4571 ) | ( n_n4587 ) | ( n_n4584 ) ;
 assign wire11654 = ( n_n4574 ) | ( n_n4550 ) | ( n_n4527 ) | ( wire99 ) ;
 assign wire11658 = ( wire22  &  n_n464  &  n_n536 ) | ( n_n464  &  n_n536  &  wire23 ) ;
 assign wire11660 = ( n_n4455 ) | ( n_n4420 ) | ( n_n4430 ) | ( n_n4429 ) ;
 assign wire11661 = ( n_n4409 ) | ( n_n4410 ) | ( n_n4394 ) | ( wire11658 ) ;
 assign wire11671 = ( n_n473  &  wire15  &  n_n325 ) | ( wire15  &  n_n482  &  n_n325 ) ;
 assign wire11677 = ( i_9_  &  n_n528  &  n_n535  &  n_n260 ) | ( (~ i_9_)  &  n_n528  &  n_n535  &  n_n260 ) ;
 assign wire11687 = ( n_n4998 ) | ( n_n4887 ) | ( n_n4915 ) ;
 assign wire11688 = ( n_n4907 ) | ( n_n4879 ) | ( n_n4936 ) | ( n_n4947 ) ;
 assign wire11693 = ( wire19  &  n_n526  &  n_n518 ) | ( wire19  &  n_n526  &  n_n535 ) ;
 assign wire11694 = ( wire19  &  n_n528  &  n_n535 ) | ( wire19  &  n_n535  &  n_n520 ) ;
 assign wire11698 = ( n_n5254 ) | ( n_n5218 ) | ( wire11694 ) ;
 assign wire11699 = ( n_n5248 ) | ( n_n5213 ) | ( n_n5227 ) | ( wire11693 ) ;
 assign wire11703 = ( wire15  &  n_n464  &  n_n130 ) | ( n_n464  &  wire11  &  n_n130 ) ;
 assign wire11705 = ( n_n5206 ) | ( n_n5186 ) | ( n_n5182 ) | ( n_n5172 ) ;
 assign wire11706 = ( n_n5191 ) | ( n_n5209 ) | ( n_n5192 ) | ( wire11703 ) ;
 assign wire11707 = ( n_n532  &  wire12  &  n_n500 ) | ( n_n520  &  wire12  &  n_n500 ) ;
 assign wire11710 = ( i_9_  &  n_n509  &  n_n528  &  n_n130 ) | ( (~ i_9_)  &  n_n509  &  n_n528  &  n_n130 ) ;
 assign wire11712 = ( n_n5113 ) | ( n_n5155 ) | ( n_n5161 ) | ( n_n5127 ) ;
 assign wire11713 = ( n_n5108 ) | ( wire11707 ) | ( wire11710 ) ;
 assign wire11715 = ( wire15  &  n_n535  &  n_n130 ) | ( wire11  &  n_n535  &  n_n130 ) ;
 assign wire11731 = ( n_n5318 ) | ( n_n5320 ) | ( n_n5307 ) | ( n_n5329 ) ;
 assign wire11732 = ( n_n5302 ) | ( n_n5335 ) | ( n_n5304 ) | ( n_n5289 ) ;
 assign wire11738 = ( n_n522  &  wire16  &  n_n518 ) | ( n_n522  &  wire16  &  n_n535 ) ;
 assign wire11739 = ( n_n526  &  n_n491  &  wire16 ) | ( n_n491  &  wire16  &  n_n520 ) ;
 assign wire11743 = ( n_n1002 ) | ( wire11738 ) | ( wire11739 ) | ( _23316 ) ;
 assign wire11748 = ( n_n522  &  n_n491  &  wire14 ) | ( n_n491  &  wire14  &  n_n520 ) ;
 assign wire11751 = ( n_n4770 ) | ( n_n4769 ) | ( n_n4765 ) | ( n_n4766 ) ;
 assign wire11752 = ( n_n4767 ) | ( n_n4764 ) | ( n_n4771 ) | ( wire11748 ) ;
 assign wire11753 = ( n_n473  &  n_n526  &  wire14 ) | ( n_n473  &  wire14  &  n_n528 ) ;
 assign wire11754 = ( n_n473  &  n_n524  &  wire14 ) | ( n_n473  &  wire14  &  n_n520 ) ;
 assign wire11756 = ( n_n4810 ) | ( wire773 ) | ( wire11753 ) ;
 assign wire11757 = ( n_n4803 ) | ( n_n4804 ) | ( n_n4807 ) | ( wire11754 ) ;
 assign wire11759 = ( n_n524  &  n_n464  &  wire14 ) | ( n_n464  &  wire14  &  n_n520 ) ;
 assign wire11761 = ( _22359 ) | ( _22360 ) ;
 assign wire11762 = ( wire186 ) | ( wire85 ) | ( wire11759 ) ;
 assign wire11765 = ( n_n4787 ) | ( n_n4792 ) | ( n_n4793 ) | ( wire179 ) ;
 assign wire11766 = ( wire313 ) | ( wire292 ) | ( wire11765 ) ;
 assign wire11767 = ( wire11756 ) | ( wire11757 ) | ( wire11761 ) | ( wire11762 ) ;
 assign wire11768 = ( wire22  &  n_n518  &  n_n260 ) | ( n_n518  &  wire21  &  n_n260 ) ;
 assign wire11772 = ( n_n4862 ) | ( wire245 ) | ( n_n4861 ) ;
 assign wire11773 = ( n_n4856 ) | ( wire102 ) | ( n_n4853 ) | ( n_n4860 ) ;
 assign wire11774 = ( n_n518  &  wire24  &  n_n260 ) | ( wire24  &  n_n535  &  n_n260 ) ;
 assign wire11776 = ( n_n4825 ) | ( n_n4848 ) | ( n_n4826 ) ;
 assign wire11777 = ( n_n4842 ) | ( n_n4841 ) | ( wire11774 ) ;
 assign wire11778 = ( n_n4845 ) | ( n_n4846 ) | ( n_n4852 ) | ( wire11768 ) ;
 assign wire11781 = ( n_n3820 ) | ( n_n4836 ) | ( wire11769 ) | ( wire11778 ) ;
 assign wire11782 = ( wire11772 ) | ( wire11773 ) | ( wire11776 ) | ( wire11777 ) ;
 assign wire11783 = ( n_n482  &  n_n522  &  wire17 ) | ( n_n482  &  wire17  &  n_n530 ) ;
 assign wire11785 = ( n_n4913 ) | ( wire352 ) | ( n_n4914 ) ;
 assign wire11786 = ( n_n4911 ) | ( n_n4912 ) | ( n_n4905 ) | ( wire11783 ) ;
 assign wire11788 = ( n_n473  &  n_n524  &  wire17 ) | ( n_n473  &  n_n532  &  wire17 ) ;
 assign wire11790 = ( n_n4924 ) | ( n_n4921 ) | ( n_n4926 ) | ( n_n4925 ) ;
 assign wire11791 = ( n_n4920 ) | ( n_n4918 ) | ( n_n4919 ) | ( wire11788 ) ;
 assign wire11795 = ( n_n4937 ) | ( n_n4938 ) | ( n_n4931 ) | ( wire180 ) ;
 assign wire11797 = ( wire11785 ) | ( wire11786 ) | ( wire11790 ) | ( wire11791 ) ;
 assign wire11801 = ( n_n4963 ) | ( n_n4966 ) | ( wire771 ) | ( wire772 ) ;
 assign wire11802 = ( wire250 ) | ( n_n4968 ) | ( n_n4962 ) | ( n_n4971 ) ;
 assign wire11803 = ( n_n464  &  n_n528  &  wire17 ) | ( n_n464  &  wire17  &  n_n520 ) ;
 assign wire11804 = ( wire22  &  n_n464  &  n_n260 ) | ( n_n464  &  wire11  &  n_n260 ) ;
 assign wire11805 = ( n_n522  &  n_n464  &  wire17 ) | ( n_n524  &  n_n464  &  wire17 ) ;
 assign wire11807 = ( wire11803 ) | ( wire11804 ) ;
 assign wire11808 = ( n_n4955 ) | ( wire141 ) | ( wire11805 ) ;
 assign wire11809 = ( n_n518  &  n_n528  &  wire18 ) | ( n_n518  &  wire18  &  n_n530 ) ;
 assign wire11810 = ( wire22  &  n_n518  &  n_n195 ) | ( n_n518  &  wire11  &  n_n195 ) ;
 assign wire11811 = ( n_n518  &  wire21  &  n_n195 ) | ( n_n518  &  n_n195  &  wire20 ) ;
 assign wire11812 = ( n_n522  &  n_n518  &  wire18 ) | ( n_n524  &  n_n518  &  wire18 ) ;
 assign wire11814 = ( n_n4973 ) | ( wire11809 ) | ( wire11812 ) ;
 assign wire11816 = ( wire11801 ) | ( wire11802 ) | ( wire11807 ) | ( wire11808 ) ;
 assign wire11824 = ( wire40 ) | ( n_n4864 ) | ( n_n4867 ) | ( n_n4873 ) ;
 assign wire11825 = ( n_n491  &  n_n524  &  wire17 ) | ( n_n491  &  wire17  &  n_n520 ) ;
 assign wire11826 = ( n_n491  &  n_n260  &  wire20 ) | ( n_n491  &  n_n260  &  wire23 ) ;
 assign wire11829 = ( n_n4900 ) | ( n_n4899 ) | ( n_n4897 ) | ( wire11826 ) ;
 assign wire11834 = ( i_9_  &  n_n522  &  n_n325  &  n_n500 ) | ( (~ i_9_)  &  n_n522  &  n_n325  &  n_n500 ) ;
 assign wire11836 = ( n_n4760 ) | ( n_n4758 ) | ( n_n4761 ) | ( n_n4762 ) ;
 assign wire11837 = ( n_n4763 ) | ( wire11834 ) | ( _22321 ) ;
 assign wire11839 = ( i_9_  &  n_n325  &  n_n528  &  n_n500 ) | ( (~ i_9_)  &  n_n325  &  n_n528  &  n_n500 ) ;
 assign wire11841 = ( n_n4754 ) | ( n_n4753 ) | ( wire47 ) ;
 assign wire11842 = ( n_n4748 ) | ( n_n4747 ) | ( n_n4745 ) | ( wire11839 ) ;
 assign wire11846 = ( n_n4732 ) | ( n_n4725 ) | ( n_n4726 ) | ( wire767 ) ;
 assign wire11847 = ( n_n4737 ) | ( n_n4738 ) | ( wire293 ) ;
 assign wire11848 = ( n_n4733 ) | ( n_n4728 ) | ( n_n4743 ) | ( n_n4730 ) ;
 assign wire11855 = ( n_n4675 ) | ( n_n4676 ) | ( wire417 ) ;
 assign wire11859 = ( n_n4673 ) | ( n_n4662 ) | ( wire157 ) ;
 assign wire11870 = ( wire22  &  n_n325  &  n_n535 ) | ( n_n325  &  n_n535  &  wire20 ) ;
 assign wire11877 = ( wire25  &  n_n482  &  n_n390 ) | ( n_n482  &  wire21  &  n_n390 ) ;
 assign wire11880 = ( wire81 ) | ( wire418 ) | ( wire11877 ) ;
 assign wire11881 = ( n_n4652 ) | ( wire140 ) | ( wire391 ) | ( wire431 ) ;
 assign wire11886 = ( n_n482  &  n_n524  &  wire14 ) | ( n_n482  &  wire14  &  n_n528 ) ;
 assign wire11888 = ( n_n4784 ) | ( n_n4783 ) | ( wire315 ) ;
 assign wire11889 = ( n_n4779 ) | ( n_n4780 ) | ( n_n4775 ) | ( wire11886 ) ;
 assign wire11891 = ( wire11751 ) | ( wire11752 ) | ( wire11836 ) | ( wire11837 ) ;
 assign wire11893 = ( wire11766 ) | ( wire11767 ) | ( wire11781 ) | ( wire11782 ) ;
 assign wire11899 = ( n_n5162 ) | ( n_n5154 ) | ( wire287 ) ;
 assign wire11900 = ( n_n5152 ) | ( wire406 ) | ( n_n5159 ) | ( n_n5160 ) ;
 assign wire11902 = ( n_n482  &  wire22  &  n_n130 ) | ( n_n482  &  wire24  &  n_n130 ) ;
 assign wire11906 = ( wire114 ) | ( wire44 ) | ( _22749 ) ;
 assign wire11907 = ( wire33 ) | ( wire107 ) | ( wire113 ) | ( wire254 ) ;
 assign wire11909 = ( wire11899 ) | ( wire11900 ) | ( wire11907 ) ;
 assign wire11916 = ( n_n526  &  n_n509  &  wire12 ) | ( n_n534  &  n_n509  &  wire12 ) ;
 assign wire11917 = ( wire15  &  n_n509  &  n_n130 ) | ( wire22  &  n_n509  &  n_n130 ) ;
 assign wire11924 = ( wire25  &  n_n65  &  n_n500 ) | ( n_n65  &  wire20  &  n_n500 ) ;
 assign wire11928 = ( n_n65  &  n_n491  &  wire21 ) | ( n_n65  &  n_n491  &  wire23 ) ;
 assign wire11939 = ( n_n5299 ) | ( n_n5290 ) | ( n_n5291 ) | ( wire63 ) ;
 assign wire11947 = ( i_9_  &  n_n65  &  n_n464  &  n_n528 ) | ( (~ i_9_)  &  n_n65  &  n_n464  &  n_n528 ) ;
 assign wire11951 = ( n_n5322 ) | ( n_n5333 ) | ( n_n5319 ) | ( wire11946 ) ;
 assign wire11952 = ( wire148 ) | ( wire115 ) | ( wire175 ) | ( wire11947 ) ;
 assign wire11955 = ( wire25  &  n_n65  &  n_n509 ) | ( n_n65  &  wire24  &  n_n509 ) ;
 assign wire11959 = ( n_n5230 ) | ( n_n5233 ) | ( n_n5236 ) | ( wire320 ) ;
 assign wire11964 = ( wire19  &  n_n522  &  n_n535 ) | ( wire19  &  n_n535  &  n_n530 ) ;
 assign wire11967 = ( wire181 ) | ( wire11964 ) ;
 assign wire11968 = ( n_n5226 ) | ( n_n5225 ) | ( n_n5215 ) | ( wire384 ) ;
 assign wire11970 = ( n_n5189 ) | ( n_n5190 ) | ( wire452 ) ;
 assign wire11971 = ( n_n5200 ) | ( n_n5188 ) | ( n_n5194 ) | ( wire453 ) ;
 assign wire11972 = ( n_n464  &  wire21  &  n_n130 ) | ( n_n464  &  n_n130  &  wire23 ) ;
 assign wire11973 = ( wire19  &  n_n532  &  n_n535 ) | ( wire19  &  n_n534  &  n_n535 ) ;
 assign wire11978 = ( wire11967 ) | ( wire11968 ) | ( wire11970 ) | ( wire11971 ) ;
 assign wire11981 = ( wire248 ) | ( wire299 ) ;
 assign wire11982 = ( wire103 ) | ( n_n4994 ) | ( n_n5003 ) | ( n_n5006 ) ;
 assign wire11986 = ( n_n5017 ) | ( n_n5010 ) | ( n_n5019 ) | ( n_n5020 ) ;
 assign wire11987 = ( wire135 ) | ( n_n5012 ) | ( n_n5009 ) | ( n_n5007 ) ;
 assign wire11992 = ( n_n5050 ) | ( n_n5055 ) | ( n_n5059 ) | ( n_n5045 ) ;
 assign wire11993 = ( n_n5046 ) | ( n_n5056 ) | ( n_n5057 ) | ( wire166 ) ;
 assign wire11994 = ( n_n491  &  n_n524  &  wire18 ) | ( n_n491  &  n_n528  &  wire18 ) ;
 assign wire11995 = ( n_n5027 ) | ( n_n5028 ) | ( wire296 ) ;
 assign wire11996 = ( wire50 ) | ( n_n5029 ) | ( wire11994 ) ;
 assign wire11997 = ( n_n482  &  n_n532  &  wire18 ) | ( n_n482  &  n_n528  &  wire18 ) ;
 assign wire11999 = ( n_n482  &  wire22  &  n_n195 ) | ( n_n482  &  wire21  &  n_n195 ) ;
 assign wire12007 = ( n_n518  &  wire21  &  n_n130 ) | ( n_n518  &  wire20  &  n_n130 ) ;
 assign wire12018 = ( n_n5060 ) | ( n_n5067 ) | ( n_n5064 ) | ( wire755 ) ;
 assign wire12023 = ( n_n4983 ) | ( n_n4985 ) | ( n_n4984 ) ;
 assign wire12024 = ( n_n4988 ) | ( n_n4987 ) | ( wire104 ) ;
 assign wire12027 = ( wire11981 ) | ( wire11982 ) | ( wire11986 ) | ( wire11987 ) ;
 assign wire12033 = ( n_n5149 ) | ( n_n5138 ) | ( wire125 ) | ( n_n5143 ) ;
 assign wire12058 = ( n_n526  &  wire13  &  n_n500 ) | ( wire13  &  n_n500  &  n_n530 ) ;
 assign wire12060 = ( n_n4546 ) | ( n_n4555 ) | ( n_n4562 ) | ( n_n4506 ) ;
 assign wire12061 = ( n_n4512 ) | ( n_n4526 ) | ( n_n4535 ) | ( wire12058 ) ;
 assign wire12080 = ( n_n4790 ) | ( n_n4835 ) | ( n_n4788 ) ;
 assign wire12081 = ( n_n4774 ) | ( n_n4845 ) | ( n_n4796 ) | ( n_n4822 ) ;
 assign wire12089 = ( n_n4920 ) | ( n_n4907 ) | ( n_n4950 ) | ( n_n4894 ) ;
 assign wire12090 = ( n_n4916 ) | ( n_n4930 ) | ( n_n4947 ) | ( wire96 ) ;
 assign wire12091 = ( wire25  &  n_n130  &  n_n500 ) | ( wire24  &  n_n130  &  n_n500 ) ;
 assign wire12092 = ( i_9_  &  n_n526  &  n_n130  &  n_n500 ) | ( (~ i_9_)  &  n_n526  &  n_n130  &  n_n500 ) ;
 assign wire12093 = ( n_n526  &  n_n464  &  wire12 ) | ( n_n464  &  n_n520  &  wire12 ) ;
 assign wire12096 = ( wire12092 ) | ( wire12093 ) ;
 assign wire12097 = ( n_n5146 ) | ( n_n5204 ) | ( n_n5191 ) | ( wire12091 ) ;
 assign wire12099 = ( wire25  &  n_n535  &  n_n130 ) | ( wire22  &  n_n535  &  n_n130 ) ;
 assign wire12101 = ( n_n5096 ) | ( n_n5113 ) | ( n_n5066 ) | ( n_n5063 ) ;
 assign wire12102 = ( n_n5124 ) | ( wire335 ) | ( wire12099 ) ;
 assign wire12106 = ( wire19  &  n_n526  &  n_n535 ) | ( wire19  &  n_n535  &  n_n520 ) ;
 assign wire12108 = ( n_n5274 ) | ( n_n5232 ) | ( n_n5255 ) | ( n_n5267 ) ;
 assign wire12109 = ( n_n5244 ) | ( n_n5258 ) | ( n_n5212 ) | ( wire12106 ) ;
 assign wire12111 = ( wire12096 ) | ( wire12097 ) | ( wire12101 ) | ( wire12102 ) ;
 assign wire12113 = ( n_n522  &  n_n491  &  wire18 ) | ( n_n491  &  n_n528  &  wire18 ) ;
 assign wire12114 = ( n_n482  &  wire21  &  n_n195 ) | ( n_n482  &  n_n195  &  wire20 ) ;
 assign wire12115 = ( n_n473  &  wire15  &  n_n195 ) | ( n_n473  &  wire22  &  n_n195 ) ;
 assign wire12117 = ( wire12113 ) | ( wire12114 ) ;
 assign wire12118 = ( n_n5025 ) | ( n_n5048 ) | ( n_n5009 ) | ( wire12115 ) ;
 assign wire12120 = ( n_n522  &  n_n518  &  wire18 ) | ( n_n518  &  n_n528  &  wire18 ) ;
 assign wire12126 = ( n_n482  &  wire19  &  n_n528 ) | ( n_n482  &  wire19  &  n_n520 ) ;
 assign wire12128 = ( n_n5321 ) | ( n_n5326 ) | ( n_n5335 ) | ( wire12126 ) ;
 assign wire12129 = ( wire12089 ) | ( wire12090 ) | ( wire12128 ) ;
 assign wire12131 = ( n_n1333 ) | ( wire12117 ) | ( wire12118 ) | ( wire12129 ) ;
 assign wire12134 = ( wire25  &  n_n473  &  n_n536 ) | ( n_n473  &  wire22  &  n_n536 ) ;
 assign wire12136 = ( n_n4407 ) | ( n_n4430 ) | ( _23965 ) ;
 assign wire12137 = ( wire84 ) | ( n_n4410 ) | ( wire12134 ) ;
 assign wire12141 = ( n_n4340 ) | ( n_n4345 ) | ( wire399 ) ;
 assign wire12142 = ( n_n4331 ) | ( n_n4312 ) | ( n_n4326 ) | ( wire156 ) ;
 assign wire12146 = ( n_n4400 ) | ( n_n4383 ) | ( n_n4369 ) | ( n_n4372 ) ;
 assign wire12147 = ( n_n4397 ) | ( n_n4360 ) | ( wire423 ) | ( n_n4375 ) ;
 assign wire12149 = ( wire12136 ) | ( wire12137 ) | ( wire12141 ) | ( wire12142 ) ;
 assign wire12152 = ( wire12131 ) | ( wire12149 ) | ( _23986 ) | ( _23987 ) ;
 assign wire12162 = ( wire15  &  n_n535  &  n_n195 ) | ( wire22  &  n_n535  &  n_n195 ) ;
 assign wire12164 = ( n_n4951 ) | ( n_n4952 ) | ( n_n4959 ) | ( n_n4960 ) ;
 assign wire12165 = ( wire250 ) | ( n_n4953 ) | ( wire12162 ) ;
 assign wire12167 = ( n_n464  &  wire24  &  n_n260 ) | ( n_n464  &  n_n260  &  wire20 ) ;
 assign wire12168 = ( n_n4937 ) | ( n_n4938 ) | ( n_n4944 ) ;
 assign wire12169 = ( wire59 ) | ( wire12166 ) | ( wire12167 ) ;
 assign wire12170 = ( n_n473  &  n_n528  &  wire17 ) | ( n_n473  &  wire17  &  n_n520 ) ;
 assign wire12171 = ( n_n524  &  n_n464  &  wire17 ) | ( n_n464  &  n_n534  &  wire17 ) ;
 assign wire12172 = ( n_n473  &  wire21  &  n_n260 ) | ( n_n473  &  n_n260  &  wire20 ) ;
 assign wire12175 = ( wire31 ) | ( wire42 ) | ( wire12172 ) ;
 assign wire12176 = ( wire12170 ) | ( wire12171 ) | ( wire12175 ) ;
 assign wire12177 = ( wire12164 ) | ( wire12165 ) | ( wire12168 ) | ( wire12169 ) ;
 assign wire12181 = ( wire260 ) | ( wire49 ) ;
 assign wire12182 = ( n_n4888 ) | ( n_n4895 ) | ( n_n4889 ) | ( wire12179 ) ;
 assign wire12183 = ( wire25  &  n_n482  &  n_n260 ) | ( n_n482  &  wire22  &  n_n260 ) ;
 assign wire12186 = ( n_n4911 ) | ( n_n4912 ) | ( n_n4901 ) | ( n_n4904 ) ;
 assign wire12187 = ( wire305 ) | ( wire12183 ) ;
 assign wire12188 = ( n_n4917 ) | ( n_n4914 ) | ( n_n4915 ) | ( n_n4910 ) ;
 assign wire12191 = ( n_n3810 ) | ( n_n1592 ) | ( wire12188 ) ;
 assign wire12192 = ( wire12181 ) | ( wire12182 ) | ( wire12186 ) | ( wire12187 ) ;
 assign wire12196 = ( n_n4964 ) | ( n_n4968 ) | ( wire342 ) | ( n_n4973 ) ;
 assign wire12202 = ( n_n482  &  wire21  &  n_n325 ) | ( n_n482  &  n_n325  &  wire20 ) ;
 assign wire12204 = ( n_n4784 ) | ( n_n4791 ) | ( wire158 ) ;
 assign wire12205 = ( wire179 ) | ( n_n4799 ) | ( wire12202 ) ;
 assign wire12210 = ( n_n534  &  n_n509  &  wire17 ) | ( n_n509  &  wire17  &  n_n530 ) ;
 assign wire12213 = ( wire277 ) | ( wire12210 ) ;
 assign wire12214 = ( wire245 ) | ( n_n4864 ) | ( n_n4865 ) | ( n_n4854 ) ;
 assign wire12217 = ( wire21  &  n_n509  &  n_n260 ) | ( n_n509  &  n_n260  &  wire23 ) ;
 assign wire12218 = ( n_n4882 ) | ( n_n4881 ) | ( wire330 ) ;
 assign wire12219 = ( n_n4868 ) | ( n_n4880 ) | ( wire324 ) ;
 assign wire12220 = ( n_n4877 ) | ( n_n4870 ) | ( wire12217 ) ;
 assign wire12226 = ( i_9_  &  n_n528  &  n_n535  &  n_n260 ) | ( (~ i_9_)  &  n_n528  &  n_n535  &  n_n260 ) ;
 assign wire12232 = ( wire22  &  n_n518  &  n_n260 ) | ( n_n518  &  wire24  &  n_n260 ) ;
 assign wire12239 = ( n_n4817 ) | ( n_n4824 ) | ( wire85 ) | ( wire12225 ) ;
 assign wire12243 = ( n_n4803 ) | ( n_n4804 ) | ( n_n4807 ) | ( n_n4808 ) ;
 assign wire12245 = ( n_n4802 ) | ( n_n4805 ) | ( n_n4197 ) | ( wire12243 ) ;
 assign wire12253 = ( n_n5026 ) | ( n_n5017 ) | ( wire135 ) | ( n_n5016 ) ;
 assign wire12262 = ( n_n5157 ) | ( n_n5152 ) | ( n_n5149 ) | ( wire195 ) ;
 assign wire12266 = ( n_n5135 ) | ( n_n5148 ) | ( wire125 ) | ( n_n5144 ) ;
 assign wire12268 = ( wire22  &  n_n464  &  n_n130 ) | ( n_n464  &  wire11  &  n_n130 ) ;
 assign wire12269 = ( wire15  &  n_n464  &  n_n130 ) | ( n_n464  &  wire21  &  n_n130 ) ;
 assign wire12271 = ( wire453 ) | ( wire12268 ) ;
 assign wire12272 = ( wire452 ) | ( n_n5192 ) | ( wire12269 ) ;
 assign wire12276 = ( _1230 ) | ( wire19  &  n_n524  &  n_n518 ) ;
 assign wire12277 = ( n_n5207 ) | ( n_n5208 ) | ( n_n5205 ) ;
 assign wire12278 = ( n_n5230 ) | ( n_n5223 ) | ( n_n5233 ) | ( n_n5220 ) ;
 assign wire12282 = ( n_n1530 ) | ( n_n1532 ) | ( n_n763 ) | ( wire12276 ) ;
 assign wire12283 = ( wire12271 ) | ( wire12272 ) | ( wire12277 ) | ( wire12278 ) ;
 assign wire12285 = ( i_9_  &  n_n482  &  n_n528  &  n_n130 ) | ( (~ i_9_)  &  n_n482  &  n_n528  &  n_n130 ) ;
 assign wire12288 = ( n_n5163 ) | ( wire33 ) | ( wire12285 ) ;
 assign wire12290 = ( wire25  &  n_n473  &  n_n130 ) | ( n_n473  &  wire21  &  n_n130 ) ;
 assign wire12292 = ( n_n5189 ) | ( n_n5190 ) | ( wire332 ) ;
 assign wire12293 = ( n_n5171 ) | ( n_n5186 ) | ( wire12290 ) ;
 assign wire12296 = ( n_n4129 ) | ( wire44 ) | ( n_n5176 ) | ( wire12293 ) ;
 assign wire12297 = ( wire12288 ) | ( wire12292 ) | ( _24373 ) ;
 assign wire12300 = ( n_n5128 ) | ( n_n5121 ) | ( n_n5122 ) ;
 assign wire12301 = ( n_n5130 ) | ( n_n5120 ) | ( wire286 ) ;
 assign wire12304 = ( wire12262 ) | ( wire12266 ) | ( _24317 ) ;
 assign wire12306 = ( wire12282 ) | ( wire12283 ) | ( wire12296 ) | ( wire12297 ) ;
 assign wire12317 = ( wire15  &  n_n464  &  n_n195 ) | ( wire22  &  n_n464  &  n_n195 ) ;
 assign wire12318 = ( n_n526  &  n_n464  &  wire18 ) | ( n_n524  &  n_n464  &  wire18 ) ;
 assign wire12319 = ( n_n522  &  n_n464  &  wire18 ) | ( n_n464  &  n_n528  &  wire18 ) ;
 assign wire12323 = ( n_n5075 ) | ( n_n5068 ) | ( n_n5071 ) | ( wire12317 ) ;
 assign wire12326 = ( wire15  &  n_n509  &  n_n130 ) | ( wire24  &  n_n509  &  n_n130 ) ;
 assign wire12335 = ( wire21  &  n_n535  &  n_n130 ) | ( n_n535  &  wire20  &  n_n130 ) ;
 assign wire12337 = ( n_n5098 ) | ( n_n5095 ) | ( wire88 ) ;
 assign wire12342 = ( n_n65  &  wire15  &  n_n482 ) | ( n_n65  &  n_n482  &  wire11 ) ;
 assign wire12345 = ( n_n5289 ) | ( wire12342 ) | ( _24448 ) ;
 assign wire12355 = ( wire19  &  n_n528  &  n_n500 ) | ( wire19  &  n_n500  &  n_n530 ) ;
 assign wire12356 = ( i_9_  &  n_n65  &  n_n526  &  n_n500 ) | ( (~ i_9_)  &  n_n65  &  n_n526  &  n_n500 ) ;
 assign wire12358 = ( n_n5272 ) | ( n_n5271 ) | ( n_n5270 ) | ( wire12356 ) ;
 assign wire12359 = ( wire77 ) | ( wire12355 ) | ( wire12358 ) ;
 assign wire12361 = ( n_n65  &  n_n464  &  wire11 ) | ( n_n65  &  n_n464  &  wire24 ) ;
 assign wire12366 = ( n_n473  &  n_n65  &  wire15 ) | ( n_n473  &  n_n65  &  wire11 ) ;
 assign wire12376 = ( n_n5303 ) | ( n_n5304 ) | ( wire63 ) ;
 assign wire12380 = ( wire12345 ) | ( wire12376 ) | ( _24456 ) ;
 assign wire12382 = ( n_n1435 ) | ( n_n1436 ) | ( wire12359 ) | ( wire12380 ) ;
 assign wire12384 = ( n_n491  &  n_n195  &  wire20 ) | ( n_n491  &  n_n195  &  wire23 ) ;
 assign wire12386 = ( n_n5038 ) | ( n_n5035 ) | ( n_n5037 ) | ( wire12384 ) ;
 assign wire12389 = ( n_n1454 ) | ( wire12386 ) | ( _24285 ) | ( _24286 ) ;
 assign wire12391 = ( n_n1409 ) | ( n_n1408 ) | ( wire12389 ) ;
 assign wire12392 = ( wire12306 ) | ( wire12382 ) | ( _24460 ) ;
 assign wire12395 = ( n_n4765 ) | ( n_n4766 ) | ( n_n4762 ) ;
 assign wire12398 = ( i_9_  &  n_n522  &  n_n509  &  n_n325 ) | ( (~ i_9_)  &  n_n522  &  n_n509  &  n_n325 ) ;
 assign wire12399 = ( n_n4738 ) | ( n_n4744 ) | ( n_n4739 ) | ( n_n4745 ) ;
 assign wire12400 = ( wire95 ) | ( n_n4736 ) | ( wire12398 ) ;
 assign wire12401 = ( wire25  &  n_n325  &  n_n535 ) | ( wire11  &  n_n325  &  n_n535 ) ;
 assign wire12413 = ( n_n4718 ) | ( n_n4717 ) | ( n_n4713 ) ;
 assign wire12414 = ( n_n4704 ) | ( n_n4711 ) | ( n_n4710 ) | ( n_n4709 ) ;
 assign wire12420 = ( n_n4673 ) | ( n_n4670 ) | ( wire417 ) ;
 assign wire12421 = ( n_n4674 ) | ( n_n4671 ) | ( wire81 ) | ( wire418 ) ;
 assign wire12422 = ( n_n522  &  n_n464  &  wire10 ) | ( n_n464  &  wire10  &  n_n520 ) ;
 assign wire12425 = ( wire157 ) | ( wire225 ) ;
 assign wire12426 = ( n_n4667 ) | ( n_n4662 ) | ( n_n4660 ) | ( wire72 ) ;
 assign wire12428 = ( wire15  &  n_n464  &  n_n390 ) | ( n_n464  &  wire11  &  n_n390 ) ;
 assign wire12435 = ( n_n4748 ) | ( n_n4747 ) | ( n_n4761 ) ;
 assign wire12436 = ( n_n4754 ) | ( n_n4757 ) | ( n_n4749 ) | ( n_n4760 ) ;
 assign wire12439 = ( wire447 ) | ( wire12395 ) | ( wire12399 ) | ( wire12400 ) ;
 assign wire12442 = ( wire21  &  n_n536  &  n_n500 ) | ( n_n536  &  wire20  &  n_n500 ) ;
 assign wire12445 = ( n_n4367 ) | ( n_n4368 ) | ( wire12442 ) ;
 assign wire12446 = ( n_n4374 ) | ( wire280 ) | ( n_n4365 ) | ( n_n4370 ) ;
 assign wire12448 = ( n_n522  &  n_n491  &  wire16 ) | ( n_n491  &  wire16  &  n_n520 ) ;
 assign wire12451 = ( _23507 ) | ( _23508 ) ;
 assign wire12453 = ( n_n4386 ) | ( wire12447 ) | ( n_n4387 ) | ( wire12448 ) ;
 assign wire12456 = ( wire27 ) | ( wire12445 ) | ( wire12446 ) | ( wire12451 ) ;
 assign wire12461 = ( n_n482  &  wire16  &  n_n534 ) | ( n_n482  &  wire16  &  n_n528 ) ;
 assign wire12467 = ( wire98 ) | ( n_n4421 ) | ( wire215 ) | ( n_n4429 ) ;
 assign wire12472 = ( wire13  &  n_n534  &  n_n535 ) | ( wire13  &  n_n535  &  n_n530 ) ;
 assign wire12475 = ( n_n4445 ) | ( n_n4446 ) | ( wire12472 ) ;
 assign wire12476 = ( n_n4437 ) | ( n_n4447 ) | ( n_n4435 ) | ( wire421 ) ;
 assign wire12478 = ( i_9_  &  n_n522  &  n_n455  &  n_n535 ) | ( (~ i_9_)  &  n_n522  &  n_n455  &  n_n535 ) ;
 assign wire12479 = ( _1428 ) | ( wire21  &  n_n455  &  n_n535 ) ;
 assign wire12480 = ( n_n4464 ) | ( n_n4463 ) | ( n_n4465 ) ;
 assign wire12481 = ( wire128 ) | ( wire12478 ) ;
 assign wire12485 = ( n_n3162 ) | ( wire55 ) | ( n_n2058 ) | ( wire12479 ) ;
 assign wire12486 = ( wire12475 ) | ( wire12476 ) | ( wire12480 ) | ( wire12481 ) ;
 assign wire12488 = ( wire15  &  n_n455  &  n_n500 ) | ( wire22  &  n_n455  &  n_n500 ) ;
 assign wire12490 = ( n_n4488 ) | ( n_n4487 ) | ( n_n4486 ) | ( wire12488 ) ;
 assign wire12497 = ( wire416 ) | ( wire201 ) ;
 assign wire12498 = ( n_n4547 ) | ( n_n4538 ) | ( wire212 ) | ( n_n4545 ) ;
 assign wire12499 = ( wire25  &  n_n482  &  n_n455 ) | ( n_n482  &  wire21  &  n_n455 ) ;
 assign wire12500 = ( i_9_  &  n_n473  &  n_n455  &  n_n534 ) | ( (~ i_9_)  &  n_n473  &  n_n455  &  n_n534 ) ;
 assign wire12501 = ( n_n482  &  n_n526  &  wire13 ) | ( n_n482  &  wire13  &  n_n520 ) ;
 assign wire12502 = ( wire170 ) | ( n_n4529 ) | ( wire724 ) ;
 assign wire12503 = ( wire361 ) | ( wire12499 ) ;
 assign wire12507 = ( n_n4247 ) | ( n_n3879 ) | ( wire12500 ) | ( wire12501 ) ;
 assign wire12508 = ( wire12497 ) | ( wire12498 ) | ( wire12502 ) | ( wire12503 ) ;
 assign wire12510 = ( wire15  &  n_n491  &  n_n455 ) | ( n_n491  &  n_n455  &  wire24 ) ;
 assign wire12514 = ( wire308 ) | ( n_n4505 ) | ( n_n4501 ) | ( n_n4499 ) ;
 assign wire12518 = ( wire12485 ) | ( wire12486 ) | ( wire12507 ) | ( wire12508 ) ;
 assign wire12519 = ( i_9_  &  n_n390  &  n_n509  &  n_n528 ) | ( (~ i_9_)  &  n_n390  &  n_n509  &  n_n528 ) ;
 assign wire12520 = ( i_9_  &  n_n518  &  n_n532  &  n_n390 ) | ( (~ i_9_)  &  n_n518  &  n_n532  &  n_n390 ) ;
 assign wire12521 = ( i_9_  &  n_n532  &  n_n390  &  n_n535 ) | ( (~ i_9_)  &  n_n532  &  n_n390  &  n_n535 ) ;
 assign wire12525 = ( n_n4561 ) | ( n_n4568 ) | ( n_n4572 ) | ( wire238 ) ;
 assign wire12530 = ( n_n4557 ) | ( n_n4560 ) | ( n_n4582 ) | ( n_n4581 ) ;
 assign wire12531 = ( n_n4554 ) | ( n_n4584 ) | ( n_n4577 ) | ( n_n4556 ) ;
 assign wire12534 = ( n_n3871 ) | ( n_n4585 ) | ( wire12520 ) | ( wire12531 ) ;
 assign wire12535 = ( wire12525 ) | ( wire12530 ) | ( _23708 ) ;
 assign wire12539 = ( n_n4616 ) | ( n_n4612 ) | ( n_n4611 ) | ( n_n4619 ) ;
 assign wire12540 = ( n_n4608 ) | ( wire465 ) | ( n_n4620 ) | ( n_n4609 ) ;
 assign wire12541 = ( n_n518  &  wire10  &  n_n528 ) | ( n_n518  &  wire10  &  n_n520 ) ;
 assign wire12543 = ( n_n4593 ) | ( n_n4594 ) | ( wire255 ) ;
 assign wire12544 = ( wire365 ) | ( n_n4595 ) | ( wire12541 ) ;
 assign wire12545 = ( n_n526  &  wire10  &  n_n500 ) | ( n_n524  &  wire10  &  n_n500 ) ;
 assign wire12546 = ( i_9_  &  n_n522  &  n_n390  &  n_n500 ) | ( (~ i_9_)  &  n_n522  &  n_n390  &  n_n500 ) ;
 assign wire12547 = ( wire25  &  n_n491  &  n_n390 ) | ( wire15  &  n_n491  &  n_n390 ) ;
 assign wire12551 = ( n_n4648 ) | ( n_n4646 ) | ( wire391 ) ;
 assign wire12552 = ( n_n4644 ) | ( wire311 ) | ( n_n4650 ) | ( n_n4654 ) ;
 assign wire12554 = ( n_n4630 ) | ( n_n4631 ) | ( n_n4632 ) ;
 assign wire12555 = ( wire310 ) | ( wire401 ) ;
 assign wire12556 = ( n_n4640 ) | ( n_n4621 ) | ( n_n4625 ) | ( wire12545 ) ;
 assign wire12557 = ( n_n4639 ) | ( n_n4627 ) | ( wire12546 ) | ( wire12547 ) ;
 assign wire12559 = ( wire12556 ) | ( wire12557 ) ;
 assign wire12560 = ( wire12551 ) | ( wire12552 ) | ( wire12554 ) | ( wire12555 ) ;
 assign wire12561 = ( i_9_  &  n_n390  &  n_n534  &  n_n509 ) | ( (~ i_9_)  &  n_n390  &  n_n534  &  n_n509 ) ;
 assign wire12564 = ( n_n4599 ) | ( wire12519 ) | ( _23648 ) ;
 assign wire12566 = ( wire12539 ) | ( wire12540 ) | ( wire12543 ) | ( wire12544 ) ;
 assign wire12568 = ( wire12534 ) | ( wire12535 ) | ( wire12559 ) | ( wire12560 ) ;
 assign wire12569 = ( n_n522  &  wire16  &  n_n535 ) | ( n_n524  &  wire16  &  n_n535 ) ;
 assign wire12570 = ( i_9_  &  n_n526  &  n_n518  &  n_n536 ) | ( (~ i_9_)  &  n_n526  &  n_n518  &  n_n536 ) ;
 assign wire12573 = ( n_n4335 ) | ( n_n4344 ) | ( n_n4341 ) | ( wire12570 ) ;
 assign wire12574 = ( n_n526  &  wire16  &  n_n535 ) | ( wire16  &  n_n528  &  n_n535 ) ;
 assign wire12577 = ( n_n4313 ) | ( wire171 ) | ( wire12574 ) ;
 assign wire12578 = ( wire16  &  n_n518  &  n_n534 ) | ( wire16  &  n_n518  &  n_n530 ) ;
 assign wire12579 = ( n_n4330 ) | ( n_n4329 ) | ( wire106 ) ;
 assign wire12582 = ( wire12573 ) | ( wire12577 ) | ( _23538 ) ;
 assign wire12602 = ( n_n473  &  n_n455  &  wire24 ) | ( n_n482  &  n_n455  &  wire24 ) ;
 assign wire12607 = ( n_n4557 ) | ( n_n4572 ) | ( n_n4531 ) | ( n_n4555 ) ;
 assign wire12608 = ( n_n4528 ) | ( n_n4549 ) | ( n_n4559 ) | ( wire12602 ) ;
 assign wire12613 = ( n_n4756 ) | ( n_n4753 ) | ( n_n4765 ) | ( n_n4766 ) ;
 assign wire12614 = ( wire131 ) | ( n_n4792 ) | ( n_n4764 ) | ( n_n4763 ) ;
 assign wire12615 = ( n_n473  &  wire10  &  n_n528 ) | ( n_n473  &  wire10  &  n_n530 ) ;
 assign wire12620 = ( n_n4656 ) | ( n_n4676 ) | ( n_n4703 ) | ( n_n4698 ) ;
 assign wire12621 = ( n_n4672 ) | ( n_n4692 ) | ( n_n4686 ) | ( wire12615 ) ;
 assign wire12626 = ( n_n4735 ) | ( n_n4749 ) | ( n_n4740 ) ;
 assign wire12627 = ( n_n4718 ) | ( n_n4727 ) | ( n_n4733 ) | ( n_n4730 ) ;
 assign wire12629 = ( n_n4750 ) | ( n_n4736 ) | ( wire12626 ) | ( wire12627 ) ;
 assign wire12630 = ( wire12613 ) | ( wire12614 ) | ( wire12620 ) | ( wire12621 ) ;
 assign wire12634 = ( n_n5258 ) | ( n_n5212 ) | ( n_n5262 ) | ( n_n5259 ) ;
 assign wire12635 = ( n_n5266 ) | ( n_n5236 ) | ( n_n5235 ) | ( wire320 ) ;
 assign wire12638 = ( n_n482  &  n_n526  &  wire12 ) | ( n_n482  &  n_n528  &  wire12 ) ;
 assign wire12640 = ( n_n5183 ) | ( n_n5204 ) | ( n_n5182 ) | ( n_n5173 ) ;
 assign wire12641 = ( wire114 ) | ( n_n5211 ) | ( wire12638 ) ;
 assign wire12642 = ( n_n491  &  wire21  &  n_n130 ) | ( wire21  &  n_n509  &  n_n130 ) ;
 assign wire12643 = ( wire15  &  n_n482  &  n_n130 ) | ( wire15  &  n_n509  &  n_n130 ) ;
 assign wire12648 = ( n_n5121 ) | ( n_n5134 ) | ( n_n5151 ) | ( wire12642 ) ;
 assign wire12649 = ( n_n5135 ) | ( n_n5158 ) | ( wire12643 ) | ( wire12648 ) ;
 assign wire12650 = ( wire12634 ) | ( wire12635 ) | ( wire12640 ) | ( wire12641 ) ;
 assign wire12651 = ( n_n518  &  n_n534  &  wire12 ) | ( n_n518  &  wire12  &  n_n530 ) ;
 assign wire12653 = ( wire22  &  n_n518  &  n_n130 ) | ( n_n518  &  wire11  &  n_n130 ) ;
 assign wire12656 = ( n_n5089 ) | ( n_n5098 ) | ( wire12653 ) ;
 assign wire12657 = ( n_n5104 ) | ( n_n5078 ) | ( n_n5090 ) | ( wire12651 ) ;
 assign wire12658 = ( n_n526  &  n_n518  &  wire18 ) | ( n_n526  &  n_n509  &  wire18 ) ;
 assign wire12659 = ( n_n491  &  wire24  &  n_n195 ) | ( wire24  &  n_n509  &  n_n195 ) ;
 assign wire12663 = ( n_n5010 ) | ( n_n4966 ) | ( wire12659 ) ;
 assign wire12664 = ( n_n5011 ) | ( n_n4961 ) | ( wire706 ) | ( wire12658 ) ;
 assign wire12669 = ( n_n5027 ) | ( n_n5048 ) | ( wire695 ) ;
 assign wire12670 = ( n_n5042 ) | ( n_n5022 ) | ( n_n5067 ) | ( n_n5020 ) ;
 assign wire12672 = ( n_n5072 ) | ( n_n5075 ) | ( wire12669 ) | ( wire12670 ) ;
 assign wire12673 = ( wire12656 ) | ( wire12657 ) | ( wire12663 ) | ( wire12664 ) ;
 assign wire12675 = ( n_n491  &  wire11  &  n_n260 ) | ( n_n491  &  n_n260  &  wire23 ) ;
 assign wire12678 = ( n_n4885 ) | ( n_n4911 ) | ( wire12675 ) ;
 assign wire12679 = ( n_n4886 ) | ( n_n4890 ) | ( n_n4892 ) | ( wire324 ) ;
 assign wire12688 = ( n_n4918 ) | ( n_n4917 ) | ( n_n4954 ) ;
 assign wire12689 = ( n_n4928 ) | ( n_n4950 ) | ( n_n4936 ) | ( n_n4956 ) ;
 assign wire12691 = ( n_n4931 ) | ( n_n4948 ) | ( wire12688 ) | ( wire12689 ) ;
 assign wire12693 = ( n_n554 ) | ( wire12678 ) | ( wire12679 ) | ( wire12691 ) ;
 assign wire12694 = ( wire12649 ) | ( wire12650 ) | ( wire12672 ) | ( wire12673 ) ;
 assign wire12710 = ( n_n536  &  wire24  &  n_n509 ) | ( n_n536  &  wire24  &  n_n500 ) ;
 assign wire12722 = ( wire15  &  n_n491  &  n_n260 ) | ( n_n491  &  wire22  &  n_n260 ) ;
 assign wire12724 = ( n_n4898 ) | ( n_n4901 ) | ( n_n4904 ) | ( n_n4899 ) ;
 assign wire12729 = ( n_n4869 ) | ( n_n4876 ) | ( wire330 ) ;
 assign wire12730 = ( wire295 ) | ( n_n4871 ) | ( n_n4875 ) | ( n_n4874 ) ;
 assign wire12732 = ( n_n526  &  n_n509  &  wire17 ) | ( n_n509  &  wire17  &  n_n530 ) ;
 assign wire12735 = ( n_n4857 ) | ( n_n4862 ) | ( wire12732 ) ;
 assign wire12736 = ( wire277 ) | ( n_n4861 ) | ( n_n4851 ) | ( n_n4863 ) ;
 assign wire12740 = ( wire22  &  n_n535  &  n_n260 ) | ( n_n535  &  n_n260  &  wire20 ) ;
 assign wire12742 = ( n_n4835 ) | ( n_n4832 ) | ( n_n4828 ) | ( n_n4839 ) ;
 assign wire12743 = ( n_n4838 ) | ( wire304 ) | ( wire12740 ) ;
 assign wire12744 = ( wire15  &  n_n518  &  n_n260 ) | ( n_n518  &  wire24  &  n_n260 ) ;
 assign wire12745 = ( n_n518  &  n_n534  &  wire17 ) | ( n_n518  &  wire17  &  n_n530 ) ;
 assign wire12747 = ( wire52 ) | ( wire150 ) ;
 assign wire12748 = ( n_n4827 ) | ( n_n4824 ) | ( wire12744 ) ;
 assign wire12749 = ( n_n4822 ) | ( n_n4826 ) | ( wire12745 ) ;
 assign wire12759 = ( wire25  &  n_n482  &  n_n325 ) | ( n_n482  &  wire24  &  n_n325 ) ;
 assign wire12760 = ( n_n482  &  n_n522  &  wire14 ) | ( n_n482  &  n_n532  &  wire14 ) ;
 assign wire12766 = ( n_n4789 ) | ( n_n4793 ) | ( n_n4797 ) | ( wire179 ) ;
 assign wire12770 = ( n_n4884 ) | ( n_n4883 ) | ( n_n4891 ) ;
 assign wire12771 = ( n_n4882 ) | ( n_n4881 ) | ( wire261 ) ;
 assign wire12774 = ( wire12729 ) | ( wire12730 ) | ( wire12735 ) | ( wire12736 ) ;
 assign wire12787 = ( wire15  &  n_n518  &  n_n325 ) | ( n_n518  &  wire11  &  n_n325 ) ;
 assign wire12788 = ( n_n518  &  wire21  &  n_n325 ) | ( n_n518  &  wire24  &  n_n325 ) ;
 assign wire12792 = ( wire25  &  n_n325  &  n_n535 ) | ( wire24  &  n_n325  &  n_n535 ) ;
 assign wire12794 = ( n_n4695 ) | ( n_n4696 ) | ( wire12792 ) ;
 assign wire12799 = ( n_n4683 ) | ( n_n4684 ) | ( wire417 ) ;
 assign wire12800 = ( n_n4677 ) | ( wire81 ) | ( wire418 ) | ( n_n4685 ) ;
 assign wire12801 = ( i_9_  &  n_n473  &  n_n532  &  n_n390 ) | ( (~ i_9_)  &  n_n473  &  n_n532  &  n_n390 ) ;
 assign wire12802 = ( n_n473  &  wire15  &  n_n390 ) | ( n_n473  &  wire21  &  n_n390 ) ;
 assign wire12804 = ( wire225 ) | ( wire12801 ) ;
 assign wire12805 = ( n_n4674 ) | ( n_n4673 ) | ( n_n4671 ) | ( wire12802 ) ;
 assign wire12810 = ( n_n4644 ) | ( n_n4649 ) | ( n_n4657 ) ;
 assign wire12811 = ( n_n4662 ) | ( n_n4659 ) | ( n_n4655 ) | ( n_n4658 ) ;
 assign wire12815 = ( wire21  &  n_n325  &  n_n500 ) | ( n_n325  &  wire20  &  n_n500 ) ;
 assign wire12819 = ( n_n4758 ) | ( n_n4747 ) | ( wire12815 ) ;
 assign wire12820 = ( n_n4752 ) | ( wire47 ) | ( n_n4751 ) | ( n_n4745 ) ;
 assign wire12822 = ( n_n4760 ) | ( n_n4769 ) | ( n_n4762 ) ;
 assign wire12826 = ( n_n856 ) | ( wire12819 ) | ( wire12820 ) | ( wire12822 ) ;
 assign wire12831 = ( wire15  &  n_n535  &  n_n195 ) | ( wire11  &  n_n535  &  n_n195 ) ;
 assign wire12832 = ( wire25  &  n_n535  &  n_n195 ) | ( wire24  &  n_n535  &  n_n195 ) ;
 assign wire12833 = ( n_n4952 ) | ( n_n4949 ) | ( wire12831 ) ;
 assign wire12834 = ( n_n4945 ) | ( n_n4946 ) | ( n_n4947 ) | ( wire12832 ) ;
 assign wire12835 = ( n_n526  &  n_n535  &  wire18 ) | ( n_n522  &  n_n535  &  wire18 ) ;
 assign wire12838 = ( n_n4940 ) | ( n_n4939 ) | ( wire342 ) ;
 assign wire12839 = ( wire341 ) | ( wire362 ) ;
 assign wire12841 = ( wire59 ) | ( wire12166 ) | ( wire180 ) | ( n_n4971 ) ;
 assign wire12843 = ( n_n4938 ) | ( n_n4933 ) | ( wire12835 ) | ( wire12841 ) ;
 assign wire12844 = ( wire12833 ) | ( wire12834 ) | ( wire12838 ) | ( wire12839 ) ;
 assign wire12845 = ( wire21  &  n_n509  &  n_n195 ) | ( wire11  &  n_n509  &  n_n195 ) ;
 assign wire12848 = ( n_n4983 ) | ( n_n4984 ) | ( wire12845 ) ;
 assign wire12849 = ( n_n4993 ) | ( n_n4994 ) | ( wire134 ) | ( n_n4986 ) ;
 assign wire12852 = ( wire103 ) | ( wire252 ) ;
 assign wire12853 = ( n_n4998 ) | ( wire57 ) | ( wire743 ) ;
 assign wire12854 = ( n_n4975 ) | ( n_n4999 ) | ( n_n4981 ) | ( n_n5002 ) ;
 assign wire12857 = ( n_n4973 ) | ( n_n801 ) | ( wire11809 ) | ( wire12854 ) ;
 assign wire12858 = ( wire12848 ) | ( wire12849 ) | ( wire12852 ) | ( wire12853 ) ;
 assign wire12859 = ( n_n482  &  n_n522  &  wire17 ) | ( n_n482  &  wire17  &  n_n530 ) ;
 assign wire12862 = ( n_n4913 ) | ( n_n4914 ) | ( n_n4915 ) | ( wire12859 ) ;
 assign wire12875 = ( _1120 ) | ( n_n65  &  wire15  &  n_n518 ) ;
 assign wire12883 = ( i_9_  &  n_n526  &  n_n130  &  n_n500 ) | ( (~ i_9_)  &  n_n526  &  n_n130  &  n_n500 ) ;
 assign wire12888 = ( n_n5167 ) | ( n_n5162 ) | ( wire168 ) ;
 assign wire12889 = ( n_n5163 ) | ( n_n5159 ) | ( wire287 ) | ( n_n5169 ) ;
 assign wire12892 = ( n_n5142 ) | ( n_n5144 ) | ( wire679 ) ;
 assign wire12893 = ( n_n5150 ) | ( n_n5149 ) | ( wire407 ) ;
 assign wire12904 = ( i_9_  &  n_n473  &  n_n528  &  n_n195 ) | ( (~ i_9_)  &  n_n473  &  n_n528  &  n_n195 ) ;
 assign wire12909 = ( wire25  &  n_n535  &  n_n130 ) | ( wire15  &  n_n535  &  n_n130 ) ;
 assign wire12914 = ( n_n5079 ) | ( n_n5083 ) | ( n_n5080 ) | ( wire209 ) ;
 assign wire12917 = ( i_9_  &  n_n522  &  n_n535  &  n_n130 ) | ( (~ i_9_)  &  n_n522  &  n_n535  &  n_n130 ) ;
 assign wire12921 = ( n_n5129 ) | ( n_n5120 ) | ( wire336 ) ;
 assign wire12922 = ( n_n5127 ) | ( n_n5128 ) | ( wire414 ) | ( n_n5122 ) ;
 assign wire12924 = ( n_n524  &  n_n518  &  wire12 ) | ( n_n518  &  n_n528  &  wire12 ) ;
 assign wire12925 = ( n_n5107 ) | ( wire122 ) | ( n_n5108 ) ;
 assign wire12926 = ( n_n5112 ) | ( n_n5086 ) | ( n_n5087 ) | ( n_n5088 ) ;
 assign wire12931 = ( n_n522  &  wire18  &  n_n500 ) | ( n_n520  &  wire18  &  n_n500 ) ;
 assign wire12934 = ( n_n5016 ) | ( n_n5013 ) | ( n_n5007 ) | ( wire12931 ) ;
 assign wire12935 = ( n_n522  &  n_n491  &  wire18 ) | ( n_n491  &  n_n524  &  wire18 ) ;
 assign wire12936 = ( n_n491  &  wire11  &  n_n195 ) | ( n_n491  &  n_n195  &  wire23 ) ;
 assign wire12939 = ( n_n5029 ) | ( wire253 ) | ( wire12936 ) ;
 assign wire12940 = ( n_n482  &  n_n526  &  wire18 ) | ( n_n482  &  wire18  &  n_n530 ) ;
 assign wire12941 = ( wire15  &  n_n482  &  n_n195 ) | ( n_n482  &  wire22  &  n_n195 ) ;
 assign wire12943 = ( n_n5043 ) | ( n_n5044 ) | ( wire12940 ) ;
 assign wire12946 = ( wire12934 ) | ( wire12939 ) | ( _24803 ) ;
 assign wire12949 = ( wire25  &  n_n65  &  n_n491 ) | ( n_n65  &  n_n491  &  wire20 ) ;
 assign wire12952 = ( n_n5277 ) | ( n_n5280 ) | ( n_n5283 ) | ( wire12371 ) ;
 assign wire12953 = ( n_n65  &  wire21  &  n_n509 ) | ( n_n65  &  wire21  &  n_n500 ) ;
 assign wire12954 = ( wire19  &  n_n522  &  n_n509 ) | ( wire19  &  n_n509  &  n_n520 ) ;
 assign wire12958 = ( n_n5260 ) | ( n_n5253 ) | ( wire12954 ) ;
 assign wire12960 = ( wire77 ) | ( wire446 ) | ( wire205 ) | ( wire12953 ) ;
 assign wire12961 = ( n_n5255 ) | ( wire433 ) | ( n_n1521 ) | ( wire12958 ) ;
 assign wire12963 = ( n_n65  &  n_n464  &  wire20 ) | ( n_n65  &  n_n464  &  wire23 ) ;
 assign wire12972 = ( n_n473  &  n_n65  &  wire22 ) | ( n_n473  &  n_n65  &  wire23 ) ;
 assign wire12976 = ( n_n65  &  n_n482  &  wire21 ) | ( n_n65  &  n_n482  &  wire11 ) ;
 assign wire12978 = ( n_n5291 ) | ( n_n5292 ) | ( n_n5298 ) ;
 assign wire12979 = ( n_n5288 ) | ( n_n5286 ) | ( wire12976 ) ;
 assign wire12981 = ( n_n5290 ) | ( n_n5289 ) | ( wire12978 ) | ( wire12979 ) ;
 assign wire12984 = ( n_n632 ) | ( n_n662 ) | ( n_n661 ) | ( wire12981 ) ;
 assign wire12985 = ( n_n464  &  wire11  &  n_n130 ) | ( n_n464  &  n_n130  &  wire23 ) ;
 assign wire12986 = ( wire15  &  n_n464  &  n_n130 ) | ( n_n464  &  wire21  &  n_n130 ) ;
 assign wire12988 = ( wire452 ) | ( wire12985 ) ;
 assign wire12989 = ( wire761 ) | ( wire12986 ) | ( _24874 ) ;
 assign wire12991 = ( wire112 ) | ( n_n5189 ) | ( n_n5190 ) ;
 assign wire12992 = ( n_n5188 ) | ( n_n5194 ) | ( wire453 ) | ( n_n5192 ) ;
 assign wire12996 = ( n_n5177 ) | ( n_n5172 ) | ( wire44 ) | ( n_n5176 ) ;
 assign wire12998 = ( wire12988 ) | ( wire12989 ) | ( wire12991 ) | ( wire12992 ) ;
 assign wire13003 = ( n_n526  &  wire13  &  n_n535 ) | ( n_n522  &  wire13  &  n_n535 ) ;
 assign wire13005 = ( n_n4445 ) | ( n_n4446 ) | ( wire128 ) ;
 assign wire13006 = ( wire368 ) | ( n_n4447 ) | ( wire13003 ) ;
 assign wire13008 = ( n_n464  &  wire16  &  n_n532 ) | ( n_n464  &  wire16  &  n_n528 ) ;
 assign wire13013 = ( n_n4436 ) | ( n_n4443 ) | ( n_n4428 ) | ( n_n4427 ) ;
 assign wire13015 = ( wire233 ) | ( wire234 ) | ( wire37 ) | ( wire13008 ) ;
 assign wire13022 = ( wire25  &  n_n455  &  n_n500 ) | ( n_n455  &  wire24  &  n_n500 ) ;
 assign wire13025 = ( wire70 ) | ( wire13022 ) ;
 assign wire13026 = ( n_n4487 ) | ( wire66 ) | ( n_n4492 ) | ( n_n4486 ) ;
 assign wire13027 = ( i_9_  &  n_n526  &  n_n455  &  n_n500 ) | ( (~ i_9_)  &  n_n526  &  n_n455  &  n_n500 ) ;
 assign wire13036 = ( n_n4522 ) | ( n_n4525 ) | ( n_n4505 ) | ( n_n4499 ) ;
 assign wire13044 = ( n_n2058 ) | ( _24946 ) | ( _24947 ) | ( _24948 ) ;
 assign wire13048 = ( n_n524  &  wire16  &  n_n535 ) | ( wire16  &  n_n528  &  n_n535 ) ;
 assign wire13049 = ( wire171 ) | ( wire364 ) ;
 assign wire13050 = ( n_n4313 ) | ( wire11583 ) | ( wire13048 ) ;
 assign wire13053 = ( n_n4325 ) | ( n_n4329 ) | ( n_n4334 ) | ( wire677 ) ;
 assign wire13054 = ( n_n4335 ) | ( n_n4330 ) | ( n_n4323 ) | ( wire12570 ) ;
 assign wire13057 = ( wire15  &  n_n536  &  n_n509 ) | ( n_n536  &  n_n509  &  wire23 ) ;
 assign wire13059 = ( n_n4355 ) | ( n_n4352 ) | ( n_n4351 ) | ( n_n4356 ) ;
 assign wire13060 = ( n_n4357 ) | ( n_n4358 ) | ( n_n4354 ) | ( wire13057 ) ;
 assign wire13062 = ( n_n4374 ) | ( n_n4373 ) | ( wire345 ) ;
 assign wire13063 = ( n_n4378 ) | ( n_n4361 ) | ( n_n4370 ) | ( wire423 ) ;
 assign wire13067 = ( n_n473  &  n_n522  &  wire16 ) | ( n_n473  &  wire16  &  n_n532 ) ;
 assign wire13078 = ( n_n4408 ) | ( n_n4397 ) | ( _24971 ) ;
 assign wire13085 = ( n_n4339 ) | ( n_n4344 ) | ( n_n4348 ) | ( wire156 ) ;
 assign wire13087 = ( wire13049 ) | ( wire13050 ) | ( wire13053 ) | ( wire13054 ) ;
 assign wire13090 = ( n_n473  &  wire13  &  n_n532 ) | ( n_n473  &  wire13  &  n_n530 ) ;
 assign wire13091 = ( i_9_  &  n_n473  &  n_n524  &  n_n455 ) | ( (~ i_9_)  &  n_n473  &  n_n524  &  n_n455 ) ;
 assign wire13093 = ( n_n473  &  wire13  &  n_n528 ) | ( n_n473  &  wire13  &  n_n520 ) ;
 assign wire13095 = ( n_n4544 ) | ( n_n4541 ) | ( wire13093 ) ;
 assign wire13096 = ( n_n4548 ) | ( wire13091 ) | ( _25076 ) ;
 assign wire13104 = ( n_n522  &  wire10  &  n_n535 ) | ( wire10  &  n_n528  &  n_n535 ) ;
 assign wire13105 = ( n_n4570 ) | ( n_n4569 ) | ( wire91 ) ;
 assign wire13108 = ( n_n4571 ) | ( n_n4582 ) | ( wire13104 ) ;
 assign wire13113 = ( _25047 ) | ( wire22  &  n_n390  &  n_n509 ) ;
 assign wire13114 = ( wire465 ) | ( wire12519 ) | ( _25048 ) ;
 assign wire13117 = ( n_n4639 ) | ( n_n4642 ) | ( n_n4632 ) ;
 assign wire13118 = ( n_n4637 ) | ( n_n4638 ) | ( wire190 ) ;
 assign wire13119 = ( n_n4616 ) | ( n_n4629 ) | ( n_n4630 ) | ( n_n4619 ) ;
 assign wire13120 = ( n_n4617 ) | ( n_n4634 ) | ( n_n4628 ) | ( n_n4640 ) ;
 assign wire13126 = ( n_n464  &  wire13  &  n_n528 ) | ( n_n464  &  wire13  &  n_n530 ) ;
 assign wire13127 = ( n_n4561 ) | ( n_n4532 ) | ( n_n4529 ) | ( wire724 ) ;
 assign wire13128 = ( n_n4536 ) | ( wire13090 ) | ( wire13126 ) ;
 assign wire13132 = ( n_n3875 ) | ( wire13095 ) | ( wire13096 ) | ( wire13127 ) ;
 assign wire13140 = ( n_n5305 ) | ( n_n5293 ) | ( n_n5297 ) ;
 assign wire13141 = ( n_n5296 ) | ( n_n5284 ) | ( wire13140 ) ;
 assign wire13144 = ( n_n562 ) | ( n_n561 ) | ( n_n563 ) | ( wire13141 ) ;
 assign wire13146 = ( n_n543 ) | ( wire12629 ) | ( wire12630 ) | ( wire13144 ) ;
 assign wire13149 = ( n_n4767 ) | ( n_n4764 ) | ( n_n4766 ) ;
 assign wire13151 = ( i_9_  &  n_n473  &  n_n325  &  n_n530 ) | ( (~ i_9_)  &  n_n473  &  n_n325  &  n_n530 ) ;
 assign wire13153 = ( n_n4790 ) | ( n_n4798 ) | ( wire158 ) ;
 assign wire13154 = ( wire179 ) | ( n_n4799 ) | ( wire13151 ) ;
 assign wire13171 = ( n_n4857 ) | ( n_n4862 ) | ( n_n4856 ) | ( wire40 ) ;
 assign wire13172 = ( n_n518  &  wire21  &  n_n260 ) | ( n_n518  &  wire11  &  n_n260 ) ;
 assign wire13174 = ( n_n4849 ) | ( n_n4850 ) | ( n_n4848 ) | ( wire13172 ) ;
 assign wire13182 = ( n_n482  &  n_n526  &  wire14 ) | ( n_n482  &  wire14  &  n_n528 ) ;
 assign wire13183 = ( n_n482  &  wire24  &  n_n325 ) | ( n_n482  &  n_n325  &  wire20 ) ;
 assign wire13185 = ( n_n4776 ) | ( n_n4774 ) | ( n_n4775 ) | ( wire13183 ) ;
 assign wire13187 = ( wire447 ) | ( wire13149 ) | ( wire13153 ) | ( wire13154 ) ;
 assign wire13193 = ( n_n4885 ) | ( n_n4882 ) | ( wire330 ) ;
 assign wire13194 = ( n_n4883 ) | ( wire260 ) | ( n_n4880 ) | ( n_n4889 ) ;
 assign wire13198 = ( n_n4898 ) | ( n_n4895 ) | ( wire49 ) ;
 assign wire13199 = ( n_n4894 ) | ( wire96 ) | ( n_n4897 ) | ( n_n4891 ) ;
 assign wire13213 = ( wire31 ) | ( n_n1592 ) | ( wire42 ) | ( _25642 ) ;
 assign wire13215 = ( n_n522  &  n_n535  &  wire18 ) | ( n_n535  &  n_n520  &  wire18 ) ;
 assign wire13216 = ( i_9_  &  n_n535  &  n_n195  &  n_n530 ) | ( (~ i_9_)  &  n_n535  &  n_n195  &  n_n530 ) ;
 assign wire13217 = ( n_n518  &  wire11  &  n_n195 ) | ( n_n518  &  wire24  &  n_n195 ) ;
 assign wire13218 = ( i_9_  &  n_n518  &  n_n195  &  n_n530 ) | ( (~ i_9_)  &  n_n518  &  n_n195  &  n_n530 ) ;
 assign wire13222 = ( n_n4959 ) | ( n_n4960 ) | ( wire771 ) | ( wire772 ) ;
 assign wire13223 = ( wire141 ) | ( wire317 ) ;
 assign wire13224 = ( n_n4967 ) | ( n_n4962 ) | ( n_n4948 ) | ( n_n4953 ) ;
 assign wire13234 = ( wire13193 ) | ( wire13194 ) | ( wire13198 ) | ( wire13199 ) ;
 assign wire13237 = ( i_9_  &  n_n509  &  n_n325  &  n_n528 ) | ( (~ i_9_)  &  n_n509  &  n_n325  &  n_n528 ) ;
 assign wire13239 = ( n_n4737 ) | ( n_n4738 ) | ( n_n4732 ) | ( wire767 ) ;
 assign wire13240 = ( wire374 ) | ( n_n4743 ) | ( wire13237 ) ;
 assign wire13248 = ( wire25  &  n_n518  &  n_n325 ) | ( n_n518  &  wire21  &  n_n325 ) ;
 assign wire13251 = ( n_n4708 ) | ( n_n4716 ) | ( wire13248 ) ;
 assign wire13256 = ( i_9_  &  n_n473  &  n_n532  &  n_n390 ) | ( (~ i_9_)  &  n_n473  &  n_n532  &  n_n390 ) ;
 assign wire13259 = ( n_n4658 ) | ( wire775 ) | ( wire13256 ) ;
 assign wire13260 = ( n_n4664 ) | ( n_n4662 ) | ( wire72 ) | ( n_n4657 ) ;
 assign wire13261 = ( i_9_  &  n_n473  &  n_n390  &  n_n528 ) | ( (~ i_9_)  &  n_n473  &  n_n390  &  n_n528 ) ;
 assign wire13263 = ( n_n4674 ) | ( n_n4673 ) | ( wire157 ) ;
 assign wire13264 = ( wire80 ) | ( n_n4680 ) | ( wire13261 ) ;
 assign wire13265 = ( n_n526  &  n_n464  &  wire10 ) | ( n_n524  &  n_n464  &  wire10 ) ;
 assign wire13266 = ( wire15  &  n_n464  &  n_n390 ) | ( n_n464  &  wire11  &  n_n390 ) ;
 assign wire13268 = ( n_n4683 ) | ( wire81 ) | ( n_n4684 ) | ( wire13266 ) ;
 assign wire13272 = ( wire22  &  n_n325  &  n_n500 ) | ( wire24  &  n_n325  &  n_n500 ) ;
 assign wire13274 = ( n_n4754 ) | ( n_n4749 ) | ( wire47 ) ;
 assign wire13277 = ( wire11836 ) | ( wire11837 ) | ( wire13239 ) | ( wire13240 ) ;
 assign wire13283 = ( n_n5142 ) | ( n_n5135 ) | ( wire407 ) ;
 assign wire13284 = ( n_n5150 ) | ( wire76 ) | ( n_n5140 ) | ( n_n5143 ) ;
 assign wire13285 = ( n_n491  &  wire20  &  n_n130 ) | ( n_n491  &  n_n130  &  wire23 ) ;
 assign wire13287 = ( wire358 ) | ( wire168 ) ;
 assign wire13288 = ( wire196 ) | ( n_n5151 ) | ( wire13285 ) ;
 assign wire13291 = ( n_n473  &  n_n532  &  wire12 ) | ( n_n473  &  n_n534  &  wire12 ) ;
 assign wire13292 = ( n_n5174 ) | ( n_n5183 ) | ( wire113 ) ;
 assign wire13293 = ( n_n5181 ) | ( n_n5182 ) | ( wire732 ) | ( wire13291 ) ;
 assign wire13294 = ( n_n482  &  n_n526  &  wire12 ) | ( n_n482  &  n_n532  &  wire12 ) ;
 assign wire13296 = ( wire254 ) | ( wire332 ) ;
 assign wire13297 = ( n_n5169 ) | ( wire33 ) | ( wire13294 ) ;
 assign wire13298 = ( i_9_  &  n_n473  &  n_n522  &  n_n130 ) | ( (~ i_9_)  &  n_n473  &  n_n522  &  n_n130 ) ;
 assign wire13301 = ( n_n5187 ) | ( n_n5196 ) | ( wire13298 ) ;
 assign wire13303 = ( n_n5195 ) | ( n_n2670 ) | ( n_n5192 ) | ( wire13301 ) ;
 assign wire13304 = ( wire13292 ) | ( wire13293 ) | ( wire13296 ) | ( wire13297 ) ;
 assign wire13308 = ( n_n5113 ) | ( n_n5108 ) | ( _25791 ) ;
 assign wire13310 = ( n_n518  &  n_n532  &  wire12 ) | ( n_n518  &  wire12  &  n_n530 ) ;
 assign wire13311 = ( i_9_  &  n_n528  &  n_n535  &  n_n130 ) | ( (~ i_9_)  &  n_n528  &  n_n535  &  n_n130 ) ;
 assign wire13313 = ( wire289 ) | ( wire279 ) ;
 assign wire13314 = ( n_n5099 ) | ( n_n5085 ) | ( wire13310 ) ;
 assign wire13317 = ( n_n5106 ) | ( n_n5095 ) | ( wire144 ) | ( wire13311 ) ;
 assign wire13318 = ( wire28 ) | ( wire13308 ) | ( wire13313 ) | ( wire13314 ) ;
 assign wire13320 = ( n_n509  &  n_n528  &  wire12 ) | ( n_n528  &  wire12  &  n_n500 ) ;
 assign wire13334 = ( n_n5276 ) | ( n_n5281 ) | ( n_n5277 ) | ( wire218 ) ;
 assign wire13350 = ( wire19  &  n_n524  &  n_n535 ) | ( wire19  &  n_n528  &  n_n535 ) ;
 assign wire13351 = ( wire19  &  n_n518  &  n_n528 ) | ( wire19  &  n_n518  &  n_n520 ) ;
 assign wire13352 = ( n_n65  &  n_n518  &  wire21 ) | ( n_n65  &  n_n518  &  wire20 ) ;
 assign wire13354 = ( wire181 ) | ( wire13351 ) ;
 assign wire13355 = ( wire87 ) | ( wire182 ) | ( wire13352 ) ;
 assign wire13359 = ( n_n5210 ) | ( wire384 ) | ( n_n5209 ) ;
 assign wire13360 = ( n_n5204 ) | ( n_n5201 ) | ( n_n5207 ) | ( n_n5208 ) ;
 assign wire13361 = ( n_n5220 ) | ( n_n5203 ) | ( n_n5211 ) | ( n_n5205 ) ;
 assign wire13368 = ( i_9_  &  n_n65  &  n_n482  &  n_n532 ) | ( (~ i_9_)  &  n_n65  &  n_n482  &  n_n532 ) ;
 assign wire13370 = ( n_n5294 ) | ( n_n5299 ) | ( n_n5287 ) | ( n_n5288 ) ;
 assign wire13372 = ( n_n5292 ) | ( wire441 ) | ( wire13368 ) | ( wire13370 ) ;
 assign wire13378 = ( n_n509  &  n_n528  &  wire18 ) | ( n_n509  &  n_n520  &  wire18 ) ;
 assign wire13380 = ( n_n4991 ) | ( n_n4996 ) | ( n_n4992 ) | ( n_n4995 ) ;
 assign wire13381 = ( n_n4999 ) | ( wire103 ) | ( wire13378 ) ;
 assign wire13384 = ( wire393 ) | ( wire343 ) ;
 assign wire13385 = ( n_n5004 ) | ( wire136 ) | ( n_n5013 ) | ( n_n5008 ) ;
 assign wire13390 = ( n_n5081 ) | ( n_n5082 ) | ( n_n5084 ) | ( n_n5079 ) ;
 assign wire13391 = ( n_n473  &  wire21  &  n_n195 ) | ( n_n473  &  wire11  &  n_n195 ) ;
 assign wire13392 = ( n_n5067 ) | ( n_n5057 ) | ( n_n5058 ) ;
 assign wire13393 = ( n_n5061 ) | ( wire160 ) | ( wire669 ) ;
 assign wire13394 = ( n_n5073 ) | ( n_n5074 ) | ( n_n5072 ) | ( wire13391 ) ;
 assign wire13397 = ( n_n1952 ) | ( n_n789 ) | ( wire13394 ) ;
 assign wire13398 = ( wire90 ) | ( wire13390 ) | ( wire13392 ) | ( wire13393 ) ;
 assign wire13399 = ( i_9_  &  n_n491  &  n_n524  &  n_n195 ) | ( (~ i_9_)  &  n_n491  &  n_n524  &  n_n195 ) ;
 assign wire13400 = ( i_9_  &  n_n491  &  n_n528  &  n_n195 ) | ( (~ i_9_)  &  n_n491  &  n_n528  &  n_n195 ) ;
 assign wire13401 = ( n_n473  &  n_n534  &  wire18 ) | ( n_n473  &  n_n528  &  wire18 ) ;
 assign wire13404 = ( n_n5050 ) | ( n_n5049 ) | ( wire13401 ) ;
 assign wire13405 = ( n_n5045 ) | ( wire166 ) | ( n_n5051 ) | ( n_n5044 ) ;
 assign wire13406 = ( n_n482  &  n_n526  &  wire18 ) | ( n_n482  &  n_n528  &  wire18 ) ;
 assign wire13408 = ( i_9_  &  n_n482  &  n_n524  &  n_n195 ) | ( (~ i_9_)  &  n_n482  &  n_n524  &  n_n195 ) ;
 assign wire13409 = ( n_n5034 ) | ( n_n5041 ) | ( wire13406 ) ;
 assign wire13410 = ( wire50 ) | ( n_n5029 ) | ( wire13408 ) ;
 assign wire13411 = ( i_9_  &  n_n491  &  n_n532  &  n_n195 ) | ( (~ i_9_)  &  n_n491  &  n_n532  &  n_n195 ) ;
 assign wire13413 = ( n_n5025 ) | ( n_n5024 ) | ( wire13399 ) | ( wire13400 ) ;
 assign wire13414 = ( n_n5014 ) | ( wire13411 ) | ( wire13413 ) ;
 assign wire13415 = ( wire13404 ) | ( wire13405 ) | ( wire13409 ) | ( wire13410 ) ;
 assign wire13417 = ( i_9_  &  n_n534  &  n_n509  &  n_n195 ) | ( (~ i_9_)  &  n_n534  &  n_n509  &  n_n195 ) ;
 assign wire13422 = ( wire13380 ) | ( wire13381 ) | ( wire13384 ) | ( wire13385 ) ;
 assign wire13424 = ( wire13397 ) | ( wire13398 ) | ( wire13414 ) | ( wire13415 ) ;
 assign wire13425 = ( i_9_  &  n_n522  &  n_n455  &  n_n535 ) | ( (~ i_9_)  &  n_n522  &  n_n455  &  n_n535 ) ;
 assign wire13428 = ( wire233 ) | ( wire236 ) ;
 assign wire13429 = ( n_n4440 ) | ( n_n4434 ) | ( n_n4432 ) | ( wire98 ) ;
 assign wire13430 = ( wire25  &  n_n455  &  n_n535 ) | ( wire22  &  n_n455  &  n_n535 ) ;
 assign wire13431 = ( n_n4448 ) | ( n_n4447 ) | ( wire421 ) ;
 assign wire13432 = ( n_n4445 ) | ( n_n4444 ) | ( n_n4446 ) | ( wire13430 ) ;
 assign wire13436 = ( n_n4430 ) | ( n_n4425 ) | ( n_n4423 ) | ( n_n4429 ) ;
 assign wire13437 = ( n_n4421 ) | ( wire84 ) | ( n_n4424 ) | ( n_n4428 ) ;
 assign wire13438 = ( wire13436 ) | ( wire13437 ) ;
 assign wire13439 = ( wire13428 ) | ( wire13429 ) | ( wire13431 ) | ( wire13432 ) ;
 assign wire13443 = ( n_n524  &  wire10  &  n_n509 ) | ( wire10  &  n_n509  &  n_n528 ) ;
 assign wire13448 = ( wire22  &  n_n390  &  n_n535 ) | ( n_n390  &  n_n535  &  wire20 ) ;
 assign wire13450 = ( n_n4575 ) | ( n_n4584 ) | ( n_n4586 ) | ( n_n4583 ) ;
 assign wire13454 = ( i_9_  &  n_n526  &  n_n491  &  n_n390 ) | ( (~ i_9_)  &  n_n526  &  n_n491  &  n_n390 ) ;
 assign wire13455 = ( i_9_  &  n_n482  &  n_n390  &  n_n534 ) | ( (~ i_9_)  &  n_n482  &  n_n390  &  n_n534 ) ;
 assign wire13457 = ( wire140 ) | ( wire13455 ) ;
 assign wire13458 = ( n_n4652 ) | ( n_n4643 ) | ( n_n4642 ) | ( wire13454 ) ;
 assign wire13459 = ( n_n491  &  wire10  &  n_n532 ) | ( n_n491  &  wire10  &  n_n528 ) ;
 assign wire13461 = ( wire22  &  n_n390  &  n_n500 ) | ( n_n390  &  wire23  &  n_n500 ) ;
 assign wire13462 = ( wire118 ) | ( n_n4633 ) | ( n_n4630 ) ;
 assign wire13463 = ( wire401 ) | ( wire13459 ) ;
 assign wire13465 = ( n_n4616 ) | ( wire465 ) | ( n_n4627 ) | ( wire12546 ) ;
 assign wire13470 = ( n_n4568 ) | ( wire455 ) | ( wire783 ) ;
 assign wire13471 = ( n_n4560 ) | ( n_n4569 ) | ( wire471 ) | ( wire91 ) ;
 assign wire13473 = ( n_n473  &  n_n522  &  wire13 ) | ( n_n473  &  wire13  &  n_n520 ) ;
 assign wire13474 = ( n_n4554 ) | ( n_n4541 ) | ( wire416 ) ;
 assign wire13475 = ( n_n4545 ) | ( wire13091 ) | ( wire13473 ) ;
 assign wire13479 = ( n_n4537 ) | ( n_n4527 ) | ( n_n4534 ) | ( wire11532 ) ;
 assign wire13481 = ( wire13470 ) | ( wire13471 ) | ( wire13474 ) | ( wire13475 ) ;
 assign wire13487 = ( n_n4482 ) | ( n_n4489 ) | ( wire199 ) ;
 assign wire13488 = ( n_n4487 ) | ( n_n4478 ) | ( wire70 ) | ( n_n4486 ) ;
 assign wire13494 = ( wire66 ) | ( n_n4496 ) | ( n_n4499 ) | ( n_n4493 ) ;
 assign wire13495 = ( _930 ) | ( n_n526  &  n_n491  &  wire13 ) ;
 assign wire13497 = ( n_n4502 ) | ( wire308 ) | ( n_n4501 ) ;
 assign wire13501 = ( n_n4247 ) | ( n_n4246 ) | ( n_n3152 ) | ( wire13495 ) ;
 assign wire13502 = ( wire13494 ) | ( wire13497 ) | ( _25438 ) ;
 assign wire13503 = ( n_n518  &  wire21  &  n_n455 ) | ( n_n518  &  n_n455  &  wire23 ) ;
 assign wire13504 = ( i_9_  &  n_n522  &  n_n518  &  n_n455 ) | ( (~ i_9_)  &  n_n522  &  n_n518  &  n_n455 ) ;
 assign wire13505 = ( n_n4464 ) | ( n_n4463 ) | ( wire13503 ) ;
 assign wire13506 = ( n_n4476 ) | ( wire13504 ) | ( _25401 ) ;
 assign wire13508 = ( i_9_  &  n_n536  &  n_n534  &  n_n509 ) | ( (~ i_9_)  &  n_n536  &  n_n534  &  n_n509 ) ;
 assign wire13509 = ( wire67 ) | ( wire156 ) ;
 assign wire13510 = ( n_n4337 ) | ( wire53 ) | ( wire13508 ) ;
 assign wire13513 = ( n_n526  &  wire16  &  n_n518 ) | ( n_n526  &  wire16  &  n_n535 ) ;
 assign wire13515 = ( wire283 ) | ( n_n4334 ) | ( wire677 ) ;
 assign wire13516 = ( n_n4316 ) | ( n_n4313 ) | ( wire13513 ) ;
 assign wire13521 = ( _25369 ) | ( n_n536  &  wire20  &  n_n500 ) ;
 assign wire13522 = ( n_n4381 ) | ( wire423 ) | ( n_n4375 ) | ( wire12449 ) ;
 assign wire13523 = ( wire22  &  n_n536  &  n_n509 ) | ( n_n536  &  n_n509  &  wire20 ) ;
 assign wire13524 = ( n_n4355 ) | ( n_n4352 ) | ( n_n4351 ) | ( n_n4356 ) ;
 assign wire13525 = ( n_n4350 ) | ( n_n4349 ) | ( n_n4348 ) | ( wire13523 ) ;
 assign wire13526 = ( wire25  &  n_n473  &  n_n536 ) | ( n_n473  &  wire22  &  n_n536 ) ;
 assign wire13534 = ( n_n482  &  wire22  &  n_n536 ) | ( n_n482  &  wire21  &  n_n536 ) ;
 assign wire13535 = ( n_n482  &  n_n526  &  wire16 ) | ( n_n482  &  n_n522  &  wire16 ) ;
 assign wire13538 = ( n_n4396 ) | ( n_n4405 ) | ( n_n4406 ) | ( wire13535 ) ;
 assign wire13541 = ( wire22  &  n_n536  &  n_n500 ) | ( n_n536  &  wire11  &  n_n500 ) ;
 assign wire13542 = ( n_n524  &  wire16  &  n_n500 ) | ( wire16  &  n_n534  &  n_n500 ) ;
 assign wire13543 = ( n_n4361 ) | ( n_n4359 ) | ( wire13541 ) ;
 assign wire13546 = ( wire13521 ) | ( wire13522 ) | ( wire13524 ) | ( wire13525 ) ;
 assign wire13550 = ( n_n4451 ) | ( n_n4462 ) | ( wire12471 ) | ( wire13425 ) ;
 assign wire13552 = ( wire13487 ) | ( wire13488 ) | ( wire13505 ) | ( wire13506 ) ;
 assign wire13559 = ( wire19  &  n_n464  &  n_n534 ) | ( wire19  &  n_n464  &  n_n528 ) ;
 assign wire13560 = ( n_n65  &  wire22  &  n_n464 ) | ( n_n65  &  n_n464  &  wire11 ) ;
 assign wire13561 = ( wire19  &  n_n526  &  n_n464 ) | ( wire19  &  n_n464  &  n_n532 ) ;
 assign wire13562 = ( i_9_  &  n_n65  &  n_n464  &  n_n520 ) | ( (~ i_9_)  &  n_n65  &  n_n464  &  n_n520 ) ;
 assign wire13577 = ( wire15  &  n_n509  &  n_n130 ) | ( wire11  &  n_n509  &  n_n130 ) ;
 assign wire13601 = ( n_n482  &  n_n534  &  wire18 ) | ( n_n482  &  wire18  &  n_n530 ) ;
 assign wire13606 = ( n_n5017 ) | ( n_n5037 ) | ( n_n5015 ) | ( n_n5056 ) ;
 assign wire13607 = ( n_n5047 ) | ( n_n5020 ) | ( n_n5021 ) | ( wire13601 ) ;
 assign wire13611 = ( n_n5156 ) | ( n_n5191 ) | ( n_n5175 ) | ( n_n5177 ) ;
 assign wire13612 = ( n_n5190 ) | ( wire107 ) | ( n_n5194 ) | ( n_n5213 ) ;
 assign wire13616 = ( wire13606 ) | ( wire13607 ) | ( wire13611 ) | ( wire13612 ) ;
 assign wire13617 = ( n_n3926 ) | ( n_n3924 ) | ( n_n3923 ) | ( n_n3928 ) ;
 assign wire13638 = ( wire15  &  n_n482  &  n_n325 ) | ( wire15  &  n_n509  &  n_n325 ) ;
 assign wire13648 = ( n_n526  &  wire10  &  n_n535 ) | ( n_n522  &  wire10  &  n_n535 ) ;
 assign wire13650 = ( n_n4570 ) | ( n_n4557 ) | ( n_n4553 ) | ( n_n4558 ) ;
 assign wire13651 = ( n_n4551 ) | ( n_n4552 ) | ( n_n4549 ) | ( wire13648 ) ;
 assign wire13656 = ( n_n4617 ) | ( n_n4637 ) | ( n_n4613 ) | ( n_n4602 ) ;
 assign wire13657 = ( n_n4611 ) | ( n_n4639 ) | ( n_n4608 ) | ( wire139 ) ;
 assign wire13660 = ( wire15  &  n_n491  &  n_n455 ) | ( n_n491  &  n_n455  &  wire24 ) ;
 assign wire13662 = ( n_n4521 ) | ( n_n4544 ) | ( n_n4520 ) ;
 assign wire13663 = ( n_n4504 ) | ( n_n4535 ) | ( wire13660 ) ;
 assign wire13666 = ( wire13650 ) | ( wire13651 ) | ( wire13656 ) | ( wire13657 ) ;
 assign wire13670 = ( n_n526  &  wire13  &  n_n509 ) | ( wire13  &  n_n534  &  n_n509 ) ;
 assign wire13673 = ( n_n4459 ) | ( n_n4420 ) | ( n_n4410 ) | ( wire13670 ) ;
 assign wire13681 = ( n_n3936 ) | ( wire13679 ) | ( _25967 ) | ( _25975 ) ;
 assign wire13683 = ( wire13616 ) | ( wire13617 ) | ( wire13681 ) ;
 assign wire13689 = ( n_n4339 ) | ( n_n4401 ) | ( n_n4314 ) | ( n_n4389 ) ;
 assign wire13690 = ( n_n4369 ) | ( n_n4381 ) | ( n_n4340 ) | ( wire280 ) ;
 assign wire13694 = ( wire25  &  n_n491  &  n_n130 ) | ( wire25  &  n_n130  &  n_n500 ) ;
 assign wire13696 = ( n_n5142 ) | ( n_n5107 ) | ( n_n5130 ) | ( n_n5123 ) ;
 assign wire13697 = ( n_n5101 ) | ( n_n5110 ) | ( n_n5156 ) | ( wire13694 ) ;
 assign wire13698 = ( i_9_  &  n_n65  &  n_n518  &  n_n520 ) | ( (~ i_9_)  &  n_n65  &  n_n518  &  n_n520 ) ;
 assign wire13703 = ( n_n5182 ) | ( n_n5173 ) | ( n_n5165 ) | ( n_n5230 ) ;
 assign wire13704 = ( n_n5166 ) | ( n_n5163 ) | ( n_n5214 ) | ( wire13698 ) ;
 assign wire13713 = ( n_n5305 ) | ( n_n5302 ) | ( n_n5303 ) ;
 assign wire13717 = ( n_n473  &  n_n195  &  wire23 ) | ( n_n464  &  n_n195  &  wire23 ) ;
 assign wire13719 = ( n_n5085 ) | ( n_n5072 ) | ( n_n5082 ) | ( n_n5075 ) ;
 assign wire13720 = ( n_n5096 ) | ( n_n5099 ) | ( n_n5065 ) | ( wire13717 ) ;
 assign wire13725 = ( n_n4996 ) | ( n_n4987 ) | ( n_n5006 ) ;
 assign wire13726 = ( n_n4994 ) | ( n_n5056 ) | ( n_n5002 ) | ( n_n5053 ) ;
 assign wire13735 = ( n_n4437 ) | ( n_n4409 ) | ( n_n4487 ) | ( n_n4472 ) ;
 assign wire13736 = ( n_n4484 ) | ( n_n4462 ) | ( n_n4428 ) | ( wire403 ) ;
 assign wire13741 = ( n_n4539 ) | ( n_n4544 ) | ( n_n4533 ) | ( n_n4507 ) ;
 assign wire13742 = ( n_n4532 ) | ( n_n4499 ) | ( n_n4545 ) | ( wire471 ) ;
 assign wire13755 = ( wire25  &  n_n325  &  n_n535 ) | ( wire24  &  n_n325  &  n_n535 ) ;
 assign wire13756 = ( n_n526  &  n_n491  &  wire10 ) | ( n_n491  &  wire10  &  n_n528 ) ;
 assign wire13765 = ( n_n522  &  n_n518  &  wire18 ) | ( n_n518  &  wire18  &  n_n530 ) ;
 assign wire13776 = ( n_n518  &  wire11  &  n_n260 ) | ( n_n518  &  n_n260  &  wire20 ) ;
 assign wire13777 = ( n_n482  &  n_n526  &  wire17 ) | ( n_n526  &  n_n509  &  wire17 ) ;
 assign wire13779 = ( n_n4900 ) | ( n_n4849 ) | ( n_n4896 ) ;
 assign wire13788 = ( n_n4784 ) | ( n_n4783 ) | ( wire292 ) ;
 assign wire13789 = ( n_n4782 ) | ( wire131 ) | ( n_n4789 ) | ( n_n4788 ) ;
 assign wire13790 = ( _664 ) | ( n_n325  &  wire23  &  n_n500 ) ;
 assign wire13791 = ( _26476 ) | ( n_n491  &  n_n532  &  wire14 ) ;
 assign wire13792 = ( n_n4760 ) | ( n_n4758 ) | ( wire164 ) ;
 assign wire13798 = ( n_n473  &  n_n526  &  wire14 ) | ( n_n473  &  n_n532  &  wire14 ) ;
 assign wire13800 = ( n_n4801 ) | ( n_n4802 ) | ( wire380 ) ;
 assign wire13807 = ( i_9_  &  n_n518  &  n_n534  &  n_n260 ) | ( (~ i_9_)  &  n_n518  &  n_n534  &  n_n260 ) ;
 assign wire13810 = ( wire21  &  n_n509  &  n_n260 ) | ( n_n509  &  n_n260  &  wire20 ) ;
 assign wire13815 = ( wire15  &  n_n518  &  n_n260 ) | ( n_n518  &  wire24  &  n_n260 ) ;
 assign wire13816 = ( n_n526  &  n_n518  &  wire17 ) | ( n_n518  &  n_n528  &  wire17 ) ;
 assign wire13823 = ( n_n4806 ) | ( n_n4810 ) | ( n_n4805 ) | ( wire773 ) ;
 assign wire13824 = ( wire85 ) | ( n_n4807 ) | ( n_n4808 ) | ( wire12225 ) ;
 assign wire13827 = ( n_n3330 ) | ( wire13823 ) | ( wire13824 ) | ( _26515 ) ;
 assign wire13833 = ( n_n4976 ) | ( n_n4981 ) | ( wire251 ) ;
 assign wire13834 = ( n_n4988 ) | ( n_n4985 ) | ( n_n4984 ) | ( wire57 ) ;
 assign wire13836 = ( n_n4975 ) | ( n_n4968 ) | ( wire771 ) | ( wire772 ) ;
 assign wire13837 = ( n_n464  &  wire21  &  n_n260 ) | ( n_n464  &  n_n260  &  wire20 ) ;
 assign wire13840 = ( wire342 ) | ( wire13837 ) ;
 assign wire13841 = ( n_n4974 ) | ( n_n4948 ) | ( n_n4957 ) | ( n_n4971 ) ;
 assign wire13854 = ( wire25  &  n_n482  &  n_n260 ) | ( wire25  &  n_n491  &  n_n260 ) ;
 assign wire13857 = ( n_n4909 ) | ( n_n4894 ) | ( wire13854 ) ;
 assign wire13865 = ( n_n4927 ) | ( n_n4926 ) | ( n_n4925 ) | ( n_n4934 ) ;
 assign wire13866 = ( wire31 ) | ( n_n4930 ) | ( n_n4933 ) | ( n_n4931 ) ;
 assign wire13870 = ( n_n4911 ) | ( n_n4916 ) | ( n_n4918 ) | ( n_n4917 ) ;
 assign wire13872 = ( wire25  &  n_n473  &  n_n260 ) | ( n_n473  &  n_n260  &  wire23 ) ;
 assign wire13873 = ( n_n4923 ) | ( n_n4924 ) | ( n_n4937 ) | ( n_n4938 ) ;
 assign wire13874 = ( n_n4942 ) | ( wire59 ) | ( n_n4940 ) | ( wire13872 ) ;
 assign wire13877 = ( wire58 ) | ( wire13865 ) | ( wire13866 ) | ( wire13873 ) ;
 assign wire13880 = ( n_n524  &  wire14  &  n_n500 ) | ( n_n534  &  wire14  &  n_n500 ) ;
 assign wire13881 = ( wire15  &  n_n325  &  n_n500 ) | ( n_n325  &  wire20  &  n_n500 ) ;
 assign wire13883 = ( n_n4748 ) | ( n_n4747 ) | ( wire13880 ) ;
 assign wire13884 = ( n_n4756 ) | ( wire109 ) | ( wire13881 ) ;
 assign wire13885 = ( wire25  &  n_n482  &  n_n390 ) | ( n_n482  &  wire11  &  n_n390 ) ;
 assign wire13887 = ( wire140 ) | ( wire391 ) ;
 assign wire13888 = ( wire311 ) | ( n_n4654 ) | ( wire13885 ) ;
 assign wire13891 = ( n_n4669 ) | ( n_n4670 ) | ( wire72 ) ;
 assign wire13892 = ( n_n4671 ) | ( wire418 ) | ( n_n4672 ) ;
 assign wire13893 = ( n_n4673 ) | ( n_n4658 ) | ( n_n4684 ) | ( n_n4665 ) ;
 assign wire13895 = ( n_n4674 ) | ( n_n4677 ) | ( wire11855 ) | ( wire13893 ) ;
 assign wire13896 = ( wire13887 ) | ( wire13888 ) | ( wire13891 ) | ( wire13892 ) ;
 assign wire13900 = ( n_n526  &  n_n464  &  wire10 ) | ( n_n464  &  wire10  &  n_n528 ) ;
 assign wire13902 = ( n_n4690 ) | ( n_n4689 ) | ( wire442 ) ;
 assign wire13903 = ( n_n4694 ) | ( wire445 ) | ( wire13900 ) ;
 assign wire13905 = ( n_n4718 ) | ( n_n4717 ) | ( n_n4716 ) ;
 assign wire13906 = ( n_n4710 ) | ( n_n4709 ) | ( wire366 ) ;
 assign wire13910 = ( wire13897 ) | ( n_n2378 ) | ( _672 ) | ( _26451 ) ;
 assign wire13911 = ( wire13902 ) | ( wire13903 ) | ( wire13905 ) | ( wire13906 ) ;
 assign wire13913 = ( n_n4725 ) | ( n_n4726 ) | ( n_n4729 ) ;
 assign wire13914 = ( wire244 ) | ( n_n4732 ) | ( wire767 ) ;
 assign wire13915 = ( n_n4727 ) | ( wire95 ) | ( n_n4733 ) | ( n_n4736 ) ;
 assign wire13918 = ( wire13883 ) | ( wire13884 ) | ( wire13913 ) | ( wire13914 ) ;
 assign wire13919 = ( wire456 ) | ( wire13915 ) | ( wire13918 ) ;
 assign wire13920 = ( wire13895 ) | ( wire13896 ) | ( wire13910 ) | ( wire13911 ) ;
 assign wire13931 = ( n_n473  &  wire19  &  n_n528 ) | ( n_n473  &  wire19  &  n_n520 ) ;
 assign wire13932 = ( n_n473  &  wire19  &  n_n522 ) | ( n_n473  &  wire19  &  n_n524 ) ;
 assign wire13934 = ( wire459 ) | ( wire13931 ) ;
 assign wire13935 = ( n_n5320 ) | ( n_n5321 ) | ( n_n5319 ) | ( wire13932 ) ;
 assign wire13938 = ( n_n65  &  n_n482  &  wire22 ) | ( n_n65  &  n_n482  &  wire21 ) ;
 assign wire13940 = ( n_n473  &  wire19  &  n_n534 ) | ( n_n473  &  wire19  &  n_n530 ) ;
 assign wire13942 = ( n_n5306 ) | ( n_n5309 ) | ( wire13938 ) ;
 assign wire13943 = ( wire200 ) | ( wire656 ) | ( wire13940 ) ;
 assign wire13944 = ( i_9_  &  n_n65  &  n_n526  &  n_n464 ) | ( (~ i_9_)  &  n_n65  &  n_n526  &  n_n464 ) ;
 assign wire13947 = ( n_n2274 ) | ( n_n2643 ) | ( n_n5330 ) | ( wire13944 ) ;
 assign wire13948 = ( wire13934 ) | ( wire13935 ) | ( wire13942 ) | ( wire13943 ) ;
 assign wire13952 = ( n_n5222 ) | ( n_n5225 ) | ( wire385 ) | ( wire87 ) ;
 assign wire13955 = ( wire433 ) | ( n_n5250 ) | ( _26108 ) ;
 assign wire13957 = ( i_9_  &  n_n65  &  n_n524  &  n_n518 ) | ( (~ i_9_)  &  n_n65  &  n_n524  &  n_n518 ) ;
 assign wire13960 = ( n_n5244 ) | ( n_n5243 ) | ( n_n5246 ) | ( wire13957 ) ;
 assign wire13961 = ( n_n5232 ) | ( n_n5241 ) | ( wire386 ) | ( wire13960 ) ;
 assign wire13962 = ( wire13952 ) | ( wire13955 ) | ( _26110 ) ;
 assign wire13963 = ( i_9_  &  n_n65  &  n_n524  &  n_n500 ) | ( (~ i_9_)  &  n_n65  &  n_n524  &  n_n500 ) ;
 assign wire13964 = ( wire19  &  n_n528  &  n_n500 ) | ( wire19  &  n_n500  &  n_n530 ) ;
 assign wire13966 = ( n_n5270 ) | ( n_n5269 ) | ( wire13963 ) ;
 assign wire13967 = ( wire62 ) | ( wire92 ) | ( wire13964 ) ;
 assign wire13968 = ( wire218 ) | ( wire19  &  n_n526  &  n_n491 ) ;
 assign wire13969 = ( i_9_  &  n_n65  &  n_n482  &  n_n528 ) | ( (~ i_9_)  &  n_n65  &  n_n482  &  n_n528 ) ;
 assign wire13971 = ( n_n5290 ) | ( n_n5286 ) | ( n_n5289 ) ;
 assign wire13972 = ( wire441 ) | ( wire13969 ) ;
 assign wire13975 = ( wire204 ) | ( wire13966 ) | ( wire13967 ) | ( wire13968 ) ;
 assign wire13977 = ( wire13947 ) | ( wire13948 ) | ( wire13961 ) | ( wire13962 ) ;
 assign wire13978 = ( n_n473  &  n_n522  &  wire18 ) | ( n_n473  &  n_n532  &  wire18 ) ;
 assign wire13979 = ( i_9_  &  n_n473  &  n_n528  &  n_n195 ) | ( (~ i_9_)  &  n_n473  &  n_n528  &  n_n195 ) ;
 assign wire13981 = ( n_n5057 ) | ( n_n5058 ) | ( wire13978 ) ;
 assign wire13982 = ( n_n5059 ) | ( n_n5064 ) | ( wire755 ) | ( wire13979 ) ;
 assign wire13985 = ( n_n473  &  n_n534  &  wire18 ) | ( n_n482  &  n_n534  &  wire18 ) ;
 assign wire13989 = ( n_n5025 ) | ( n_n5028 ) | ( n_n5036 ) | ( wire13399 ) ;
 assign wire13990 = ( wire50 ) | ( wire231 ) | ( wire356 ) | ( wire13985 ) ;
 assign wire13991 = ( n_n5039 ) | ( wire97 ) | ( wire13983 ) | ( wire13989 ) ;
 assign wire13992 = ( wire13981 ) | ( wire13982 ) | ( wire13990 ) ;
 assign wire13995 = ( n_n5018 ) | ( n_n5019 ) | ( n_n5015 ) | ( n_n5020 ) ;
 assign wire13996 = ( n_n5021 ) | ( wire13400 ) | ( _26122 ) ;
 assign wire13997 = ( i_9_  &  n_n509  &  n_n528  &  n_n195 ) | ( (~ i_9_)  &  n_n509  &  n_n528  &  n_n195 ) ;
 assign wire13999 = ( wire103 ) | ( wire248 ) ;
 assign wire14000 = ( n_n4998 ) | ( n_n4993 ) | ( n_n4989 ) | ( wire13997 ) ;
 assign wire14001 = ( i_9_  &  n_n526  &  n_n518  &  n_n130 ) | ( (~ i_9_)  &  n_n526  &  n_n518  &  n_n130 ) ;
 assign wire14003 = ( n_n522  &  n_n464  &  wire18 ) | ( n_n524  &  n_n464  &  wire18 ) ;
 assign wire14006 = ( n_n5081 ) | ( n_n5069 ) | ( wire14003 ) ;
 assign wire14007 = ( n_n5083 ) | ( wire160 ) | ( n_n5077 ) | ( n_n5071 ) ;
 assign wire14009 = ( i_9_  &  n_n528  &  n_n535  &  n_n130 ) | ( (~ i_9_)  &  n_n528  &  n_n535  &  n_n130 ) ;
 assign wire14010 = ( n_n5098 ) | ( n_n5084 ) | ( n_n5095 ) ;
 assign wire14011 = ( n_n5097 ) | ( n_n5089 ) | ( wire232 ) ;
 assign wire14012 = ( n_n5106 ) | ( wire14001 ) | ( wire14009 ) ;
 assign wire14015 = ( n_n1167 ) | ( wire88 ) | ( wire12917 ) | ( wire14012 ) ;
 assign wire14016 = ( wire14006 ) | ( wire14007 ) | ( wire14010 ) | ( wire14011 ) ;
 assign wire14018 = ( wire21  &  n_n195  &  n_n500 ) | ( wire24  &  n_n195  &  n_n500 ) ;
 assign wire14021 = ( n_n5013 ) | ( n_n5008 ) | ( n_n5007 ) | ( wire12931 ) ;
 assign wire14023 = ( wire13995 ) | ( wire13996 ) | ( wire13999 ) | ( wire14000 ) ;
 assign wire14025 = ( wire13991 ) | ( wire13992 ) | ( wire14015 ) | ( wire14016 ) ;
 assign wire14027 = ( n_n473  &  wire22  &  n_n130 ) | ( n_n473  &  wire11  &  n_n130 ) ;
 assign wire14028 = ( n_n5181 ) | ( n_n5184 ) | ( wire112 ) ;
 assign wire14029 = ( wire114 ) | ( wire765 ) | ( wire14027 ) ;
 assign wire14031 = ( n_n491  &  n_n524  &  wire12 ) | ( n_n491  &  n_n528  &  wire12 ) ;
 assign wire14033 = ( n_n5157 ) | ( n_n5158 ) | ( wire196 ) ;
 assign wire14034 = ( n_n5147 ) | ( wire76 ) | ( wire14031 ) ;
 assign wire14036 = ( wire25  &  n_n482  &  n_n130 ) | ( n_n482  &  wire11  &  n_n130 ) ;
 assign wire14037 = ( n_n482  &  n_n532  &  wire12 ) | ( n_n482  &  wire12  &  n_n530 ) ;
 assign wire14040 = ( n_n5175 ) | ( n_n5177 ) | ( n_n5176 ) | ( wire14037 ) ;
 assign wire14042 = ( wire14028 ) | ( wire14029 ) | ( wire14033 ) | ( wire14034 ) ;
 assign wire14043 = ( wire19  &  n_n522  &  n_n535 ) | ( wire19  &  n_n524  &  n_n535 ) ;
 assign wire14045 = ( wire449 ) | ( n_n5210 ) | ( n_n5209 ) ;
 assign wire14046 = ( n_n5212 ) | ( n_n5219 ) | ( n_n5211 ) | ( wire14043 ) ;
 assign wire14047 = ( n_n526  &  n_n464  &  wire12 ) | ( n_n464  &  n_n520  &  wire12 ) ;
 assign wire14049 = ( n_n5208 ) | ( wire761 ) | ( _26036 ) ;
 assign wire14050 = ( n_n5203 ) | ( wire220 ) | ( wire14047 ) ;
 assign wire14055 = ( n_n5193 ) | ( n_n5189 ) | ( n_n5188 ) | ( n_n5199 ) ;
 assign wire14056 = ( n_n5197 ) | ( wire451 ) | ( n_n5198 ) | ( n_n5192 ) ;
 assign wire14058 = ( wire14045 ) | ( wire14046 ) | ( wire14049 ) | ( wire14050 ) ;
 assign wire14061 = ( n_n5146 ) | ( n_n5138 ) | ( wire211 ) ;
 assign wire14062 = ( n_n5133 ) | ( n_n5144 ) | ( n_n5143 ) | ( wire12883 ) ;
 assign wire14079 = ( n_n4641 ) | ( n_n4634 ) | ( n_n4648 ) | ( n_n4618 ) ;
 assign wire14080 = ( n_n4628 ) | ( wire26 ) | ( n_n4625 ) | ( wire12545 ) ;
 assign wire14094 = ( wire22  &  n_n390  &  n_n535 ) | ( wire11  &  n_n390  &  n_n535 ) ;
 assign wire14097 = ( i_9_  &  n_n390  &  n_n535  &  n_n530 ) | ( (~ i_9_)  &  n_n390  &  n_n535  &  n_n530 ) ;
 assign wire14099 = ( n_n4576 ) | ( n_n4569 ) | ( n_n4574 ) | ( n_n4581 ) ;
 assign wire14103 = ( i_9_  &  n_n526  &  n_n464  &  n_n455 ) | ( (~ i_9_)  &  n_n526  &  n_n464  &  n_n455 ) ;
 assign wire14105 = ( n_n4568 ) | ( wire430 ) | ( wire783 ) ;
 assign wire14106 = ( wire213 ) | ( n_n4556 ) | ( wire14103 ) ;
 assign wire14111 = ( wire15  &  n_n482  &  n_n455 ) | ( n_n482  &  wire21  &  n_n455 ) ;
 assign wire14112 = ( n_n4526 ) | ( n_n4538 ) | ( n_n4535 ) | ( n_n4536 ) ;
 assign wire14128 = ( n_n4488 ) | ( n_n4483 ) | ( n_n4471 ) | ( n_n4490 ) ;
 assign wire14133 = ( n_n526  &  wire13  &  n_n535 ) | ( n_n524  &  wire13  &  n_n535 ) ;
 assign wire14134 = ( n_n526  &  n_n464  &  wire16 ) | ( n_n524  &  n_n464  &  wire16 ) ;
 assign wire14138 = ( n_n4431 ) | ( n_n4441 ) | ( wire14134 ) ;
 assign wire14139 = ( n_n4436 ) | ( n_n4439 ) | ( n_n4435 ) | ( wire421 ) ;
 assign wire14141 = ( n_n473  &  n_n536  &  wire20 ) | ( n_n473  &  n_n536  &  wire23 ) ;
 assign wire14142 = ( wire37 ) | ( n_n473  &  wire16  &  n_n520 ) ;
 assign wire14143 = ( n_n4420 ) | ( n_n4430 ) | ( wire84 ) ;
 assign wire14144 = ( n_n4451 ) | ( wire13425 ) | ( wire14141 ) ;
 assign wire14148 = ( wire14138 ) | ( wire14139 ) | ( wire14142 ) | ( wire14143 ) ;
 assign wire14149 = ( i_9_  &  n_n536  &  n_n534  &  n_n500 ) | ( (~ i_9_)  &  n_n536  &  n_n534  &  n_n500 ) ;
 assign wire14150 = ( i_9_  &  n_n522  &  n_n536  &  n_n509 ) | ( (~ i_9_)  &  n_n522  &  n_n536  &  n_n509 ) ;
 assign wire14153 = ( wire14149 ) | ( wire14150 ) ;
 assign wire14154 = ( n_n4353 ) | ( n_n4358 ) | ( wire399 ) | ( n_n4354 ) ;
 assign wire14155 = ( i_9_  &  n_n491  &  n_n536  &  n_n528 ) | ( (~ i_9_)  &  n_n491  &  n_n536  &  n_n528 ) ;
 assign wire14157 = ( i_9_  &  n_n524  &  n_n536  &  n_n500 ) | ( (~ i_9_)  &  n_n524  &  n_n536  &  n_n500 ) ;
 assign wire14158 = ( n_n4374 ) | ( n_n4373 ) | ( n_n4368 ) ;
 assign wire14159 = ( n_n4380 ) | ( n_n4372 ) | ( wire14155 ) ;
 assign wire14160 = ( n_n4362 ) | ( n_n4363 ) | ( n_n4364 ) | ( wire14157 ) ;
 assign wire14171 = ( n_n473  &  wire15  &  n_n536 ) | ( n_n473  &  wire22  &  n_n536 ) ;
 assign wire14177 = ( i_9_  &  n_n482  &  n_n536  &  n_n532 ) | ( (~ i_9_)  &  n_n482  &  n_n536  &  n_n532 ) ;
 assign wire14192 = ( n_n4345 ) | ( n_n4341 ) | ( wire67 ) | ( n_n4348 ) ;
 assign wire14198 = ( wire66 ) | ( n_n4502 ) | ( n_n4501 ) ;
 assign wire14199 = ( n_n4493 ) | ( wire13027 ) | ( _26339 ) ;
 assign wire14200 = ( i_9_  &  n_n491  &  n_n455  &  n_n530 ) | ( (~ i_9_)  &  n_n491  &  n_n455  &  n_n530 ) ;
 assign wire14202 = ( n_n4506 ) | ( wire129 ) | ( n_n4505 ) ;
 assign wire14203 = ( n_n4511 ) | ( n_n4503 ) | ( n_n4510 ) | ( wire14200 ) ;
 assign wire14205 = ( n_n4521 ) | ( n_n4517 ) | ( n_n4520 ) ;
 assign wire14208 = ( wire14198 ) | ( wire14199 ) | ( wire14202 ) | ( wire14203 ) ;
 assign wire14213 = ( wire149 ) | ( n_n5331 ) | ( wire12963 ) ;
 assign wire14214 = ( n_n3275 ) | ( wire13827 ) | ( _26519 ) ;
 assign wire14218 = ( wire13689 ) | ( wire13690 ) | ( wire13735 ) | ( wire13736 ) ;
 assign wire14219 = ( wire13741 ) | ( wire13742 ) | ( wire14218 ) ;
 assign wire14226 = ( n_n5124 ) | ( n_n5117 ) | ( wire125 ) ;
 assign wire14227 = ( n_n5135 ) | ( n_n5152 ) | ( n_n5153 ) | ( wire168 ) ;
 assign wire14232 = ( n_n5172 ) | ( n_n5207 ) | ( n_n5169 ) | ( n_n5197 ) ;
 assign wire14233 = ( wire254 ) | ( n_n5211 ) | ( n_n5176 ) | ( n_n5205 ) ;
 assign wire14238 = ( n_n5092 ) | ( n_n5110 ) | ( n_n5100 ) | ( n_n5097 ) ;
 assign wire14239 = ( n_n5087 ) | ( n_n5065 ) | ( n_n5077 ) | ( wire159 ) ;
 assign wire14240 = ( wire14238 ) | ( wire14239 ) ;
 assign wire14241 = ( wire14226 ) | ( wire14227 ) | ( wire14232 ) | ( wire14233 ) ;
 assign wire14245 = ( n_n5307 ) | ( n_n5266 ) | ( wire63 ) ;
 assign wire14246 = ( n_n5295 ) | ( n_n5290 ) | ( wire433 ) | ( n_n5283 ) ;
 assign wire14252 = ( n_n5320 ) | ( n_n5325 ) | ( wire435 ) ;
 assign wire14253 = ( n_n5232 ) | ( n_n5255 ) | ( n_n5212 ) | ( n_n5249 ) ;
 assign wire14254 = ( n_n5308 ) | ( n_n5237 ) | ( n_n5226 ) | ( n_n5218 ) ;
 assign wire14256 = ( wire14252 ) | ( wire14253 ) | ( wire14254 ) ;
 assign wire14272 = ( n_n4994 ) | ( n_n5061 ) | ( wire669 ) ;
 assign wire14273 = ( n_n5034 ) | ( n_n4996 ) | ( n_n5026 ) | ( n_n4988 ) ;
 assign wire14275 = ( n_n5057 ) | ( n_n4974 ) | ( wire14272 ) | ( wire14273 ) ;
 assign wire14277 = ( wire14245 ) | ( wire14246 ) | ( wire14256 ) | ( wire14275 ) ;
 assign wire14278 = ( n_n3558 ) | ( n_n3557 ) | ( wire14240 ) | ( wire14241 ) ;
 assign wire14280 = ( wire22  &  n_n455  &  n_n535 ) | ( wire21  &  n_n455  &  n_n535 ) ;
 assign wire14281 = ( n_n526  &  wire13  &  n_n509 ) | ( wire13  &  n_n509  &  n_n520 ) ;
 assign wire14283 = ( n_n4464 ) | ( n_n4467 ) | ( wire14280 ) ;
 assign wire14284 = ( n_n4432 ) | ( n_n4435 ) | ( n_n4493 ) | ( wire14281 ) ;
 assign wire14285 = ( n_n522  &  wire16  &  n_n535 ) | ( wire16  &  n_n532  &  n_n535 ) ;
 assign wire14290 = ( n_n4362 ) | ( n_n4317 ) | ( n_n4319 ) | ( n_n4336 ) ;
 assign wire14291 = ( n_n4355 ) | ( n_n4348 ) | ( n_n4321 ) | ( wire14285 ) ;
 assign wire14293 = ( wire21  &  n_n390  &  n_n500 ) | ( wire24  &  n_n390  &  n_n500 ) ;
 assign wire14295 = ( n_n4617 ) | ( n_n4637 ) | ( n_n4638 ) | ( n_n4626 ) ;
 assign wire14296 = ( n_n4613 ) | ( n_n4610 ) | ( n_n4632 ) | ( wire14293 ) ;
 assign wire14301 = ( n_n4514 ) | ( n_n4544 ) | ( n_n4561 ) | ( n_n4522 ) ;
 assign wire14302 = ( n_n4525 ) | ( wire65 ) | ( n_n4542 ) | ( n_n4559 ) ;
 assign wire14307 = ( n_n4602 ) | ( n_n4601 ) | ( n_n4595 ) ;
 assign wire14308 = ( n_n4568 ) | ( n_n4590 ) | ( n_n4582 ) | ( n_n4581 ) ;
 assign wire14311 = ( wire14295 ) | ( wire14296 ) | ( wire14301 ) | ( wire14302 ) ;
 assign wire14320 = ( n_n473  &  wire10  &  n_n528 ) | ( n_n473  &  wire10  &  n_n520 ) ;
 assign wire14329 = ( n_n4784 ) | ( n_n4787 ) | ( n_n4780 ) ;
 assign wire14330 = ( n_n4759 ) | ( n_n4778 ) | ( n_n4811 ) | ( n_n4793 ) ;
 assign wire14334 = ( wire16  &  n_n520  &  n_n500 ) | ( wire16  &  n_n500  &  n_n530 ) ;
 assign wire14338 = ( n_n4399 ) | ( n_n4409 ) | ( wire37 ) | ( n_n4370 ) ;
 assign wire14340 = ( wire14283 ) | ( wire14284 ) | ( wire14290 ) | ( wire14291 ) ;
 assign wire14343 = ( n_n3548 ) | ( wire14340 ) | ( _27085 ) | ( _27086 ) ;
 assign wire14344 = ( n_n518  &  wire14  &  n_n528 ) | ( n_n518  &  wire14  &  n_n520 ) ;
 assign wire14349 = ( n_n534  &  wire14  &  n_n535 ) | ( wire14  &  n_n528  &  n_n535 ) ;
 assign wire14355 = ( n_n4704 ) | ( n_n4711 ) | ( n_n4705 ) | ( n_n4706 ) ;
 assign wire14356 = ( n_n4710 ) | ( wire366 ) | ( n_n4707 ) | ( n_n4713 ) ;
 assign wire14365 = ( i_9_  &  n_n473  &  n_n532  &  n_n390 ) | ( (~ i_9_)  &  n_n473  &  n_n532  &  n_n390 ) ;
 assign wire14367 = ( i_9_  &  n_n482  &  n_n390  &  n_n520 ) | ( (~ i_9_)  &  n_n482  &  n_n390  &  n_n520 ) ;
 assign wire14373 = ( wire25  &  n_n491  &  n_n325 ) | ( n_n491  &  wire11  &  n_n325 ) ;
 assign wire14375 = ( n_n4760 ) | ( n_n4758 ) | ( n_n4764 ) | ( n_n4763 ) ;
 assign wire14376 = ( n_n4765 ) | ( n_n4766 ) | ( n_n4762 ) | ( wire14373 ) ;
 assign wire14377 = ( wire22  &  n_n509  &  n_n325 ) | ( wire21  &  n_n509  &  n_n325 ) ;
 assign wire14378 = ( n_n522  &  n_n509  &  wire14 ) | ( n_n509  &  wire14  &  n_n530 ) ;
 assign wire14380 = ( wire244 ) | ( wire14377 ) ;
 assign wire14381 = ( wire95 ) | ( n_n4742 ) | ( wire14378 ) ;
 assign wire14385 = ( n_n4755 ) | ( n_n4743 ) | ( n_n4745 ) | ( wire11834 ) ;
 assign wire14387 = ( wire14375 ) | ( wire14376 ) | ( wire14380 ) | ( wire14381 ) ;
 assign wire14396 = ( n_n482  &  n_n526  &  wire10 ) | ( n_n482  &  wire10  &  n_n530 ) ;
 assign wire14401 = ( n_n491  &  wire21  &  n_n390 ) | ( n_n491  &  wire24  &  n_n390 ) ;
 assign wire14403 = ( n_n4641 ) | ( n_n4644 ) | ( n_n4640 ) | ( n_n4639 ) ;
 assign wire14404 = ( n_n4631 ) | ( wire14401 ) | ( _26646 ) ;
 assign wire14408 = ( wire25  &  n_n473  &  n_n455 ) | ( n_n473  &  n_n455  &  wire11 ) ;
 assign wire14409 = ( n_n4539 ) | ( n_n4536 ) | ( wire201 ) ;
 assign wire14410 = ( n_n4545 ) | ( wire13091 ) | ( wire14408 ) ;
 assign wire14413 = ( n_n473  &  wire13  &  n_n520 ) | ( n_n464  &  wire13  &  n_n520 ) ;
 assign wire14414 = ( n_n4557 ) | ( wire212 ) | ( n_n4558 ) ;
 assign wire14415 = ( n_n4571 ) | ( n_n4560 ) | ( wire430 ) ;
 assign wire14416 = ( n_n4569 ) | ( n_n4556 ) | ( wire14413 ) ;
 assign wire14426 = ( i_9_  &  n_n518  &  n_n532  &  n_n390 ) | ( (~ i_9_)  &  n_n518  &  n_n532  &  n_n390 ) ;
 assign wire14428 = ( n_n4578 ) | ( n_n4575 ) | ( wire99 ) ;
 assign wire14429 = ( n_n4583 ) | ( wire239 ) | ( wire14426 ) ;
 assign wire14430 = ( i_9_  &  n_n390  &  n_n509  &  n_n528 ) | ( (~ i_9_)  &  n_n390  &  n_n509  &  n_n528 ) ;
 assign wire14432 = ( n_n4612 ) | ( n_n4611 ) | ( wire14430 ) ;
 assign wire14434 = ( n_n2037 ) | ( n_n4614 ) | ( n_n4609 ) | ( wire14432 ) ;
 assign wire14439 = ( n_n524  &  wire13  &  n_n509 ) | ( wire13  &  n_n509  &  n_n528 ) ;
 assign wire14440 = ( n_n4475 ) | ( n_n4476 ) | ( wire199 ) ;
 assign wire14441 = ( n_n4484 ) | ( wire14438 ) | ( wire14439 ) ;
 assign wire14442 = ( i_9_  &  n_n455  &  n_n528  &  n_n500 ) | ( (~ i_9_)  &  n_n455  &  n_n528  &  n_n500 ) ;
 assign wire14443 = ( n_n526  &  wire13  &  n_n500 ) | ( n_n522  &  wire13  &  n_n500 ) ;
 assign wire14444 = ( n_n4491 ) | ( n_n4492 ) | ( wire14442 ) ;
 assign wire14445 = ( n_n4488 ) | ( n_n4489 ) | ( n_n4490 ) | ( wire14443 ) ;
 assign wire14446 = ( wire25  &  n_n482  &  n_n455 ) | ( n_n482  &  n_n455  &  wire24 ) ;
 assign wire14452 = ( n_n4506 ) | ( n_n4505 ) | ( n_n4529 ) ;
 assign wire14455 = ( n_n4531 ) | ( n_n4507 ) | ( n_n4510 ) | ( n_n4501 ) ;
 assign wire14461 = ( wire25  &  n_n536  &  n_n500 ) | ( n_n536  &  wire24  &  n_n500 ) ;
 assign wire14464 = ( n_n522  &  wire16  &  n_n509 ) | ( wire16  &  n_n509  &  n_n520 ) ;
 assign wire14466 = ( n_n4359 ) | ( n_n4365 ) | ( n_n4360 ) | ( n_n4352 ) ;
 assign wire14467 = ( n_n4354 ) | ( wire14461 ) | ( wire14464 ) ;
 assign wire14468 = ( wire22  &  n_n536  &  n_n500 ) | ( n_n536  &  wire20  &  n_n500 ) ;
 assign wire14476 = ( wire16  &  n_n534  &  n_n535 ) | ( wire16  &  n_n535  &  n_n530 ) ;
 assign wire14479 = ( n_n4320 ) | ( n_n4315 ) | ( wire14476 ) ;
 assign wire14480 = ( n_n4313 ) | ( n_n4322 ) | ( n_n4323 ) | ( wire106 ) ;
 assign wire14484 = ( wire198 ) | ( wire156 ) ;
 assign wire14485 = ( n_n4344 ) | ( n_n4345 ) | ( n_n4347 ) | ( wire675 ) ;
 assign wire14486 = ( n_n4341 ) | ( n_n4351 ) | ( n_n4349 ) | ( n_n4334 ) ;
 assign wire14489 = ( n_n4340 ) | ( wire14473 ) | ( n_n2445 ) | ( wire14486 ) ;
 assign wire14490 = ( wire14479 ) | ( wire14480 ) | ( wire14484 ) | ( wire14485 ) ;
 assign wire14492 = ( n_n473  &  wire22  &  n_n536 ) | ( n_n473  &  n_n536  &  wire20 ) ;
 assign wire14493 = ( i_9_  &  n_n473  &  n_n536  &  n_n528 ) | ( (~ i_9_)  &  n_n473  &  n_n536  &  n_n528 ) ;
 assign wire14495 = ( n_n4420 ) | ( n_n4419 ) | ( wire14492 ) ;
 assign wire14496 = ( n_n4418 ) | ( wire328 ) | ( wire14493 ) ;
 assign wire14498 = ( n_n4393 ) | ( n_n4396 ) | ( n_n4395 ) | ( n_n4394 ) ;
 assign wire14499 = ( n_n4391 ) | ( n_n4397 ) | ( n_n4387 ) | ( wire12448 ) ;
 assign wire14500 = ( n_n482  &  wire22  &  n_n536 ) | ( n_n482  &  wire21  &  n_n536 ) ;
 assign wire14503 = ( i_9_  &  n_n473  &  n_n536  &  n_n532 ) | ( (~ i_9_)  &  n_n473  &  n_n536  &  n_n532 ) ;
 assign wire14505 = ( n_n4400 ) | ( n_n4407 ) | ( n_n4398 ) | ( n_n4405 ) ;
 assign wire14507 = ( n_n4402 ) | ( wire14500 ) | ( wire14503 ) | ( wire14505 ) ;
 assign wire14508 = ( wire14495 ) | ( wire14496 ) | ( wire14498 ) | ( wire14499 ) ;
 assign wire14510 = ( n_n4379 ) | ( n_n4382 ) | ( n_n4380 ) | ( n_n4377 ) ;
 assign wire14511 = ( n_n4386 ) | ( wire12447 ) | ( wire14460 ) | ( wire14510 ) ;
 assign wire14519 = ( i_9_  &  n_n464  &  n_n536  &  n_n530 ) | ( (~ i_9_)  &  n_n464  &  n_n536  &  n_n530 ) ;
 assign wire14520 = ( n_n524  &  n_n464  &  wire16 ) | ( n_n464  &  wire16  &  n_n532 ) ;
 assign wire14523 = ( n_n524  &  wire13  &  n_n535 ) | ( wire13  &  n_n534  &  n_n535 ) ;
 assign wire14524 = ( i_9_  &  n_n455  &  n_n535  &  n_n530 ) | ( (~ i_9_)  &  n_n455  &  n_n535  &  n_n530 ) ;
 assign wire14526 = ( n_n455  &  wire11  &  n_n535 ) | ( n_n455  &  wire24  &  n_n535 ) ;
 assign wire14533 = ( n_n4471 ) | ( n_n4468 ) | ( n_n4472 ) ;
 assign wire14534 = ( n_n4463 ) | ( n_n4470 ) | ( n_n4466 ) | ( n_n4469 ) ;
 assign wire14536 = ( n_n4474 ) | ( n_n4465 ) | ( wire14533 ) | ( wire14534 ) ;
 assign wire14537 = ( wire14440 ) | ( wire14441 ) | ( wire14444 ) | ( wire14445 ) ;
 assign wire14542 = ( i_9_  &  n_n65  &  n_n491  &  n_n520 ) | ( (~ i_9_)  &  n_n65  &  n_n491  &  n_n520 ) ;
 assign wire14550 = ( n_n5267 ) | ( n_n5262 ) | ( wire77 ) | ( wire92 ) ;
 assign wire14551 = ( n_n473  &  wire19  &  n_n524 ) | ( n_n473  &  wire19  &  n_n528 ) ;
 assign wire14552 = ( n_n473  &  n_n65  &  wire11 ) | ( n_n473  &  n_n65  &  wire20 ) ;
 assign wire14554 = ( n_n5305 ) | ( n_n5306 ) | ( wire14551 ) ;
 assign wire14555 = ( wire459 ) | ( n_n5315 ) | ( wire14552 ) ;
 assign wire14557 = ( n_n65  &  wire22  &  n_n464 ) | ( n_n65  &  n_n464  &  wire11 ) ;
 assign wire14558 = ( wire19  &  n_n464  &  n_n532 ) | ( wire19  &  n_n464  &  n_n530 ) ;
 assign wire14560 = ( n_n5318 ) | ( n_n5326 ) | ( wire14557 ) ;
 assign wire14561 = ( n_n5321 ) | ( n_n5328 ) | ( n_n5319 ) | ( wire14558 ) ;
 assign wire14563 = ( n_n5293 ) | ( n_n5294 ) | ( n_n5292 ) ;
 assign wire14564 = ( n_n5303 ) | ( n_n5304 ) | ( wire200 ) ;
 assign wire14566 = ( n_n5302 ) | ( n_n5299 ) | ( wire14563 ) | ( wire14564 ) ;
 assign wire14567 = ( wire14554 ) | ( wire14555 ) | ( wire14560 ) | ( wire14561 ) ;
 assign wire14570 = ( n_n65  &  wire15  &  n_n518 ) | ( n_n65  &  n_n518  &  wire21 ) ;
 assign wire14572 = ( n_n5240 ) | ( n_n5238 ) | ( n_n5244 ) | ( n_n5233 ) ;
 assign wire14573 = ( n_n5241 ) | ( n_n5234 ) | ( n_n5242 ) | ( wire14570 ) ;
 assign wire14577 = ( n_n5228 ) | ( n_n5225 ) | ( wire62 ) ;
 assign wire14578 = ( wire183 ) | ( wire434 ) ;
 assign wire14579 = ( n_n5245 ) | ( n_n5254 ) | ( n_n5217 ) | ( n_n5248 ) ;
 assign wire14580 = ( wire318 ) | ( n_n5224 ) | ( wire12874 ) | ( n_n5227 ) ;
 assign wire14582 = ( wire14579 ) | ( wire14580 ) ;
 assign wire14583 = ( wire14572 ) | ( wire14573 ) | ( wire14577 ) | ( wire14578 ) ;
 assign wire14587 = ( n_n5284 ) | ( n_n5281 ) | ( n_n5288 ) | ( n_n5291 ) ;
 assign wire14588 = ( n_n5285 ) | ( n_n5289 ) | ( n_n5282 ) | ( wire14542 ) ;
 assign wire14591 = ( n_n3664 ) | ( wire14587 ) | ( wire14588 ) | ( _27156 ) ;
 assign wire14592 = ( wire14566 ) | ( wire14567 ) | ( wire14582 ) | ( wire14583 ) ;
 assign wire14594 = ( n_n5142 ) | ( wire76 ) | ( wire679 ) ;
 assign wire14595 = ( n_n5140 ) | ( n_n5144 ) | ( n_n5143 ) | ( wire12884 ) ;
 assign wire14598 = ( wire406 ) | ( wire287 ) ;
 assign wire14599 = ( n_n5155 ) | ( n_n5163 ) | ( n_n5154 ) | ( wire195 ) ;
 assign wire14601 = ( n_n526  &  n_n509  &  wire12 ) | ( n_n509  &  wire12  &  n_n530 ) ;
 assign wire14603 = ( wire22  &  n_n509  &  n_n130 ) | ( wire11  &  n_n509  &  n_n130 ) ;
 assign wire14605 = ( n_n5115 ) | ( n_n5118 ) | ( wire14601 ) ;
 assign wire14606 = ( n_n5122 ) | ( wire286 ) | ( wire14603 ) ;
 assign wire14609 = ( n_n5111 ) | ( n_n5112 ) | ( n_n5107 ) | ( n_n5108 ) ;
 assign wire14610 = ( n_n5113 ) | ( n_n5114 ) | ( n_n5106 ) | ( wire14001 ) ;
 assign wire14621 = ( n_n473  &  wire22  &  n_n130 ) | ( n_n473  &  wire11  &  n_n130 ) ;
 assign wire14622 = ( n_n522  &  n_n464  &  wire12 ) | ( n_n464  &  n_n520  &  wire12 ) ;
 assign wire14623 = ( _514 ) | ( n_n473  &  n_n130  &  wire23 ) ;
 assign wire14631 = ( n_n482  &  wire21  &  n_n130 ) | ( n_n482  &  wire20  &  n_n130 ) ;
 assign wire14635 = ( wire114 ) | ( n_n5175 ) | ( n_n5177 ) | ( n_n5170 ) ;
 assign wire14637 = ( wire14594 ) | ( wire14595 ) | ( wire14598 ) | ( wire14599 ) ;
 assign wire14641 = ( n_n464  &  wire21  &  n_n195 ) | ( n_n464  &  n_n195  &  wire23 ) ;
 assign wire14644 = ( n_n5081 ) | ( n_n5076 ) | ( wire14641 ) ;
 assign wire14645 = ( n_n5088 ) | ( n_n5078 ) | ( n_n5083 ) | ( wire123 ) ;
 assign wire14646 = ( wire22  &  n_n535  &  n_n130 ) | ( n_n535  &  wire20  &  n_n130 ) ;
 assign wire14648 = ( wire122 ) | ( wire232 ) ;
 assign wire14649 = ( n_n5098 ) | ( n_n5103 ) | ( n_n5095 ) | ( wire14646 ) ;
 assign wire14652 = ( n_n5060 ) | ( n_n5070 ) | ( wire160 ) ;
 assign wire14656 = ( n_n473  &  n_n532  &  wire18 ) | ( n_n473  &  n_n528  &  wire18 ) ;
 assign wire14665 = ( n_n5025 ) | ( wire97 ) | ( n_n5042 ) ;
 assign wire14669 = ( i_9_  &  n_n532  &  n_n195  &  n_n500 ) | ( (~ i_9_)  &  n_n532  &  n_n195  &  n_n500 ) ;
 assign wire14671 = ( wire136 ) | ( wire299 ) ;
 assign wire14672 = ( wire103 ) | ( n_n5008 ) | ( wire14669 ) ;
 assign wire14673 = ( wire21  &  n_n509  &  n_n195 ) | ( n_n509  &  n_n195  &  wire23 ) ;
 assign wire14674 = ( n_n4998 ) | ( wire104 ) | ( wire743 ) ;
 assign wire14675 = ( n_n4989 ) | ( wire13997 ) | ( wire14673 ) ;
 assign wire14678 = ( wire21  &  n_n195  &  n_n500 ) | ( n_n195  &  wire20  &  n_n500 ) ;
 assign wire14680 = ( n_n5018 ) | ( n_n5017 ) | ( n_n5014 ) | ( n_n5020 ) ;
 assign wire14681 = ( n_n5021 ) | ( wire343 ) | ( wire14678 ) ;
 assign wire14683 = ( wire14671 ) | ( wire14672 ) | ( wire14674 ) | ( wire14675 ) ;
 assign wire14690 = ( n_n4862 ) | ( wire40 ) | ( n_n4871 ) | ( n_n4867 ) ;
 assign wire14691 = ( wire15  &  n_n518  &  n_n260 ) | ( n_n518  &  wire24  &  n_n260 ) ;
 assign wire14692 = ( n_n526  &  n_n518  &  wire17 ) | ( n_n518  &  n_n532  &  wire17 ) ;
 assign wire14695 = ( n_n4844 ) | ( wire52 ) | ( wire14692 ) ;
 assign wire14706 = ( i_9_  &  n_n524  &  n_n464  &  n_n325 ) | ( (~ i_9_)  &  n_n524  &  n_n464  &  n_n325 ) ;
 assign wire14714 = ( n_n4801 ) | ( n_n4802 ) | ( wire380 ) ;
 assign wire14715 = ( n_n4791 ) | ( n_n4803 ) | ( wire179 ) | ( n_n4799 ) ;
 assign wire14718 = ( wire313 ) | ( n_n482  &  wire22  &  n_n325 ) ;
 assign wire14719 = ( n_n4782 ) | ( n_n4779 ) | ( n_n4790 ) | ( n_n4781 ) ;
 assign wire14724 = ( i_9_  &  n_n534  &  n_n509  &  n_n260 ) | ( (~ i_9_)  &  n_n534  &  n_n509  &  n_n260 ) ;
 assign wire14726 = ( wire102 ) | ( wire14724 ) ;
 assign wire14730 = ( wire14690 ) | ( wire14695 ) | ( _26926 ) | ( _26929 ) ;
 assign wire14735 = ( wire15  &  n_n482  &  n_n260 ) | ( n_n482  &  wire11  &  n_n260 ) ;
 assign wire14738 = ( n_n4900 ) | ( n_n4903 ) | ( n_n4908 ) | ( n_n4899 ) ;
 assign wire14739 = ( n_n4905 ) | ( n_n4901 ) | ( n_n4910 ) | ( wire14735 ) ;
 assign wire14740 = ( n_n473  &  wire21  &  n_n260 ) | ( n_n473  &  wire11  &  n_n260 ) ;
 assign wire14742 = ( n_n4926 ) | ( n_n4925 ) | ( wire180 ) ;
 assign wire14743 = ( wire31 ) | ( n_n4932 ) | ( wire14740 ) ;
 assign wire14745 = ( n_n482  &  n_n526  &  wire17 ) | ( n_n482  &  wire17  &  n_n520 ) ;
 assign wire14747 = ( n_n4920 ) | ( n_n4919 ) | ( wire42 ) ;
 assign wire14748 = ( n_n4924 ) | ( n_n4947 ) | ( wire14745 ) ;
 assign wire14756 = ( i_9_  &  n_n526  &  n_n518  &  n_n195 ) | ( (~ i_9_)  &  n_n526  &  n_n518  &  n_n195 ) ;
 assign wire14759 = ( n_n522  &  n_n518  &  wire18 ) | ( n_n524  &  n_n518  &  wire18 ) ;
 assign wire14762 = ( n_n4985 ) | ( n_n4986 ) | ( wire14759 ) ;
 assign wire14766 = ( n_n526  &  wire17  &  n_n500 ) | ( n_n528  &  wire17  &  n_n500 ) ;
 assign wire14768 = ( n_n4882 ) | ( n_n4881 ) | ( wire14766 ) ;
 assign wire14770 = ( n_n4884 ) | ( n_n4877 ) | ( n_n3815 ) | ( wire14768 ) ;
 assign wire14774 = ( wire148 ) | ( wire149 ) | ( wire12963 ) ;
 assign wire14775 = ( n_n3649 ) | ( wire14387 ) | ( _27243 ) | ( _27245 ) ;
 assign wire14782 = ( wire25  &  n_n509  &  n_n130 ) | ( wire25  &  n_n535  &  n_n130 ) ;
 assign wire14784 = ( n_n5131 ) | ( n_n5087 ) | ( n_n5132 ) | ( n_n5088 ) ;
 assign wire14785 = ( n_n5095 ) | ( wire14782 ) | ( _27741 ) ;
 assign wire14790 = ( n_n5174 ) | ( n_n5184 ) | ( n_n5212 ) | ( n_n5172 ) ;
 assign wire14791 = ( n_n5234 ) | ( n_n5170 ) | ( n_n5148 ) | ( wire385 ) ;
 assign wire14795 = ( n_n5059 ) | ( wire231 ) | ( n_n5018 ) | ( n_n5045 ) ;
 assign wire14796 = ( n_n5048 ) | ( wire97 ) | ( n_n5047 ) | ( wire14795 ) ;
 assign wire14797 = ( wire14784 ) | ( wire14785 ) | ( wire14790 ) | ( wire14791 ) ;
 assign wire14808 = ( n_n518  &  wire11  &  n_n195 ) | ( n_n518  &  n_n195  &  wire23 ) ;
 assign wire14816 = ( n_n518  &  wire17  &  n_n530 ) | ( wire17  &  n_n535  &  n_n530 ) ;
 assign wire14817 = ( n_n491  &  wire22  &  n_n260 ) | ( n_n491  &  wire21  &  n_n260 ) ;
 assign wire14825 = ( n_n4925 ) | ( n_n4907 ) | ( n_n4901 ) | ( n_n4904 ) ;
 assign wire14826 = ( n_n4913 ) | ( n_n4922 ) | ( n_n4934 ) | ( wire31 ) ;
 assign wire14829 = ( n_n2451 ) | ( wire14825 ) | ( wire14826 ) ;
 assign wire14830 = ( n_n2462 ) | ( n_n2464 ) | ( wire14796 ) | ( wire14797 ) ;
 assign wire14831 = ( n_n522  &  wire10  &  n_n500 ) | ( wire10  &  n_n534  &  n_n500 ) ;
 assign wire14836 = ( n_n518  &  wire13  &  n_n520 ) | ( n_n518  &  wire13  &  n_n530 ) ;
 assign wire14843 = ( wire15  &  n_n518  &  n_n390 ) | ( n_n518  &  wire24  &  n_n390 ) ;
 assign wire14845 = ( n_n4593 ) | ( n_n4571 ) | ( n_n4527 ) ;
 assign wire14846 = ( n_n4557 ) | ( n_n4533 ) | ( wire14843 ) ;
 assign wire14859 = ( wire25  &  n_n325  &  n_n500 ) | ( wire24  &  n_n325  &  n_n500 ) ;
 assign wire14867 = ( n_n4790 ) | ( n_n4800 ) | ( n_n4826 ) ;
 assign wire14868 = ( n_n4803 ) | ( n_n4770 ) | ( n_n4772 ) | ( n_n4771 ) ;
 assign wire14873 = ( wire21  &  n_n536  &  n_n500 ) | ( n_n536  &  wire20  &  n_n500 ) ;
 assign wire14886 = ( n_n4416 ) | ( n_n4415 ) | ( n_n4448 ) | ( n_n4447 ) ;
 assign wire14887 = ( n_n4453 ) | ( n_n4420 ) | ( n_n4407 ) | ( wire234 ) ;
 assign wire14890 = ( n_n2472 ) | ( n_n2473 ) | ( wire14886 ) | ( wire14887 ) ;
 assign wire14892 = ( n_n2455 ) | ( n_n2454 ) | ( wire14890 ) ;
 assign wire14896 = ( wire25  &  n_n535  &  n_n260 ) | ( wire24  &  n_n535  &  n_n260 ) ;
 assign wire14903 = ( n_n526  &  n_n518  &  wire17 ) | ( n_n518  &  n_n532  &  wire17 ) ;
 assign wire14909 = ( n_n532  &  wire17  &  n_n500 ) | ( wire17  &  n_n500  &  n_n530 ) ;
 assign wire14910 = ( n_n4880 ) | ( wire174 ) | ( n_n4879 ) ;
 assign wire14911 = ( n_n4883 ) | ( wire14909 ) | ( _27589 ) ;
 assign wire14914 = ( n_n473  &  n_n522  &  wire14 ) | ( n_n473  &  wire14  &  n_n528 ) ;
 assign wire14915 = ( wire25  &  n_n473  &  n_n325 ) | ( n_n473  &  wire24  &  n_n325 ) ;
 assign wire14920 = ( n_n482  &  n_n524  &  wire14 ) | ( n_n482  &  wire14  &  n_n528 ) ;
 assign wire14924 = ( n_n4817 ) | ( n_n4792 ) | ( wire14920 ) ;
 assign wire14931 = ( n_n4872 ) | ( n_n4867 ) | ( _27591 ) ;
 assign wire14933 = ( n_n4866 ) | ( n_n4863 ) | ( n_n2727 ) | ( wire14931 ) ;
 assign wire14937 = ( wire22  &  n_n509  &  n_n195 ) | ( wire24  &  n_n509  &  n_n195 ) ;
 assign wire14938 = ( wire134 ) | ( wire252 ) ;
 assign wire14939 = ( n_n4996 ) | ( n_n4995 ) | ( n_n4994 ) | ( wire14937 ) ;
 assign wire14940 = ( i_9_  &  n_n195  &  n_n500  &  n_n530 ) | ( (~ i_9_)  &  n_n195  &  n_n500  &  n_n530 ) ;
 assign wire14942 = ( n_n4998 ) | ( wire393 ) | ( wire743 ) ;
 assign wire14943 = ( n_n5000 ) | ( wire136 ) | ( wire14940 ) ;
 assign wire14944 = ( n_n473  &  wire11  &  n_n260 ) | ( n_n473  &  wire24  &  n_n260 ) ;
 assign wire14946 = ( n_n473  &  n_n524  &  wire17 ) | ( n_n473  &  n_n528  &  wire17 ) ;
 assign wire14948 = ( n_n4924 ) | ( n_n4921 ) | ( wire14944 ) ;
 assign wire14949 = ( n_n4920 ) | ( n_n4919 ) | ( n_n4931 ) | ( wire14946 ) ;
 assign wire14954 = ( n_n4898 ) | ( n_n4903 ) | ( n_n4895 ) | ( n_n4908 ) ;
 assign wire14955 = ( wire96 ) | ( n_n4905 ) | ( n_n4906 ) | ( n_n4896 ) ;
 assign wire14956 = ( n_n482  &  n_n526  &  wire17 ) | ( n_n482  &  n_n522  &  wire17 ) ;
 assign wire14957 = ( i_9_  &  n_n482  &  n_n524  &  n_n260 ) | ( (~ i_9_)  &  n_n482  &  n_n524  &  n_n260 ) ;
 assign wire14960 = ( n_n4910 ) | ( wire14735 ) | ( _27623 ) ;
 assign wire14961 = ( wire14948 ) | ( wire14949 ) | ( wire14954 ) | ( wire14955 ) ;
 assign wire14962 = ( i_9_  &  n_n524  &  n_n464  &  n_n260 ) | ( (~ i_9_)  &  n_n524  &  n_n464  &  n_n260 ) ;
 assign wire14964 = ( n_n4959 ) | ( n_n4960 ) | ( wire250 ) ;
 assign wire14965 = ( n_n4964 ) | ( n_n4957 ) | ( n_n4953 ) | ( wire14752 ) ;
 assign wire14967 = ( wire25  &  n_n464  &  n_n260 ) | ( n_n464  &  n_n260  &  wire20 ) ;
 assign wire14969 = ( wire382 ) | ( n_n464  &  wire24  &  n_n260 ) ;
 assign wire14970 = ( n_n4952 ) | ( n_n4950 ) | ( wire14967 ) ;
 assign wire14971 = ( n_n4936 ) | ( n_n4935 ) | ( n_n4948 ) | ( wire14962 ) ;
 assign wire14974 = ( n_n4944 ) | ( n_n2710 ) | ( wire13867 ) | ( wire14971 ) ;
 assign wire14975 = ( wire14964 ) | ( wire14965 ) | ( wire14969 ) | ( wire14970 ) ;
 assign wire14978 = ( n_n4978 ) | ( n_n4965 ) | ( n_n4973 ) | ( wire11809 ) ;
 assign wire14979 = ( wire228 ) | ( wire771 ) | ( wire772 ) | ( wire14978 ) ;
 assign wire14980 = ( wire14938 ) | ( wire14939 ) | ( wire14942 ) | ( wire14943 ) ;
 assign wire14982 = ( wire14960 ) | ( wire14961 ) | ( wire14974 ) | ( wire14975 ) ;
 assign wire14983 = ( wire15  &  n_n325  &  n_n500 ) | ( wire22  &  n_n325  &  n_n500 ) ;
 assign wire14985 = ( wire47 ) | ( wire293 ) ;
 assign wire14986 = ( wire109 ) | ( n_n4742 ) | ( wire14983 ) ;
 assign wire14987 = ( wire21  &  n_n325  &  n_n500 ) | ( n_n325  &  wire23  &  n_n500 ) ;
 assign wire14988 = ( wire15  &  n_n491  &  n_n325 ) | ( n_n491  &  wire11  &  n_n325 ) ;
 assign wire14990 = ( n_n4764 ) | ( n_n4763 ) | ( wire14987 ) ;
 assign wire14991 = ( wire164 ) | ( n_n4761 ) | ( wire14988 ) ;
 assign wire14992 = ( n_n473  &  wire10  &  n_n532 ) | ( n_n473  &  wire10  &  n_n528 ) ;
 assign wire14993 = ( n_n473  &  n_n522  &  wire10 ) | ( n_n473  &  n_n524  &  wire10 ) ;
 assign wire14995 = ( wire157 ) | ( wire14992 ) ;
 assign wire14996 = ( n_n4671 ) | ( wire80 ) | ( wire14993 ) ;
 assign wire14999 = ( n_n4695 ) | ( n_n4696 ) | ( n_n4694 ) ;
 assign wire15000 = ( n_n4685 ) | ( n_n4686 ) | ( wire417 ) ;
 assign wire15001 = ( wire445 ) | ( wire442 ) ;
 assign wire15002 = ( n_n4698 ) | ( n_n4688 ) | ( n_n4687 ) | ( n_n4680 ) ;
 assign wire15007 = ( wire21  &  n_n325  &  n_n535 ) | ( n_n325  &  n_n535  &  wire23 ) ;
 assign wire15020 = ( n_n4779 ) | ( n_n4780 ) | ( n_n4775 ) ;
 assign wire15021 = ( n_n4774 ) | ( n_n4781 ) | ( wire315 ) ;
 assign wire15024 = ( wire14985 ) | ( wire14986 ) | ( wire14990 ) | ( wire14991 ) ;
 assign wire15035 = ( n_n491  &  wire22  &  n_n536 ) | ( n_n491  &  n_n536  &  wire20 ) ;
 assign wire15038 = ( wire425 ) | ( wire15035 ) ;
 assign wire15042 = ( n_n473  &  wire22  &  n_n536 ) | ( n_n473  &  wire21  &  n_n536 ) ;
 assign wire15043 = ( n_n473  &  wire16  &  n_n532 ) | ( n_n473  &  wire16  &  n_n528 ) ;
 assign wire15046 = ( i_9_  &  n_n482  &  n_n526  &  n_n536 ) | ( (~ i_9_)  &  n_n482  &  n_n526  &  n_n536 ) ;
 assign wire15052 = ( n_n464  &  wire16  &  n_n532 ) | ( n_n464  &  wire16  &  n_n528 ) ;
 assign wire15057 = ( n_n473  &  wire21  &  n_n455 ) | ( n_n473  &  n_n455  &  wire24 ) ;
 assign wire15058 = ( n_n473  &  n_n526  &  wire13 ) | ( n_n473  &  wire13  &  n_n532 ) ;
 assign wire15059 = ( wire25  &  n_n473  &  n_n455 ) | ( n_n473  &  wire15  &  n_n455 ) ;
 assign wire15061 = ( wire15057 ) | ( wire15058 ) ;
 assign wire15062 = ( n_n4543 ) | ( n_n4535 ) | ( n_n4536 ) | ( wire15059 ) ;
 assign wire15063 = ( n_n518  &  wire13  &  n_n532 ) | ( n_n518  &  wire13  &  n_n534 ) ;
 assign wire15071 = ( wire25  &  n_n455  &  n_n535 ) | ( wire15  &  n_n455  &  n_n535 ) ;
 assign wire15077 = ( n_n526  &  n_n491  &  wire13 ) | ( n_n491  &  n_n524  &  wire13 ) ;
 assign wire15082 = ( wire25  &  n_n455  &  n_n509 ) | ( wire15  &  n_n455  &  n_n509 ) ;
 assign wire15083 = ( n_n522  &  wire13  &  n_n509 ) | ( wire13  &  n_n532  &  n_n509 ) ;
 assign wire15084 = ( wire70 ) | ( wire15082 ) ;
 assign wire15085 = ( wire184 ) | ( wire787 ) | ( wire15083 ) ;
 assign wire15089 = ( n_n4489 ) | ( wire65 ) | ( n_n4490 ) ;
 assign wire15090 = ( n_n4497 ) | ( n_n4502 ) | ( wire347 ) ;
 assign wire15091 = ( n_n4492 ) | ( n_n4507 ) | ( n_n4505 ) | ( n_n4501 ) ;
 assign wire15097 = ( n_n482  &  n_n526  &  wire13 ) | ( n_n482  &  n_n522  &  wire13 ) ;
 assign wire15099 = ( n_n4526 ) | ( n_n4531 ) | ( n_n4529 ) | ( wire724 ) ;
 assign wire15101 = ( wire170 ) | ( n_n4534 ) | ( wire15097 ) | ( wire15099 ) ;
 assign wire15108 = ( n_n4602 ) | ( n_n4601 ) | ( wire45 ) ;
 assign wire15109 = ( wire108 ) | ( n_n4607 ) | ( n_n4600 ) | ( n_n4603 ) ;
 assign wire15111 = ( wire10  &  n_n528  &  n_n500 ) | ( wire10  &  n_n500  &  n_n530 ) ;
 assign wire15112 = ( n_n4617 ) | ( n_n4612 ) | ( n_n4611 ) | ( n_n4610 ) ;
 assign wire15113 = ( n_n4613 ) | ( wire465 ) | ( wire15111 ) ;
 assign wire15115 = ( n_n524  &  n_n518  &  wire10 ) | ( n_n518  &  wire10  &  n_n532 ) ;
 assign wire15117 = ( n_n518  &  wire21  &  n_n390 ) | ( n_n518  &  wire11  &  n_n390 ) ;
 assign wire15120 = ( n_n4597 ) | ( n_n4590 ) | ( n_n4585 ) | ( wire15117 ) ;
 assign wire15121 = ( n_n4583 ) | ( n_n4588 ) | ( wire15115 ) | ( wire15120 ) ;
 assign wire15122 = ( wire15108 ) | ( wire15109 ) | ( wire15112 ) | ( wire15113 ) ;
 assign wire15123 = ( n_n524  &  wire10  &  n_n535 ) | ( wire10  &  n_n528  &  n_n535 ) ;
 assign wire15125 = ( n_n4582 ) | ( n_n4581 ) | ( wire99 ) ;
 assign wire15126 = ( n_n4580 ) | ( wire238 ) | ( wire15123 ) ;
 assign wire15127 = ( wire25  &  n_n482  &  n_n390 ) | ( n_n482  &  wire24  &  n_n390 ) ;
 assign wire15130 = ( wire431 ) | ( wire15127 ) ;
 assign wire15131 = ( n_n4663 ) | ( n_n4652 ) | ( wire72 ) | ( n_n4657 ) ;
 assign wire15132 = ( n_n526  &  n_n491  &  wire10 ) | ( n_n491  &  wire10  &  n_n528 ) ;
 assign wire15133 = ( i_9_  &  n_n491  &  n_n532  &  n_n390 ) | ( (~ i_9_)  &  n_n491  &  n_n532  &  n_n390 ) ;
 assign wire15135 = ( wire26 ) | ( n_n4633 ) | ( n_n4630 ) ;
 assign wire15136 = ( wire310 ) | ( wire190 ) ;
 assign wire15137 = ( n_n4642 ) | ( n_n4623 ) | ( wire15133 ) ;
 assign wire15140 = ( n_n4639 ) | ( n_n2761 ) | ( wire15132 ) | ( wire15137 ) ;
 assign wire15141 = ( wire15130 ) | ( wire15131 ) | ( wire15135 ) | ( wire15136 ) ;
 assign wire15142 = ( i_9_  &  n_n526  &  n_n464  &  n_n455 ) | ( (~ i_9_)  &  n_n526  &  n_n464  &  n_n455 ) ;
 assign wire15143 = ( _462 ) | ( wire10  &  n_n535  &  n_n530 ) ;
 assign wire15144 = ( wire212 ) | ( n_n473  &  n_n455  &  wire23 ) ;
 assign wire15145 = ( n_n4570 ) | ( n_n4569 ) | ( wire15142 ) ;
 assign wire15149 = ( wire15125 ) | ( wire15126 ) | ( wire15144 ) | ( wire15145 ) ;
 assign wire15153 = ( i_9_  &  n_n518  &  n_n536  &  n_n528 ) | ( (~ i_9_)  &  n_n518  &  n_n536  &  n_n528 ) ;
 assign wire15154 = ( n_n4336 ) | ( wire198 ) | ( n_n4329 ) ;
 assign wire15155 = ( n_n4337 ) | ( wire53 ) | ( wire15153 ) ;
 assign wire15159 = ( n_n4324 ) | ( n_n4319 ) | ( wire106 ) ;
 assign wire15160 = ( n_n4326 ) | ( wire283 ) | ( n_n4321 ) | ( n_n4322 ) ;
 assign wire15162 = ( n_n4348 ) | ( n_n4353 ) | ( n_n4354 ) ;
 assign wire15163 = ( n_n4345 ) | ( wire156 ) | ( wire675 ) ;
 assign wire15165 = ( n_n4350 ) | ( n_n4340 ) | ( wire15162 ) | ( wire15163 ) ;
 assign wire15166 = ( wire15154 ) | ( wire15155 ) | ( wire15159 ) | ( wire15160 ) ;
 assign wire15174 = ( n_n5258 ) | ( n_n5255 ) | ( wire433 ) ;
 assign wire15175 = ( n_n5251 ) | ( n_n5254 ) | ( wire435 ) | ( n_n5253 ) ;
 assign wire15178 = ( n_n5244 ) | ( n_n5243 ) | ( wire320 ) ;
 assign wire15179 = ( n_n5238 ) | ( wire318 ) | ( n_n5249 ) | ( n_n5242 ) ;
 assign wire15180 = ( i_9_  &  n_n65  &  n_n526  &  n_n500 ) | ( (~ i_9_)  &  n_n65  &  n_n526  &  n_n500 ) ;
 assign wire15184 = ( n_n5270 ) | ( wire77 ) | ( _27489 ) ;
 assign wire15185 = ( wire15174 ) | ( wire15175 ) | ( wire15178 ) | ( wire15179 ) ;
 assign wire15186 = ( wire19  &  n_n526  &  n_n464 ) | ( wire19  &  n_n464  &  n_n532 ) ;
 assign wire15188 = ( n_n5321 ) | ( wire149 ) | ( n_n5319 ) ;
 assign wire15189 = ( n_n5326 ) | ( n_n5325 ) | ( n_n5327 ) | ( wire15186 ) ;
 assign wire15192 = ( wire148 ) | ( n_n3019 ) | ( n_n5312 ) | ( wire15189 ) ;
 assign wire15200 = ( i_9_  &  n_n65  &  n_n482  &  n_n532 ) | ( (~ i_9_)  &  n_n65  &  n_n482  &  n_n532 ) ;
 assign wire15203 = ( n_n5293 ) | ( n_n5294 ) | ( n_n5285 ) | ( wire15200 ) ;
 assign wire15208 = ( wire19  &  n_n522  &  n_n518 ) | ( wire19  &  n_n518  &  n_n528 ) ;
 assign wire15211 = ( n_n5228 ) | ( n_n5225 ) | ( wire15208 ) ;
 assign wire15212 = ( n_n5229 ) | ( n_n5224 ) | ( wire87 ) | ( wire182 ) ;
 assign wire15216 = ( n_n5210 ) | ( wire220 ) | ( n_n5209 ) ;
 assign wire15217 = ( wire384 ) | ( wire454 ) ;
 assign wire15218 = ( n_n5206 ) | ( n_n5222 ) | ( n_n5214 ) | ( n_n5207 ) ;
 assign wire15221 = ( wire449 ) | ( wire14043 ) | ( wire15218 ) | ( _27519 ) ;
 assign wire15222 = ( wire15211 ) | ( wire15212 ) | ( wire15216 ) | ( wire15217 ) ;
 assign wire15223 = ( n_n473  &  n_n522  &  wire18 ) | ( n_n473  &  n_n532  &  wire18 ) ;
 assign wire15224 = ( n_n473  &  wire22  &  n_n195 ) | ( n_n473  &  n_n195  &  wire20 ) ;
 assign wire15226 = ( n_n5055 ) | ( n_n5056 ) | ( wire15223 ) ;
 assign wire15227 = ( wire166 ) | ( n_n5058 ) | ( wire15224 ) ;
 assign wire15230 = ( n_n5066 ) | ( wire123 ) | ( n_n5063 ) ;
 assign wire15231 = ( n_n5070 ) | ( n_n5082 ) | ( wire159 ) ;
 assign wire15241 = ( wire15  &  n_n518  &  n_n130 ) | ( n_n518  &  wire21  &  n_n130 ) ;
 assign wire15243 = ( n_n524  &  n_n518  &  wire12 ) | ( n_n518  &  n_n528  &  wire12 ) ;
 assign wire15247 = ( n_n5091 ) | ( n_n5108 ) | ( wire13305 ) | ( wire88 ) ;
 assign wire15252 = ( wire15  &  n_n482  &  n_n195 ) | ( n_n482  &  wire21  &  n_n195 ) ;
 assign wire15254 = ( n_n5036 ) | ( n_n5049 ) | ( wire253 ) ;
 assign wire15255 = ( n_n5039 ) | ( wire356 ) | ( wire15252 ) ;
 assign wire15257 = ( n_n5027 ) | ( n_n5028 ) | ( wire265 ) ;
 assign wire15258 = ( n_n5026 ) | ( wire50 ) | ( n_n5023 ) | ( n_n5029 ) ;
 assign wire15261 = ( n_n5022 ) | ( n_n5011 ) | ( n_n5013 ) | ( wire12931 ) ;
 assign wire15263 = ( wire15254 ) | ( wire15255 ) | ( wire15257 ) | ( wire15258 ) ;
 assign wire15266 = ( n_n473  &  wire15  &  n_n130 ) | ( n_n473  &  wire22  &  n_n130 ) ;
 assign wire15269 = ( n_n5191 ) | ( n_n5192 ) | ( wire15266 ) ;
 assign wire15270 = ( wire112 ) | ( n_n5193 ) | ( n_n5182 ) | ( n_n5190 ) ;
 assign wire15273 = ( n_n5201 ) | ( wire437 ) | ( wire761 ) ;
 assign wire15274 = ( n_n5175 ) | ( n_n5177 ) | ( wire451 ) ;
 assign wire15275 = ( n_n5173 ) | ( n_n5203 ) | ( n_n5197 ) | ( n_n5176 ) ;
 assign wire15278 = ( wire114 ) | ( n_n2670 ) | ( wire765 ) | ( wire15275 ) ;
 assign wire15279 = ( wire15269 ) | ( wire15270 ) | ( wire15273 ) | ( wire15274 ) ;
 assign wire15280 = ( n_n482  &  n_n532  &  wire12 ) | ( n_n482  &  wire12  &  n_n530 ) ;
 assign wire15284 = ( n_n5163 ) | ( n_n5157 ) | ( wire195 ) | ( n_n5160 ) ;
 assign wire15285 = ( wire25  &  n_n491  &  n_n130 ) | ( n_n491  &  wire21  &  n_n130 ) ;
 assign wire15288 = ( wire196 ) | ( n_n5149 ) | ( wire15285 ) ;
 assign wire15289 = ( wire22  &  n_n130  &  n_n500 ) | ( wire11  &  n_n130  &  n_n500 ) ;
 assign wire15290 = ( i_9_  &  n_n524  &  n_n130  &  n_n500 ) | ( (~ i_9_)  &  n_n524  &  n_n130  &  n_n500 ) ;
 assign wire15292 = ( n_n5130 ) | ( n_n5133 ) | ( n_n5134 ) | ( wire15290 ) ;
 assign wire15294 = ( wire15284 ) | ( wire15288 ) | ( _27515 ) ;
 assign wire15296 = ( wire15221 ) | ( wire15222 ) | ( wire15278 ) | ( wire15279 ) ;
 assign wire15304 = ( n_n491  &  n_n536  &  wire23 ) | ( n_n536  &  n_n509  &  wire23 ) ;
 assign wire15310 = ( wire21  &  n_n455  &  n_n535 ) | ( n_n455  &  n_n535  &  wire20 ) ;
 assign wire15312 = ( n_n518  &  wire13  &  n_n532 ) | ( n_n518  &  wire13  &  n_n534 ) ;
 assign wire15315 = ( n_n4487 ) | ( n_n4478 ) | ( wire15312 ) ;
 assign wire15316 = ( n_n4488 ) | ( n_n4476 ) | ( n_n4457 ) | ( wire15310 ) ;
 assign wire15326 = ( wire10  &  n_n534  &  n_n509 ) | ( wire10  &  n_n509  &  n_n528 ) ;
 assign wire15340 = ( n_n4514 ) | ( n_n4511 ) | ( n_n4525 ) | ( n_n4528 ) ;
 assign wire15341 = ( n_n4552 ) | ( wire416 ) | ( n_n4527 ) | ( n_n4534 ) ;
 assign wire15375 = ( n_n5169 ) | ( wire33 ) | ( n_n5235 ) | ( n_n5217 ) ;
 assign wire15376 = ( n_n65  &  wire15  &  n_n464 ) | ( n_n65  &  wire22  &  n_n464 ) ;
 assign wire15382 = ( n_n5302 ) | ( n_n5273 ) | ( n_n5327 ) | ( n_n5254 ) ;
 assign wire15383 = ( n_n5278 ) | ( n_n5319 ) | ( wire200 ) | ( n_n5282 ) ;
 assign wire15385 = ( wire386 ) | ( wire15376 ) | ( wire15382 ) | ( wire15383 ) ;
 assign wire15396 = ( n_n4921 ) | ( n_n4938 ) | ( n_n4936 ) | ( n_n4917 ) ;
 assign wire15397 = ( n_n4931 ) | ( n_n4948 ) | ( n_n4957 ) | ( wire141 ) ;
 assign wire15416 = ( n_n4711 ) | ( n_n4732 ) | ( _28071 ) ;
 assign wire15421 = ( wire15  &  n_n455  &  n_n509 ) | ( n_n455  &  wire24  &  n_n509 ) ;
 assign wire15428 = ( i_9_  &  n_n455  &  n_n528  &  n_n500 ) | ( (~ i_9_)  &  n_n455  &  n_n528  &  n_n500 ) ;
 assign wire15431 = ( n_n4491 ) | ( n_n4492 ) | ( wire15428 ) ;
 assign wire15432 = ( n_n4497 ) | ( wire65 ) | ( n_n4500 ) | ( n_n4496 ) ;
 assign wire15434 = ( n_n4506 ) | ( n_n4505 ) | ( n_n4490 ) ;
 assign wire15435 = ( n_n4504 ) | ( n_n4502 ) | ( n_n4507 ) | ( n_n4501 ) ;
 assign wire15448 = ( n_n473  &  n_n524  &  wire13 ) | ( n_n473  &  wire13  &  n_n532 ) ;
 assign wire15456 = ( n_n522  &  wire13  &  n_n535 ) | ( n_n524  &  wire13  &  n_n535 ) ;
 assign wire15459 = ( n_n4463 ) | ( n_n4455 ) | ( wire15456 ) ;
 assign wire15460 = ( n_n4454 ) | ( n_n4465 ) | ( n_n4462 ) | ( wire291 ) ;
 assign wire15468 = ( n_n4666 ) | ( n_n4648 ) | ( wire139 ) ;
 assign wire15469 = ( n_n4644 ) | ( n_n4658 ) | ( n_n4642 ) | ( wire13454 ) ;
 assign wire15472 = ( wire13888 ) | ( wire15468 ) | ( _28116 ) ;
 assign wire15474 = ( n_n4568 ) | ( wire783 ) | ( wire276 ) ;
 assign wire15475 = ( n_n4574 ) | ( n_n4573 ) | ( wire455 ) | ( wire671 ) ;
 assign wire15478 = ( n_n4582 ) | ( n_n4584 ) | ( _28106 ) ;
 assign wire15479 = ( n_n4587 ) | ( wire365 ) | ( n_n4580 ) | ( n_n4585 ) ;
 assign wire15481 = ( wire10  &  n_n532  &  n_n500 ) | ( wire10  &  n_n500  &  n_n530 ) ;
 assign wire15482 = ( n_n4617 ) | ( n_n4613 ) | ( n_n4607 ) | ( n_n4610 ) ;
 assign wire15483 = ( n_n4616 ) | ( wire465 ) | ( wire15481 ) ;
 assign wire15485 = ( n_n524  &  n_n518  &  wire10 ) | ( n_n518  &  wire10  &  n_n528 ) ;
 assign wire15488 = ( n_n4593 ) | ( n_n4601 ) | ( wire15485 ) ;
 assign wire15489 = ( wire108 ) | ( n_n4603 ) | ( n_n4595 ) | ( n_n4592 ) ;
 assign wire15490 = ( i_9_  &  n_n522  &  n_n390  &  n_n500 ) | ( (~ i_9_)  &  n_n522  &  n_n390  &  n_n500 ) ;
 assign wire15493 = ( n_n4639 ) | ( n_n4621 ) | ( n_n4632 ) | ( wire12547 ) ;
 assign wire15495 = ( wire15482 ) | ( wire15483 ) | ( wire15488 ) | ( wire15489 ) ;
 assign wire15498 = ( n_n4557 ) | ( n_n4558 ) | ( n_n4559 ) ;
 assign wire15499 = ( n_n4560 ) | ( n_n4553 ) | ( wire430 ) ;
 assign wire15509 = ( wire16  &  n_n532  &  n_n500 ) | ( wire16  &  n_n528  &  n_n500 ) ;
 assign wire15525 = ( n_n4331 ) | ( n_n4336 ) | ( n_n4334 ) | ( wire677 ) ;
 assign wire15526 = ( n_n4337 ) | ( n_n4332 ) | ( n_n4329 ) | ( wire53 ) ;
 assign wire15529 = ( n_n526  &  n_n464  &  wire16 ) | ( n_n524  &  n_n464  &  wire16 ) ;
 assign wire15532 = ( n_n4430 ) | ( n_n4429 ) | ( wire15529 ) ;
 assign wire15533 = ( n_n4433 ) | ( n_n4438 ) | ( n_n4425 ) | ( wire84 ) ;
 assign wire15534 = ( n_n473  &  n_n526  &  wire16 ) | ( n_n473  &  n_n522  &  wire16 ) ;
 assign wire15536 = ( wire215 ) | ( wire79 ) ;
 assign wire15537 = ( n_n4414 ) | ( n_n4411 ) | ( n_n4412 ) | ( wire15534 ) ;
 assign wire15538 = ( n_n482  &  wire21  &  n_n536 ) | ( n_n482  &  n_n536  &  wire23 ) ;
 assign wire15539 = ( n_n482  &  n_n522  &  wire16 ) | ( n_n482  &  wire16  &  n_n520 ) ;
 assign wire15542 = ( n_n4408 ) | ( n_n4401 ) | ( n_n4402 ) | ( wire15539 ) ;
 assign wire15546 = ( n_n4378 ) | ( n_n4381 ) | ( wire423 ) | ( wire12449 ) ;
 assign wire15551 = ( n_n526  &  n_n464  &  wire12 ) | ( n_n464  &  n_n520  &  wire12 ) ;
 assign wire15554 = ( n_n5207 ) | ( n_n5208 ) | ( wire15551 ) ;
 assign wire15555 = ( n_n5199 ) | ( wire220 ) | ( n_n5209 ) | ( wire636 ) ;
 assign wire15557 = ( wire19  &  n_n522  &  n_n535 ) | ( wire19  &  n_n532  &  n_n535 ) ;
 assign wire15559 = ( n_n5191 ) | ( wire454 ) | ( n_n5192 ) ;
 assign wire15560 = ( wire183 ) | ( wire453 ) ;
 assign wire15562 = ( wire112 ) | ( n_n5215 ) | ( n_n5198 ) | ( wire14615 ) ;
 assign wire15565 = ( wire15554 ) | ( wire15555 ) | ( wire15559 ) | ( wire15560 ) ;
 assign wire15569 = ( n_n5223 ) | ( n_n5229 ) | ( wire182 ) ;
 assign wire15570 = ( n_n5228 ) | ( n_n5225 ) | ( n_n5224 ) | ( wire385 ) ;
 assign wire15573 = ( n_n5239 ) | ( n_n5240 ) | ( n_n5244 ) | ( n_n5243 ) ;
 assign wire15574 = ( wire62 ) | ( wire446 ) ;
 assign wire15575 = ( n_n5241 ) | ( n_n5262 ) | ( n_n5234 ) | ( n_n5246 ) ;
 assign wire15576 = ( wire435 ) | ( wire433 ) | ( _28280 ) ;
 assign wire15579 = ( wire15569 ) | ( wire15570 ) | ( wire15573 ) | ( wire15574 ) ;
 assign wire15582 = ( n_n482  &  wire11  &  n_n130 ) | ( n_n482  &  wire24  &  n_n130 ) ;
 assign wire15583 = ( wire15582 ) | ( n_n482  &  n_n522  &  wire12 ) ;
 assign wire15586 = ( n_n5142 ) | ( wire196 ) | ( wire679 ) ;
 assign wire15587 = ( n_n5146 ) | ( wire76 ) | ( n_n5139 ) | ( n_n5151 ) ;
 assign wire15589 = ( i_9_  &  n_n473  &  n_n534  &  n_n130 ) | ( (~ i_9_)  &  n_n473  &  n_n534  &  n_n130 ) ;
 assign wire15591 = ( n_n5181 ) | ( n_n5182 ) | ( wire732 ) | ( wire15589 ) ;
 assign wire15593 = ( wire466 ) | ( wire15583 ) | ( wire15586 ) | ( wire15587 ) ;
 assign wire15595 = ( wire15565 ) | ( wire15579 ) | ( _28289 ) ;
 assign wire15596 = ( wire15  &  n_n482  &  n_n195 ) | ( n_n482  &  n_n195  &  wire20 ) ;
 assign wire15597 = ( n_n5043 ) | ( n_n5044 ) | ( wire15596 ) ;
 assign wire15598 = ( n_n473  &  n_n532  &  wire18 ) | ( n_n473  &  n_n528  &  wire18 ) ;
 assign wire15612 = ( wire25  &  n_n535  &  n_n130 ) | ( wire15  &  n_n535  &  n_n130 ) ;
 assign wire15614 = ( i_9_  &  n_n524  &  n_n464  &  n_n195 ) | ( (~ i_9_)  &  n_n524  &  n_n464  &  n_n195 ) ;
 assign wire15620 = ( n_n518  &  wire11  &  n_n130 ) | ( n_n518  &  wire20  &  n_n130 ) ;
 assign wire15621 = ( n_n526  &  n_n518  &  wire12 ) | ( n_n518  &  n_n528  &  wire12 ) ;
 assign wire15623 = ( n_n5112 ) | ( n_n5110 ) | ( wire15620 ) ;
 assign wire15624 = ( n_n5107 ) | ( n_n5106 ) | ( n_n5108 ) | ( wire15621 ) ;
 assign wire15626 = ( wire11  &  n_n509  &  n_n130 ) | ( wire24  &  n_n509  &  n_n130 ) ;
 assign wire15627 = ( n_n524  &  wire12  &  n_n500 ) | ( n_n528  &  wire12  &  n_n500 ) ;
 assign wire15628 = ( wire335 ) | ( n_n5121 ) | ( n_n5122 ) ;
 assign wire15629 = ( n_n5136 ) | ( n_n5124 ) | ( wire286 ) ;
 assign wire15639 = ( n_n5036 ) | ( wire231 ) | ( n_n5031 ) | ( n_n5029 ) ;
 assign wire15647 = ( _226 ) | ( wire19  &  n_n464  &  n_n532 ) ;
 assign wire15648 = ( n_n5318 ) | ( n_n5320 ) | ( n_n5315 ) ;
 assign wire15649 = ( _28312 ) | ( _28313 ) ;
 assign wire15651 = ( wire19  &  n_n522  &  n_n491 ) | ( wire19  &  n_n491  &  n_n530 ) ;
 assign wire15658 = ( n_n5270 ) | ( n_n5269 ) | ( wire205 ) ;
 assign wire15659 = ( n_n5268 ) | ( n_n5271 ) | ( wire334 ) | ( wire92 ) ;
 assign wire15660 = ( n_n473  &  wire19  &  n_n524 ) | ( n_n473  &  wire19  &  n_n528 ) ;
 assign wire15666 = ( n_n5291 ) | ( n_n5292 ) | ( n_n5289 ) ;
 assign wire15667 = ( n_n5293 ) | ( n_n5294 ) | ( n_n5288 ) | ( n_n5286 ) ;
 assign wire15671 = ( n_n5328 ) | ( n_n5335 ) | ( wire149 ) | ( n_n5331 ) ;
 assign wire15672 = ( wire15647 ) | ( wire15648 ) | ( wire15649 ) | ( wire15671 ) ;
 assign wire15675 = ( n_n2939 ) | ( wire15658 ) | ( wire15659 ) | ( wire15672 ) ;
 assign wire15677 = ( wire15595 ) | ( wire15675 ) | ( _28320 ) ;
 assign wire15678 = ( n_n526  &  n_n509  &  wire17 ) | ( n_n509  &  wire17  &  n_n530 ) ;
 assign wire15680 = ( n_n4862 ) | ( n_n4869 ) | ( n_n4870 ) | ( n_n4861 ) ;
 assign wire15681 = ( wire245 ) | ( n_n4868 ) | ( wire15678 ) ;
 assign wire15683 = ( wire96 ) | ( wire49 ) ;
 assign wire15684 = ( wire12179 ) | ( n_n4896 ) | ( _27917 ) ;
 assign wire15685 = ( _298 ) | ( wire17  &  n_n535  &  n_n530 ) ;
 assign wire15686 = ( n_n4830 ) | ( n_n4827 ) | ( n_n4824 ) | ( wire693 ) ;
 assign wire15688 = ( i_9_  &  n_n534  &  n_n509  &  n_n260 ) | ( (~ i_9_)  &  n_n534  &  n_n509  &  n_n260 ) ;
 assign wire15689 = ( wire22  &  n_n518  &  n_n260 ) | ( n_n518  &  n_n260  &  wire20 ) ;
 assign wire15693 = ( n_n4855 ) | ( n_n4842 ) | ( wire15689 ) ;
 assign wire15695 = ( wire176 ) | ( wire52 ) | ( wire375 ) | ( wire15688 ) ;
 assign wire15696 = ( n_n3820 ) | ( n_n4836 ) | ( wire11769 ) | ( wire15693 ) ;
 assign wire15697 = ( n_n3461 ) | ( wire15685 ) | ( wire15686 ) | ( wire15695 ) ;
 assign wire15698 = ( n_n473  &  n_n526  &  wire17 ) | ( n_n473  &  n_n532  &  wire17 ) ;
 assign wire15700 = ( n_n4925 ) | ( n_n4919 ) | ( _27868 ) ;
 assign wire15701 = ( n_n4930 ) | ( wire382 ) | ( wire15698 ) ;
 assign wire15702 = ( n_n491  &  n_n532  &  wire18 ) | ( n_n491  &  n_n528  &  wire18 ) ;
 assign wire15704 = ( wire296 ) | ( n_n5019 ) | ( n_n5020 ) ;
 assign wire15705 = ( n_n5017 ) | ( wire135 ) | ( wire15702 ) ;
 assign wire15707 = ( n_n534  &  wire18  &  n_n500 ) | ( wire18  &  n_n500  &  n_n530 ) ;
 assign wire15709 = ( n_n4998 ) | ( wire136 ) | ( wire743 ) ;
 assign wire15710 = ( wire394 ) | ( wire104 ) ;
 assign wire15712 = ( n_n4994 ) | ( n_n5003 ) | ( wire12255 ) | ( wire12256 ) ;
 assign wire15715 = ( wire15704 ) | ( wire15705 ) | ( wire15709 ) | ( wire15710 ) ;
 assign wire15718 = ( n_n4988 ) | ( n_n4987 ) | ( wire251 ) ;
 assign wire15719 = ( n_n4991 ) | ( n_n4981 ) | ( n_n4985 ) | ( wire57 ) ;
 assign wire15721 = ( n_n524  &  n_n535  &  wire18 ) | ( n_n535  &  n_n520  &  wire18 ) ;
 assign wire15723 = ( wire25  &  n_n535  &  n_n195 ) | ( wire24  &  n_n535  &  n_n195 ) ;
 assign wire15724 = ( wire341 ) | ( wire317 ) ;
 assign wire15725 = ( n_n4958 ) | ( n_n4947 ) | ( wire15721 ) ;
 assign wire15729 = ( wire15718 ) | ( wire15719 ) | ( wire15724 ) | ( wire15725 ) ;
 assign wire15733 = ( n_n4942 ) | ( wire59 ) | ( n_n4940 ) | ( n_n4939 ) ;
 assign wire15734 = ( n_n4946 ) | ( n_n4937 ) | ( wire180 ) | ( n_n4944 ) ;
 assign wire15738 = ( n_n4913 ) | ( n_n4916 ) | ( wire305 ) ;
 assign wire15739 = ( n_n4905 ) | ( n_n4918 ) | ( n_n4914 ) | ( wire340 ) ;
 assign wire15741 = ( wire15700 ) | ( wire15701 ) | ( wire15733 ) | ( wire15734 ) ;
 assign wire15747 = ( n_n4724 ) | ( n_n4727 ) | ( n_n4739 ) | ( wire95 ) ;
 assign wire15748 = ( wire15  &  n_n518  &  n_n325 ) | ( n_n518  &  wire11  &  n_n325 ) ;
 assign wire15754 = ( wire25  &  n_n482  &  n_n325 ) | ( n_n482  &  wire22  &  n_n325 ) ;
 assign wire15756 = ( n_n4784 ) | ( n_n4779 ) | ( n_n4786 ) | ( n_n4783 ) ;
 assign wire15757 = ( n_n4782 ) | ( n_n4781 ) | ( n_n4775 ) | ( wire15754 ) ;
 assign wire15758 = ( i_9_  &  n_n325  &  n_n520  &  n_n500 ) | ( (~ i_9_)  &  n_n325  &  n_n520  &  n_n500 ) ;
 assign wire15760 = ( n_n4756 ) | ( n_n4753 ) | ( n_n4761 ) | ( n_n4762 ) ;
 assign wire15761 = ( wire109 ) | ( n_n4752 ) | ( wire15758 ) ;
 assign wire15763 = ( n_n526  &  n_n491  &  wire14 ) | ( n_n491  &  wire14  &  n_n528 ) ;
 assign wire15773 = ( i_9_  &  n_n464  &  n_n390  &  n_n520 ) | ( (~ i_9_)  &  n_n464  &  n_n390  &  n_n520 ) ;
 assign wire15776 = ( n_n4707 ) | ( n_n4696 ) | ( wire13897 ) | ( wire13755 ) ;
 assign wire15781 = ( n_n4748 ) | ( n_n4747 ) | ( n_n4742 ) ;
 assign wire15784 = ( wire374 ) | ( wire47 ) | ( wire15781 ) | ( _27859 ) ;
 assign wire15790 = ( wire158 ) | ( wire380 ) ;
 assign wire15791 = ( n_n4787 ) | ( wire292 ) | ( n_n4795 ) | ( n_n4799 ) ;
 assign wire15792 = ( n_n473  &  n_n526  &  wire14 ) | ( n_n526  &  n_n464  &  wire14 ) ;
 assign wire15794 = ( n_n4803 ) | ( n_n4804 ) | ( n_n4807 ) | ( n_n4808 ) ;
 assign wire15795 = ( n_n4801 ) | ( n_n4802 ) | ( wire15792 ) ;
 assign wire15798 = ( n_n4806 ) | ( n_n4805 ) | ( n_n4197 ) | ( wire390 ) ;
 assign wire15799 = ( wire15790 ) | ( wire15791 ) | ( wire15794 ) | ( wire15795 ) ;
 assign wire15800 = ( n_n524  &  wire17  &  n_n500 ) | ( n_n528  &  wire17  &  n_n500 ) ;
 assign wire15802 = ( wire174 ) | ( wire15800 ) ;
 assign wire15805 = ( wire15680 ) | ( wire15681 ) | ( wire15683 ) | ( wire15684 ) ;
 assign wire15807 = ( wire15696 ) | ( wire15697 ) | ( wire15798 ) | ( wire15799 ) ;
 assign wire15811 = ( n_n2845 ) | ( n_n2846 ) | ( wire15315 ) | ( wire15316 ) ;
 assign wire15813 = ( n_n2827 ) | ( n_n2826 ) | ( wire15811 ) ;
 assign wire15819 = ( n_n491  &  wire22  &  n_n455 ) | ( n_n491  &  wire21  &  n_n455 ) ;
 assign wire15834 = ( wire13  &  n_n532  &  n_n509 ) | ( wire13  &  n_n509  &  n_n520 ) ;
 assign wire15836 = ( n_n4478 ) | ( n_n4502 ) | ( n_n4509 ) | ( n_n4471 ) ;
 assign wire15837 = ( n_n4473 ) | ( n_n4497 ) | ( wire617 ) | ( wire15834 ) ;
 assign wire15841 = ( n_n482  &  wire19  &  n_n520 ) | ( wire19  &  n_n509  &  n_n520 ) ;
 assign wire15842 = ( n_n65  &  n_n482  &  wire11 ) | ( n_n65  &  n_n482  &  wire24 ) ;
 assign wire15843 = ( _198 ) | ( n_n65  &  n_n509  &  wire20 ) ;
 assign wire15844 = ( n_n5238 ) | ( n_n5245 ) | ( n_n5280 ) ;
 assign wire15845 = ( wire15841 ) | ( wire15842 ) ;
 assign wire15848 = ( n_n522  &  n_n509  &  wire17 ) | ( n_n509  &  wire17  &  n_n530 ) ;
 assign wire15864 = ( n_n4993 ) | ( n_n4994 ) | ( wire248 ) ;
 assign wire15865 = ( wire136 ) | ( n_n5009 ) | ( n_n4978 ) | ( n_n5001 ) ;
 assign wire15873 = ( i_9_  &  n_n473  &  n_n532  &  n_n130 ) | ( (~ i_9_)  &  n_n473  &  n_n532  &  n_n130 ) ;
 assign wire15876 = ( wire15  &  n_n491  &  n_n130 ) | ( wire15  &  n_n130  &  n_n500 ) ;
 assign wire15880 = ( n_n473  &  n_n532  &  wire18 ) | ( n_n482  &  n_n532  &  wire18 ) ;
 assign wire15885 = ( n_n5059 ) | ( n_n5018 ) | ( n_n5022 ) | ( n_n5046 ) ;
 assign wire15886 = ( n_n5033 ) | ( n_n5063 ) | ( n_n5052 ) | ( wire15880 ) ;
 assign wire15887 = ( wire15885 ) | ( wire15886 ) ;
 assign wire15892 = ( i_9_  &  n_n65  &  n_n524  &  n_n535 ) | ( (~ i_9_)  &  n_n65  &  n_n524  &  n_n535 ) ;
 assign wire15894 = ( n_n5214 ) | ( n_n5207 ) | ( n_n5229 ) | ( n_n5221 ) ;
 assign wire15895 = ( n_n5200 ) | ( n_n5222 ) | ( n_n5203 ) | ( wire15892 ) ;
 assign wire15897 = ( n_n65  &  n_n464  &  wire21 ) | ( n_n65  &  n_n464  &  wire20 ) ;
 assign wire15898 = ( n_n5325 ) | ( n_n5303 ) | ( wire15897 ) ;
 assign wire15899 = ( wire15843 ) | ( wire15844 ) | ( wire15845 ) | ( wire15898 ) ;
 assign wire15901 = ( wire15864 ) | ( wire15865 ) | ( wire15894 ) | ( wire15895 ) ;
 assign wire15902 = ( n_n1722 ) | ( n_n1721 ) | ( wire15899 ) ;
 assign wire15903 = ( n_n1718 ) | ( n_n1717 ) | ( wire15887 ) | ( wire15901 ) ;
 assign wire15922 = ( n_n518  &  n_n325  &  wire23 ) | ( n_n325  &  n_n535  &  wire23 ) ;
 assign wire15927 = ( wire15  &  n_n482  &  n_n325 ) | ( n_n482  &  wire21  &  n_n325 ) ;
 assign wire15937 = ( n_n4337 ) | ( n_n4314 ) | ( n_n4345 ) | ( wire675 ) ;
 assign wire15938 = ( n_n4371 ) | ( n_n4343 ) | ( n_n4320 ) | ( wire345 ) ;
 assign wire15941 = ( n_n1730 ) | ( n_n1729 ) | ( wire15937 ) | ( wire15938 ) ;
 assign wire15943 = ( n_n1712 ) | ( n_n1711 ) | ( wire15941 ) ;
 assign wire15947 = ( i_9_  &  n_n522  &  n_n535  &  n_n130 ) | ( (~ i_9_)  &  n_n522  &  n_n535  &  n_n130 ) ;
 assign wire15952 = ( n_n473  &  n_n522  &  wire18 ) | ( n_n473  &  n_n528  &  wire18 ) ;
 assign wire15954 = ( n_n5057 ) | ( n_n5058 ) | ( n_n5065 ) ;
 assign wire15964 = ( n_n518  &  wire21  &  n_n130 ) | ( n_n518  &  wire20  &  n_n130 ) ;
 assign wire15970 = ( n_n522  &  wire12  &  n_n500 ) | ( wire12  &  n_n500  &  n_n530 ) ;
 assign wire15972 = ( n_n5136 ) | ( n_n5135 ) | ( n_n5134 ) | ( wire15970 ) ;
 assign wire15975 = ( n_n482  &  n_n524  &  wire18 ) | ( n_n482  &  n_n528  &  wire18 ) ;
 assign wire15980 = ( n_n491  &  n_n524  &  wire18 ) | ( n_n491  &  n_n534  &  wire18 ) ;
 assign wire15982 = ( wire296 ) | ( wire265 ) ;
 assign wire15983 = ( wire135 ) | ( n_n5020 ) | ( wire15980 ) ;
 assign wire15985 = ( i_9_  &  n_n482  &  n_n195  &  n_n530 ) | ( (~ i_9_)  &  n_n482  &  n_n195  &  n_n530 ) ;
 assign wire15987 = ( n_n5035 ) | ( n_n5032 ) | ( n_n5027 ) | ( n_n5028 ) ;
 assign wire15989 = ( wire50 ) | ( n_n5029 ) | ( wire15985 ) | ( wire15987 ) ;
 assign wire15991 = ( n_n1842 ) | ( wire15982 ) | ( wire15983 ) | ( wire15989 ) ;
 assign wire15993 = ( n_n526  &  wire13  &  n_n500 ) | ( wire13  &  n_n500  &  n_n530 ) ;
 assign wire15999 = ( i_9_  &  n_n522  &  n_n464  &  n_n536 ) | ( (~ i_9_)  &  n_n522  &  n_n464  &  n_n536 ) ;
 assign wire16001 = ( n_n4434 ) | ( wire234 ) | ( n_n4431 ) ;
 assign wire16002 = ( wire233 ) | ( n_n4447 ) | ( wire15999 ) ;
 assign wire16003 = ( n_n4470 ) | ( n_n4472 ) | ( n_n4469 ) ;
 assign wire16004 = ( wire11505 ) | ( wire14133 ) | ( _28677 ) ;
 assign wire16007 = ( n_n4462 ) | ( wire12471 ) | ( n_n2058 ) | ( wire16004 ) ;
 assign wire16008 = ( n_n3889 ) | ( wire16001 ) | ( wire16002 ) | ( wire16003 ) ;
 assign wire16009 = ( n_n482  &  wire21  &  n_n455 ) | ( n_n482  &  n_n455  &  wire20 ) ;
 assign wire16011 = ( n_n4535 ) | ( n_n4536 ) | ( wire16009 ) ;
 assign wire16012 = ( n_n4532 ) | ( n_n4537 ) | ( n_n4529 ) | ( wire11532 ) ;
 assign wire16014 = ( wire170 ) | ( n_n491  &  n_n455  &  wire20 ) ;
 assign wire16015 = ( n_n4520 ) | ( wire361 ) | ( wire789 ) ;
 assign wire16016 = ( n_n4521 ) | ( n_n4526 ) | ( n_n4542 ) | ( wire201 ) ;
 assign wire16018 = ( wire202 ) | ( wire16016 ) ;
 assign wire16019 = ( wire16011 ) | ( wire16012 ) | ( wire16014 ) | ( wire16015 ) ;
 assign wire16020 = ( n_n526  &  n_n491  &  wire13 ) | ( n_n491  &  n_n524  &  wire13 ) ;
 assign wire16022 = ( n_n4506 ) | ( n_n4505 ) | ( wire606 ) ;
 assign wire16023 = ( n_n4504 ) | ( n_n4503 ) | ( wire16020 ) ;
 assign wire16031 = ( n_n4584 ) | ( n_n4580 ) | ( n_n4585 ) | ( wire12520 ) ;
 assign wire16032 = ( wire11  &  n_n390  &  n_n535 ) | ( wire24  &  n_n390  &  n_n535 ) ;
 assign wire16045 = ( n_n4616 ) | ( n_n4619 ) | ( n_n4623 ) ;
 assign wire16046 = ( n_n4617 ) | ( n_n4628 ) | ( n_n4621 ) | ( n_n4630 ) ;
 assign wire16056 = ( n_n482  &  n_n522  &  wire10 ) | ( n_n482  &  wire10  &  n_n530 ) ;
 assign wire16057 = ( n_n482  &  wire10  &  n_n532 ) | ( n_n482  &  wire10  &  n_n528 ) ;
 assign wire16064 = ( n_n4632 ) | ( wire15132 ) | ( _28731 ) ;
 assign wire16069 = ( n_n4560 ) | ( n_n4551 ) | ( wire471 ) | ( wire91 ) ;
 assign wire16075 = ( i_9_  &  n_n536  &  n_n509  &  n_n530 ) | ( (~ i_9_)  &  n_n536  &  n_n509  &  n_n530 ) ;
 assign wire16077 = ( n_n4344 ) | ( n_n4347 ) | ( wire53 ) ;
 assign wire16078 = ( n_n4335 ) | ( wire124 ) | ( wire16075 ) ;
 assign wire16081 = ( wire171 ) | ( wire364 ) ;
 assign wire16082 = ( n_n4334 ) | ( wire106 ) | ( wire677 ) ;
 assign wire16083 = ( n_n4331 ) | ( n_n4318 ) | ( n_n4313 ) | ( n_n4326 ) ;
 assign wire16088 = ( n_n522  &  wire16  &  n_n500 ) | ( wire16  &  n_n520  &  n_n500 ) ;
 assign wire16091 = ( n_n4380 ) | ( wire280 ) | ( n_n4377 ) ;
 assign wire16093 = ( n_n473  &  n_n524  &  wire16 ) | ( n_n473  &  wire16  &  n_n528 ) ;
 assign wire16102 = ( n_n4405 ) | ( n_n4406 ) | ( n_n4411 ) ;
 assign wire16103 = ( n_n4401 ) | ( n_n4409 ) | ( n_n4410 ) | ( n_n4402 ) ;
 assign wire16109 = ( n_n4357 ) | ( n_n4358 ) | ( n_n4354 ) ;
 assign wire16110 = ( n_n4359 ) | ( n_n4356 ) | ( _28790 ) ;
 assign wire16112 = ( n_n4350 ) | ( n_n4355 ) | ( wire16109 ) | ( wire16110 ) ;
 assign wire16119 = ( n_n4735 ) | ( n_n4744 ) | ( wire374 ) ;
 assign wire16120 = ( n_n4734 ) | ( n_n4729 ) | ( n_n4728 ) | ( wire373 ) ;
 assign wire16121 = ( wire15  &  n_n325  &  n_n500 ) | ( wire21  &  n_n325  &  n_n500 ) ;
 assign wire16124 = ( n_n4756 ) | ( n_n4753 ) | ( wire16121 ) ;
 assign wire16125 = ( wire109 ) | ( n_n4747 ) | ( n_n4752 ) | ( n_n4745 ) ;
 assign wire16130 = ( n_n4720 ) | ( n_n4719 ) | ( wire173 ) | ( _28427 ) ;
 assign wire16131 = ( wire16119 ) | ( wire16120 ) | ( wire16124 ) | ( wire16125 ) ;
 assign wire16132 = ( wire25  &  n_n325  &  n_n535 ) | ( wire15  &  n_n325  &  n_n535 ) ;
 assign wire16134 = ( wire221 ) | ( wire445 ) ;
 assign wire16135 = ( n_n4692 ) | ( n_n4695 ) | ( n_n4696 ) | ( wire16132 ) ;
 assign wire16139 = ( n_n4683 ) | ( n_n4684 ) | ( n_n4680 ) ;
 assign wire16140 = ( n_n4685 ) | ( n_n4686 ) | ( wire80 ) ;
 assign wire16141 = ( n_n4689 ) | ( n_n4712 ) | ( n_n4681 ) | ( n_n4705 ) ;
 assign wire16144 = ( n_n4219 ) | ( wire16139 ) | ( _28441 ) ;
 assign wire16145 = ( wire16134 ) | ( wire16135 ) | ( wire16140 ) | ( wire16141 ) ;
 assign wire16146 = ( n_n526  &  n_n509  &  wire18 ) | ( n_n522  &  n_n509  &  wire18 ) ;
 assign wire16148 = ( n_n4988 ) | ( n_n4987 ) | ( wire16146 ) ;
 assign wire16149 = ( n_n4999 ) | ( n_n4986 ) | ( n_n4989 ) | ( wire13997 ) ;
 assign wire16152 = ( wire252 ) | ( wire393 ) ;
 assign wire16153 = ( n_n4983 ) | ( n_n4984 ) | ( wire228 ) ;
 assign wire16155 = ( n_n4979 ) | ( n_n4985 ) | ( wire12255 ) | ( wire12256 ) ;
 assign wire16166 = ( n_n4907 ) | ( n_n4942 ) | ( n_n4936 ) | ( n_n4933 ) ;
 assign wire16171 = ( wire13867 ) | ( wire14962 ) | ( _28355 ) ;
 assign wire16174 = ( n_n4959 ) | ( n_n4960 ) | ( wire141 ) ;
 assign wire16175 = ( n_n4962 ) | ( n_n4971 ) | ( n_n4973 ) | ( wire11809 ) ;
 assign wire16179 = ( wire16171 ) | ( wire16174 ) | ( _28359 ) ;
 assign wire16182 = ( n_n491  &  wire11  &  n_n260 ) | ( n_n491  &  n_n260  &  wire23 ) ;
 assign wire16184 = ( n_n4898 ) | ( wire352 ) | ( n_n4897 ) ;
 assign wire16185 = ( wire96 ) | ( n_n4901 ) | ( wire16182 ) ;
 assign wire16186 = ( n_n473  &  n_n526  &  wire14 ) | ( n_n473  &  wire14  &  n_n520 ) ;
 assign wire16192 = ( i_9_  &  n_n534  &  n_n535  &  n_n260 ) | ( (~ i_9_)  &  n_n534  &  n_n535  &  n_n260 ) ;
 assign wire16195 = ( n_n4832 ) | ( n_n4812 ) | ( wire16192 ) ;
 assign wire16201 = ( i_9_  &  n_n518  &  n_n260  &  n_n520 ) | ( (~ i_9_)  &  n_n518  &  n_n260  &  n_n520 ) ;
 assign wire16203 = ( n_n4857 ) | ( n_n4858 ) | ( wire375 ) ;
 assign wire16204 = ( n_n4848 ) | ( wire52 ) | ( wire16201 ) ;
 assign wire16206 = ( n_n4862 ) | ( wire40 ) | ( n_n4861 ) ;
 assign wire16207 = ( n_n4859 ) | ( n_n4864 ) | ( n_n4866 ) | ( wire13810 ) ;
 assign wire16211 = ( n_n4835 ) | ( n_n4843 ) | ( n_n4839 ) | ( n_n4840 ) ;
 assign wire16215 = ( i_9_  &  n_n528  &  n_n260  &  n_n500 ) | ( (~ i_9_)  &  n_n528  &  n_n260  &  n_n500 ) ;
 assign wire16222 = ( n_n1985 ) | ( wire264 ) | ( wire261 ) | ( _28406 ) ;
 assign wire16229 = ( n_n4789 ) | ( n_n4793 ) | ( n_n4797 ) | ( wire179 ) ;
 assign wire16236 = ( n_n4782 ) | ( n_n4777 ) | ( n_n4788 ) ;
 assign wire16238 = ( n_n4204 ) | ( n_n3469 ) | ( wire16236 ) ;
 assign wire16245 = ( n_n5161 ) | ( n_n5162 ) | ( n_n5163 ) ;
 assign wire16246 = ( n_n482  &  n_n520  &  wire12 ) | ( n_n482  &  wire12  &  n_n530 ) ;
 assign wire16248 = ( wire437 ) | ( wire332 ) ;
 assign wire16249 = ( wire254 ) | ( n_n5170 ) | ( wire16246 ) ;
 assign wire16251 = ( n_n473  &  wire22  &  n_n130 ) | ( n_n473  &  wire11  &  n_n130 ) ;
 assign wire16253 = ( n_n5181 ) | ( n_n5184 ) | ( n_n5175 ) | ( n_n5177 ) ;
 assign wire16254 = ( wire112 ) | ( n_n5182 ) | ( wire16251 ) ;
 assign wire16256 = ( wire22  &  n_n464  &  n_n130 ) | ( n_n464  &  wire11  &  n_n130 ) ;
 assign wire16257 = ( wire220 ) | ( wire454 ) ;
 assign wire16258 = ( n_n5191 ) | ( wire452 ) | ( n_n5192 ) ;
 assign wire16259 = ( n_n5212 ) | ( n_n5189 ) | ( wire16256 ) ;
 assign wire16270 = ( i_9_  &  n_n65  &  n_n518  &  n_n534 ) | ( (~ i_9_)  &  n_n65  &  n_n518  &  n_n534 ) ;
 assign wire16278 = ( n_n5258 ) | ( n_n5251 ) | ( n_n5249 ) | ( n_n5252 ) ;
 assign wire16279 = ( n_n5259 ) | ( wire409 ) | ( n_n5247 ) | ( n_n5250 ) ;
 assign wire16282 = ( n_n491  &  n_n524  &  wire12 ) | ( n_n491  &  n_n532  &  wire12 ) ;
 assign wire16286 = ( n_n5150 ) | ( n_n5147 ) | ( wire196 ) | ( n_n5148 ) ;
 assign wire16288 = ( wire466 ) | ( wire16245 ) | ( wire16248 ) | ( wire16249 ) ;
 assign wire16293 = ( wire19  &  n_n491  &  n_n528 ) | ( wire19  &  n_n491  &  n_n530 ) ;
 assign wire16294 = ( n_n65  &  n_n491  &  wire22 ) | ( n_n65  &  n_n491  &  wire23 ) ;
 assign wire16297 = ( wire441 ) | ( n_n5279 ) | ( wire16294 ) ;
 assign wire16306 = ( wire25  &  n_n473  &  n_n65 ) | ( n_n473  &  n_n65  &  wire15 ) ;
 assign wire16308 = ( n_n5307 ) | ( n_n5308 ) | ( wire63 ) ;
 assign wire16309 = ( wire269 ) | ( n_n5304 ) | ( wire16306 ) ;
 assign wire16310 = ( wire19  &  n_n522  &  n_n464 ) | ( wire19  &  n_n464  &  n_n528 ) ;
 assign wire16312 = ( n_n5318 ) | ( n_n5320 ) | ( n_n5330 ) ;
 assign wire16313 = ( n_n5329 ) | ( n_n5319 ) | ( wire16310 ) ;
 assign wire16320 = ( n_n1786 ) | ( n_n1801 ) | ( n_n1800 ) | ( wire15991 ) ;
 assign wire16339 = ( n_n4877 ) | ( n_n4870 ) | ( n_n4872 ) ;
 assign wire16340 = ( n_n4881 ) | ( n_n4878 ) | ( wire174 ) ;
 assign wire16345 = ( n_n473  &  n_n522  &  wire14 ) | ( n_n473  &  n_n532  &  wire14 ) ;
 assign wire16346 = ( wire25  &  n_n473  &  n_n325 ) | ( n_n473  &  wire24  &  n_n325 ) ;
 assign wire16347 = ( i_9_  &  n_n473  &  n_n325  &  n_n530 ) | ( (~ i_9_)  &  n_n473  &  n_n325  &  n_n530 ) ;
 assign wire16349 = ( wire16345 ) | ( wire16346 ) ;
 assign wire16350 = ( n_n4791 ) | ( n_n4798 ) | ( n_n4801 ) | ( wire16347 ) ;
 assign wire16360 = ( n_n522  &  n_n464  &  wire14 ) | ( n_n524  &  n_n464  &  wire14 ) ;
 assign wire16366 = ( n_n491  &  wire11  &  n_n325 ) | ( n_n491  &  wire24  &  n_n325 ) ;
 assign wire16367 = ( wire164 ) | ( n_n4765 ) | ( n_n4766 ) ;
 assign wire16368 = ( n_n4770 ) | ( n_n4773 ) | ( n_n4771 ) | ( wire16366 ) ;
 assign wire16373 = ( n_n4776 ) | ( n_n4774 ) | ( n_n4786 ) | ( wire131 ) ;
 assign wire16378 = ( i_9_  &  n_n325  &  n_n500  &  n_n530 ) | ( (~ i_9_)  &  n_n325  &  n_n500  &  n_n530 ) ;
 assign wire16379 = ( wire22  &  n_n325  &  n_n500 ) | ( wire24  &  n_n325  &  n_n500 ) ;
 assign wire16382 = ( wire16378 ) | ( wire16379 ) ;
 assign wire16383 = ( wire373 ) | ( n_n4752 ) | ( n_n4751 ) | ( n_n4750 ) ;
 assign wire16385 = ( n_n4732 ) | ( wire293 ) | ( wire767 ) ;
 assign wire16386 = ( n_n4738 ) | ( wire95 ) | ( n_n4733 ) | ( n_n4736 ) ;
 assign wire16396 = ( n_n4709 ) | ( n_n4698 ) | ( n_n4707 ) | ( n_n4702 ) ;
 assign wire16408 = ( n_n482  &  n_n522  &  wire10 ) | ( n_n482  &  n_n524  &  wire10 ) ;
 assign wire16409 = ( n_n526  &  n_n464  &  wire10 ) | ( n_n464  &  wire10  &  n_n528 ) ;
 assign wire16412 = ( n_n4667 ) | ( n_n4664 ) | ( n_n4663 ) | ( wire16409 ) ;
 assign wire16420 = ( n_n4758 ) | ( n_n4761 ) | ( n_n4762 ) ;
 assign wire16421 = ( n_n4754 ) | ( n_n4757 ) | ( n_n4756 ) | ( n_n4755 ) ;
 assign wire16427 = ( i_9_  &  n_n509  &  n_n520  &  n_n195 ) | ( (~ i_9_)  &  n_n509  &  n_n520  &  n_n195 ) ;
 assign wire16430 = ( wire393 ) | ( wire16427 ) ;
 assign wire16431 = ( n_n4994 ) | ( n_n5004 ) | ( wire136 ) | ( n_n5001 ) ;
 assign wire16435 = ( n_n5018 ) | ( n_n5015 ) | ( wire343 ) ;
 assign wire16436 = ( n_n5016 ) | ( n_n5009 ) | ( n_n5013 ) | ( wire297 ) ;
 assign wire16438 = ( i_9_  &  n_n534  &  n_n509  &  n_n195 ) | ( (~ i_9_)  &  n_n534  &  n_n509  &  n_n195 ) ;
 assign wire16442 = ( n_n4986 ) | ( wire251 ) | ( _29219 ) ;
 assign wire16443 = ( wire16430 ) | ( wire16431 ) | ( wire16435 ) | ( wire16436 ) ;
 assign wire16447 = ( wire15  &  n_n482  &  n_n260 ) | ( n_n482  &  wire11  &  n_n260 ) ;
 assign wire16448 = ( n_n491  &  n_n260  &  wire20 ) | ( n_n491  &  n_n260  &  wire23 ) ;
 assign wire16453 = ( n_n4913 ) | ( n_n4914 ) | ( n_n4915 ) ;
 assign wire16454 = ( n_n4920 ) | ( n_n4923 ) | ( n_n4918 ) | ( n_n4917 ) ;
 assign wire16461 = ( n_n4966 ) | ( n_n4978 ) | ( wire228 ) | ( n_n4972 ) ;
 assign wire16462 = ( wire21  &  n_n535  &  n_n195 ) | ( wire11  &  n_n535  &  n_n195 ) ;
 assign wire16463 = ( n_n526  &  n_n535  &  wire18 ) | ( n_n522  &  n_n535  &  wire18 ) ;
 assign wire16465 = ( n_n4953 ) | ( wire14752 ) | ( wire16463 ) ;
 assign wire16468 = ( n_n2222 ) | ( wire16465 ) | ( _29241 ) | ( _29242 ) ;
 assign wire16470 = ( n_n2177 ) | ( wire16442 ) | ( wire16443 ) | ( wire16468 ) ;
 assign wire16479 = ( n_n526  &  wire13  &  n_n500 ) | ( wire13  &  n_n500  &  n_n530 ) ;
 assign wire16480 = ( wire13  &  n_n532  &  n_n509 ) | ( wire13  &  n_n509  &  n_n520 ) ;
 assign wire16482 = ( n_n4513 ) | ( n_n4518 ) | ( wire16479 ) ;
 assign wire16483 = ( n_n4484 ) | ( wire199 ) | ( wire16480 ) ;
 assign wire16487 = ( n_n4617 ) | ( n_n4612 ) | ( wire239 ) ;
 assign wire16488 = ( n_n4640 ) | ( n_n4581 ) | ( wire256 ) | ( n_n4623 ) ;
 assign wire16490 = ( n_n473  &  wire21  &  n_n455 ) | ( n_n473  &  n_n455  &  wire24 ) ;
 assign wire16498 = ( n_n522  &  n_n491  &  wire14 ) | ( n_n491  &  wire14  &  n_n530 ) ;
 assign wire16500 = ( n_n522  &  n_n509  &  wire14 ) | ( n_n522  &  wire14  &  n_n535 ) ;
 assign wire16506 = ( n_n473  &  wire21  &  n_n390 ) | ( n_n482  &  wire21  &  n_n390 ) ;
 assign wire16514 = ( n_n4800 ) | ( n_n4803 ) | ( n_n4783 ) | ( n_n4812 ) ;
 assign wire16518 = ( n_n473  &  wire22  &  n_n536 ) | ( n_n473  &  wire21  &  n_n536 ) ;
 assign wire16531 = ( _29003 ) | ( _29004 ) ;
 assign wire16537 = ( n_n4353 ) | ( wire399 ) | ( n_n4354 ) ;
 assign wire16538 = ( n_n4343 ) | ( n_n4352 ) | ( wire67 ) | ( n_n4349 ) ;
 assign wire16539 = ( _72 ) | ( wire15  &  n_n536  &  n_n535 ) ;
 assign wire16544 = ( n_n4336 ) | ( wire171 ) | ( wire198 ) | ( wire283 ) ;
 assign wire16548 = ( n_n4355 ) | ( n_n4356 ) | ( wire345 ) ;
 assign wire16549 = ( n_n4363 ) | ( n_n4359 ) | ( n_n4365 ) | ( wire13055 ) ;
 assign wire16551 = ( n_n4379 ) | ( n_n4372 ) | ( n_n4371 ) ;
 assign wire16552 = ( n_n4382 ) | ( n_n4373 ) | ( wire423 ) ;
 assign wire16556 = ( wire16548 ) | ( wire16549 ) | ( wire16551 ) | ( wire16552 ) ;
 assign wire16560 = ( wire13  &  n_n532  &  n_n535 ) | ( wire13  &  n_n535  &  n_n530 ) ;
 assign wire16562 = ( n_n4450 ) | ( n_n4445 ) | ( wire368 ) ;
 assign wire16563 = ( n_n4441 ) | ( n_n4448 ) | ( n_n4447 ) | ( wire16560 ) ;
 assign wire16566 = ( n_n4464 ) | ( n_n4463 ) | ( n_n4466 ) ;
 assign wire16567 = ( n_n4468 ) | ( n_n4472 ) | ( _29270 ) ;
 assign wire16568 = ( n_n4459 ) | ( n_n4470 ) | ( n_n4460 ) | ( n_n4473 ) ;
 assign wire16570 = ( n_n4454 ) | ( wire11520 ) | ( wire14517 ) | ( wire16568 ) ;
 assign wire16571 = ( wire16562 ) | ( wire16563 ) | ( wire16566 ) | ( wire16567 ) ;
 assign wire16572 = ( wire22  &  n_n455  &  n_n500 ) | ( n_n455  &  wire24  &  n_n500 ) ;
 assign wire16574 = ( n_n4488 ) | ( n_n4489 ) | ( n_n4490 ) | ( wire16572 ) ;
 assign wire16578 = ( n_n482  &  n_n455  &  wire20 ) | ( n_n482  &  n_n455  &  wire23 ) ;
 assign wire16580 = ( wire416 ) | ( wire16578 ) ;
 assign wire16581 = ( n_n4536 ) | ( n_n4532 ) | ( n_n4541 ) | ( wire13090 ) ;
 assign wire16585 = ( n_n4520 ) | ( n_n4529 ) | ( wire789 ) | ( wire724 ) ;
 assign wire16586 = ( wire361 ) | ( wire378 ) ;
 assign wire16587 = ( n_n4512 ) | ( n_n4522 ) | ( n_n4531 ) | ( n_n4517 ) ;
 assign wire16590 = ( n_n4247 ) | ( wire308 ) | ( n_n4528 ) | ( wire16587 ) ;
 assign wire16591 = ( wire16580 ) | ( wire16581 ) | ( wire16585 ) | ( wire16586 ) ;
 assign wire16593 = ( n_n522  &  wire13  &  n_n500 ) | ( wire13  &  n_n520  &  n_n500 ) ;
 assign wire16594 = ( n_n4504 ) | ( n_n4503 ) | ( n_n4506 ) | ( n_n4505 ) ;
 assign wire16596 = ( n_n4508 ) | ( wire13028 ) | ( wire16593 ) | ( wire16594 ) ;
 assign wire16598 = ( wire16576 ) | ( wire16596 ) | ( _29247 ) | ( _29258 ) ;
 assign wire16599 = ( wire16570 ) | ( wire16571 ) | ( wire16590 ) | ( wire16591 ) ;
 assign wire16601 = ( n_n4570 ) | ( n_n4569 ) | ( wire455 ) ;
 assign wire16602 = ( n_n4561 ) | ( n_n4568 ) | ( wire471 ) | ( wire91 ) ;
 assign wire16603 = ( i_9_  &  n_n526  &  n_n390  &  n_n535 ) | ( (~ i_9_)  &  n_n526  &  n_n390  &  n_n535 ) ;
 assign wire16605 = ( wire238 ) | ( wire276 ) ;
 assign wire16606 = ( n_n4584 ) | ( n_n4583 ) | ( n_n4580 ) | ( wire16603 ) ;
 assign wire16609 = ( n_n526  &  wire10  &  n_n509 ) | ( wire10  &  n_n509  &  n_n520 ) ;
 assign wire16611 = ( n_n4616 ) | ( n_n4607 ) | ( n_n4618 ) | ( n_n4611 ) ;
 assign wire16612 = ( n_n4613 ) | ( n_n4610 ) | ( n_n4609 ) | ( wire16609 ) ;
 assign wire16617 = ( n_n4598 ) | ( n_n4601 ) | ( n_n4594 ) | ( n_n4606 ) ;
 assign wire16618 = ( n_n4605 ) | ( n_n4600 ) | ( n_n4603 ) | ( wire255 ) ;
 assign wire16621 = ( n_n4593 ) | ( n_n4590 ) | ( n_n4585 ) | ( wire12520 ) ;
 assign wire16623 = ( wire16611 ) | ( wire16612 ) | ( wire16617 ) | ( wire16618 ) ;
 assign wire16627 = ( n_n4648 ) | ( n_n4646 ) | ( wire311 ) ;
 assign wire16628 = ( wire309 ) | ( n_n4644 ) | ( n_n4651 ) | ( n_n4649 ) ;
 assign wire16629 = ( n_n522  &  wire10  &  n_n500 ) | ( wire10  &  n_n500  &  n_n530 ) ;
 assign wire16631 = ( n_n4629 ) | ( n_n4630 ) | ( wire190 ) ;
 assign wire16632 = ( wire118 ) | ( n_n4626 ) | ( wire16629 ) ;
 assign wire16633 = ( wire25  &  n_n491  &  n_n390 ) | ( n_n491  &  wire22  &  n_n390 ) ;
 assign wire16635 = ( n_n4637 ) | ( n_n4634 ) | ( n_n4638 ) | ( n_n4631 ) ;
 assign wire16636 = ( n_n4642 ) | ( wire16633 ) | ( _29324 ) ;
 assign wire16638 = ( wire16627 ) | ( wire16628 ) | ( wire16631 ) | ( wire16632 ) ;
 assign wire16641 = ( n_n4551 ) | ( n_n4552 ) | ( wire213 ) ;
 assign wire16642 = ( n_n4554 ) | ( wire212 ) | ( n_n4546 ) | ( n_n4555 ) ;
 assign wire16644 = ( wire16601 ) | ( wire16602 ) | ( wire16605 ) | ( wire16606 ) ;
 assign wire16645 = ( wire16641 ) | ( wire16642 ) | ( wire16644 ) ;
 assign wire16646 = ( wire16623 ) | ( wire16638 ) | ( _29335 ) ;
 assign wire16656 = ( wire148 ) | ( n_n5318 ) | ( n_n5320 ) ;
 assign wire16657 = ( n_n5321 ) | ( n_n5307 ) | ( wire269 ) ;
 assign wire16658 = ( n_n5326 ) | ( n_n5325 ) | ( n_n5332 ) | ( n_n5329 ) ;
 assign wire16662 = ( n_n2274 ) | ( wire16656 ) | ( wire16657 ) | ( wire16658 ) ;
 assign wire16663 = ( n_n526  &  n_n491  &  wire12 ) | ( n_n491  &  n_n520  &  wire12 ) ;
 assign wire16666 = ( wire76 ) | ( n_n5140 ) | ( wire16663 ) ;
 assign wire16670 = ( n_n5171 ) | ( wire114 ) | ( n_n5181 ) | ( n_n5177 ) ;
 assign wire16673 = ( n_n5191 ) | ( wire113 ) | ( n_n5192 ) ;
 assign wire16674 = ( n_n5183 ) | ( wire112 ) | ( n_n5190 ) | ( n_n5188 ) ;
 assign wire16676 = ( wire15  &  n_n464  &  n_n130 ) | ( n_n464  &  wire24  &  n_n130 ) ;
 assign wire16677 = ( wire220 ) | ( wire454 ) ;
 assign wire16678 = ( n_n5201 ) | ( wire451 ) | ( wire761 ) ;
 assign wire16679 = ( n_n5212 ) | ( n_n5203 ) | ( wire16676 ) ;
 assign wire16690 = ( i_9_  &  n_n65  &  n_n524  &  n_n518 ) | ( (~ i_9_)  &  n_n65  &  n_n524  &  n_n518 ) ;
 assign wire16693 = ( n_n5260 ) | ( n_n5226 ) | ( wire16690 ) ;
 assign wire16698 = ( n_n482  &  n_n532  &  wire12 ) | ( n_n482  &  n_n528  &  wire12 ) ;
 assign wire16699 = ( n_n482  &  wire22  &  n_n130 ) | ( n_n482  &  wire24  &  n_n130 ) ;
 assign wire16702 = ( wire33 ) | ( n_n5170 ) | ( wire16699 ) ;
 assign wire16704 = ( wire16666 ) | ( wire16670 ) | ( _28879 ) ;
 assign wire16709 = ( n_n5066 ) | ( n_n5063 ) | ( n_n5068 ) ;
 assign wire16710 = ( wire123 ) | ( wire159 ) ;
 assign wire16711 = ( n_n5064 ) | ( n_n5082 ) | ( _28900 ) ;
 assign wire16715 = ( n_n4152 ) | ( n_n5079 ) | ( n_n5083 ) | ( wire144 ) ;
 assign wire16716 = ( wire90 ) | ( wire16709 ) | ( wire16710 ) | ( wire16711 ) ;
 assign wire16717 = ( n_n518  &  n_n534  &  wire12 ) | ( n_n518  &  wire12  &  n_n530 ) ;
 assign wire16718 = ( n_n5098 ) | ( wire289 ) | ( n_n5095 ) ;
 assign wire16719 = ( n_n5108 ) | ( wire16717 ) | ( _28912 ) ;
 assign wire16721 = ( n_n532  &  n_n509  &  wire12 ) | ( n_n509  &  wire12  &  n_n530 ) ;
 assign wire16723 = ( n_n5111 ) | ( n_n5113 ) | ( wire414 ) ;
 assign wire16724 = ( n_n5112 ) | ( n_n5110 ) | ( n_n5115 ) | ( wire16721 ) ;
 assign wire16728 = ( n_n5136 ) | ( n_n5127 ) | ( n_n5128 ) | ( n_n5135 ) ;
 assign wire16730 = ( n_n5139 ) | ( n_n5125 ) | ( n_n2304 ) | ( wire16728 ) ;
 assign wire16731 = ( wire16718 ) | ( wire16719 ) | ( wire16723 ) | ( wire16724 ) ;
 assign wire16739 = ( n_n5050 ) | ( n_n5049 ) | ( n_n5043 ) | ( n_n5044 ) ;
 assign wire16740 = ( n_n5040 ) | ( n_n5048 ) | ( n_n5036 ) | ( n_n5047 ) ;
 assign wire16742 = ( n_n5039 ) | ( n_n5029 ) | ( wire16739 ) | ( wire16740 ) ;
 assign wire16755 = ( n_n5274 ) | ( n_n5266 ) | ( n_n5275 ) | ( n_n5261 ) ;
 assign wire16760 = ( i_9_  &  n_n65  &  n_n464  &  n_n520 ) | ( (~ i_9_)  &  n_n65  &  n_n464  &  n_n520 ) ;
 assign wire16761 = ( wire16760 ) | ( n_n65  &  n_n464  &  wire20 ) ;
 assign wire16769 = ( n_n4432 ) | ( n_n4461 ) | ( n_n4438 ) | ( n_n4421 ) ;
 assign wire16770 = ( wire84 ) | ( n_n4465 ) | ( n_n4443 ) | ( n_n4429 ) ;
 assign wire16773 = ( n_n65  &  wire22  &  n_n518 ) | ( n_n65  &  wire22  &  n_n509 ) ;
 assign wire16788 = ( n_n526  &  n_n518  &  wire12 ) | ( n_n524  &  n_n518  &  wire12 ) ;
 assign wire16798 = ( n_n518  &  wire11  &  n_n195 ) | ( wire11  &  n_n509  &  n_n195 ) ;
 assign wire16799 = ( n_n526  &  n_n509  &  wire18 ) | ( n_n522  &  n_n509  &  wire18 ) ;
 assign wire16804 = ( n_n5000 ) | ( n_n4957 ) | ( n_n4973 ) | ( wire16798 ) ;
 assign wire16818 = ( n_n4934 ) | ( n_n4938 ) | ( n_n4947 ) | ( n_n4940 ) ;
 assign wire16819 = ( n_n4931 ) | ( n_n4944 ) | ( n_n4932 ) | ( wire340 ) ;
 assign wire16820 = ( wire16818 ) | ( wire16819 ) ;
 assign wire16823 = ( n_n2083 ) | ( n_n2095 ) | ( n_n2096 ) | ( wire16820 ) ;
 assign wire16825 = ( n_n2104 ) | ( wire16651 ) | ( _29086 ) | ( _29091 ) ;
 assign wire16827 = ( n_n2084 ) | ( wire16823 ) | ( wire16825 ) ;
 assign wire16829 = ( wire16598 ) | ( wire16599 ) | ( wire16645 ) | ( wire16646 ) ;
 assign _38 = ( n_n473  &  n_n260  &  wire23 ) ;
 assign _64 = ( wire19  &  n_n528  &  n_n500 ) ;
 assign _72 = ( wire16  &  n_n534  &  n_n535 ) ;
 assign _90 = ( n_n526  &  n_n464  &  wire13 ) ;
 assign _120 = ( n_n536  &  wire23  &  n_n500 ) ;
 assign _144 = ( n_n455  &  wire11  &  n_n509 ) ;
 assign _172 = ( wire19  &  n_n464  &  n_n532 ) ;
 assign _198 = ( wire25  &  n_n65  &  n_n500 ) ;
 assign _204 = ( wire21  &  n_n325  &  n_n535 ) ;
 assign _206 = ( wire14  &  n_n535  &  n_n520 ) ;
 assign _220 = ( n_n464  &  wire17  &  n_n520 ) ;
 assign _226 = ( n_n473  &  n_n65  &  wire20 ) ;
 assign _230 = ( n_n65  &  n_n491  &  wire20 ) ;
 assign _298 = ( n_n464  &  n_n325  &  wire20 ) ;
 assign _348 = ( n_n65  &  n_n518  &  wire21 ) ;
 assign _356 = ( n_n491  &  n_n325  &  wire20 ) ;
 assign _362 = ( wire25  &  n_n518  &  n_n325 ) ;
 assign _364 = ( n_n534  &  n_n509  &  wire14 ) ;
 assign _388 = ( n_n491  &  n_n528  &  wire17 ) ;
 assign _462 = ( n_n464  &  n_n455  &  wire24 ) ;
 assign _514 = ( n_n473  &  n_n522  &  wire12 ) ;
 assign _560 = ( n_n532  &  n_n509  &  wire17 ) ;
 assign _564 = ( n_n482  &  wire11  &  n_n325 ) ;
 assign _600 = ( n_n518  &  wire13  &  n_n532 ) ;
 assign _660 = ( wire17  &  n_n535  &  n_n520 ) ;
 assign _664 = ( n_n491  &  wire14  &  n_n530 ) ;
 assign _670 = ( n_n518  &  wire11  &  n_n325 ) ;
 assign _672 = ( wire21  &  n_n325  &  n_n535 ) ;
 assign _690 = ( n_n482  &  n_n528  &  wire17 ) ;
 assign _708 = ( n_n536  &  wire24  &  n_n535 ) ;
 assign _778 = ( n_n65  &  n_n482  &  wire24 ) ;
 assign _904 = ( n_n535  &  n_n260  &  wire20 ) ;
 assign _930 = ( n_n455  &  wire23  &  n_n500 ) ;
 assign _932 = ( n_n482  &  wire13  &  n_n530 ) ;
 assign _1018 = ( n_n522  &  n_n464  &  wire13 ) ;
 assign _1050 = ( n_n491  &  wire22  &  n_n455 ) ;
 assign _1120 = ( wire19  &  n_n522  &  n_n535 ) ;
 assign _1152 = ( n_n473  &  wire22  &  n_n260 ) ;
 assign _1160 = ( n_n491  &  wire21  &  n_n325 ) ;
 assign _1176 = ( n_n526  &  wire17  &  n_n500 ) ;
 assign _1190 = ( wire19  &  n_n491  &  n_n520 ) ;
 assign _1204 = ( n_n65  &  n_n482  &  wire21 ) ;
 assign _1230 = ( n_n65  &  wire21  &  n_n535 ) ;
 assign _1240 = ( wire12  &  n_n500  &  n_n530 ) ;
 assign _1244 = ( wire11  &  n_n195  &  n_n500 ) ;
 assign _1366 = ( n_n526  &  wire14  &  n_n500 ) ;
 assign _1394 = ( n_n464  &  n_n455  &  wire600 ) ;
 assign _1428 = ( n_n526  &  wire13  &  n_n535 ) ;
 assign _1490 = ( n_n536  &  wire23  &  n_n500 ) ;
 assign _1514 = ( n_n491  &  n_n536  &  wire23 ) ;
 assign _1694 = ( n_n518  &  n_n520  &  wire18 ) ;
 assign _22059 = ( n_n526  &  n_n518  &  wire14 ) | ( n_n524  &  n_n518  &  wire14 ) ;
 assign _22066 = ( wire95 ) | ( n_n526  &  n_n509  &  wire14 ) ;
 assign _22147 = ( n_n4674 ) | ( n_n473  &  n_n390  &  wire20 ) ;
 assign _22149 = ( n_n4663 ) | ( wire225 ) | ( wire11856 ) | ( wire11859 ) ;
 assign _22150 = ( wire11855 ) | ( wire11880 ) | ( wire11881 ) | ( _22147 ) ;
 assign _22151 = ( wire457 ) | ( wire11852 ) | ( wire11848 ) | ( _22066 ) ;
 assign _22193 = ( wire11825 ) | ( wire264 ) ;
 assign _22194 = ( wire295 ) | ( n_n4869 ) | ( n_n4870 ) | ( wire11824 ) ;
 assign _22212 = ( n_n4940 ) | ( n_n4939 ) | ( wire382 ) ;
 assign _22253 = ( wire11811 ) | ( wire11810 ) ;
 assign _22279 = ( wire11795 ) | ( wire11814 ) | ( _22212 ) | ( _22253 ) ;
 assign _22321 = ( wire21  &  n_n325  &  n_n500 ) | ( n_n325  &  wire23  &  n_n500 ) ;
 assign _22359 = ( n_n526  &  n_n464  &  wire14 ) | ( n_n464  &  wire14  &  n_n530 ) ;
 assign _22360 = ( n_n464  &  wire11  &  n_n325 ) | ( n_n464  &  wire24  &  n_n325 ) ;
 assign _22415 = ( wire11888 ) | ( wire11889 ) | ( wire11891 ) ;
 assign _22416 = ( wire11832 ) | ( wire11797 ) | ( wire11816 ) | ( _22279 ) ;
 assign _22433 = ( n_n5244 ) | ( n_n65  &  wire22  &  n_n509 ) ;
 assign _22464 = ( n_n5273 ) | ( wire19  &  n_n491  &  n_n528 ) ;
 assign _22478 = ( n_n65  &  n_n491  &  wire22 ) | ( n_n65  &  n_n491  &  wire11 ) ;
 assign _22494 = ( n_n5293 ) | ( n_n5294 ) | ( wire200 ) ;
 assign _22495 = ( wire11929 ) | ( n_n5280 ) | ( wire11928 ) | ( _22478 ) ;
 assign _22502 = ( n_n473  &  wire19  &  n_n528 ) | ( n_n473  &  wire19  &  n_n530 ) ;
 assign _22511 = ( n_n5303 ) | ( n_n5311 ) | ( n_n5309 ) | ( _22502 ) ;
 assign _22549 = ( n_n5240 ) | ( n_n5238 ) | ( wire11955 ) ;
 assign _22550 = ( wire11952 ) | ( wire11951 ) ;
 assign _22551 = ( wire11944 ) | ( wire11959 ) | ( _22511 ) | ( _22549 ) ;
 assign _22552 = ( n_n1050 ) | ( wire409 ) | ( wire11923 ) | ( wire11927 ) ;
 assign _22574 = ( wire25  &  n_n535  &  n_n130 ) | ( wire22  &  n_n535  &  n_n130 ) ;
 assign _22575 = ( n_n532  &  n_n535  &  wire12 ) | ( n_n535  &  wire12  &  n_n530 ) ;
 assign _22614 = ( n_n5035 ) | ( n_n5036 ) | ( wire11997 ) | ( wire11999 ) ;
 assign _22691 = ( n_n4990 ) | ( wire12023 ) | ( wire12024 ) | ( _1694 ) ;
 assign _22692 = ( n_n5039 ) | ( wire253 ) | ( wire12004 ) | ( _22614 ) ;
 assign _22732 = ( wire422 ) | ( wire211 ) ;
 assign _22733 = ( wire28 ) | ( wire11916 ) | ( wire11917 ) ;
 assign _22749 = ( n_n473  &  n_n534  &  wire12 ) | ( n_n473  &  wire12  &  n_n530 ) ;
 assign _22752 = ( n_n5181 ) | ( n_n5173 ) | ( wire11902 ) ;
 assign _22800 = ( wire220 ) | ( n_n65  &  wire24  &  n_n535 ) ;
 assign _22801 = ( n_n5201 ) | ( wire761 ) | ( wire11972 ) | ( wire11973 ) ;
 assign _22829 = ( wire11906 ) | ( _22752 ) | ( _22800 ) | ( _22801 ) ;
 assign _22846 = ( n_n4460 ) | ( wire25  &  n_n518  &  n_n455 ) ;
 assign _22891 = ( wire170 ) | ( n_n482  &  wire13  &  n_n530 ) ;
 assign _22972 = ( wire84 ) | ( wire79 ) | ( wire11527 ) ;
 assign _22973 = ( wire11502 ) | ( wire11495 ) | ( wire11498 ) | ( _22891 ) ;
 assign _22987 = ( n_n4555 ) | ( n_n464  &  wire13  &  n_n530 ) ;
 assign _23016 = ( n_n4525 ) | ( n_n4528 ) | ( n_n4529 ) ;
 assign _23017 = ( n_n4542 ) | ( wire201 ) | ( wire11535 ) | ( wire11536 ) ;
 assign _23150 = ( n_n4607 ) | ( n_n4641 ) | ( wire11642 ) | ( wire11638 ) ;
 assign _23316 = ( n_n4374 ) | ( wire21  &  n_n536  &  n_n535 ) ;
 assign _23327 = ( wire15  &  n_n482  &  n_n536 ) | ( n_n482  &  wire22  &  n_n536 ) ;
 assign _23360 = ( n_n4393 ) | ( n_n4402 ) | ( _1514 ) | ( _23327 ) ;
 assign _23446 = ( n_n518  &  n_n536  &  wire11 ) | ( n_n518  &  n_n536  &  wire20 ) ;
 assign _23478 = ( n_n4399 ) | ( n_n4428 ) | ( wire12461 ) ;
 assign _23479 = ( n_n4393 ) | ( wire37 ) | ( n_n4394 ) | ( wire12465 ) ;
 assign _23490 = ( n_n4361 ) | ( wire16  &  n_n509  &  n_n530 ) ;
 assign _23507 = ( wire21  &  n_n536  &  n_n509 ) | ( n_n536  &  n_n509  &  wire20 ) ;
 assign _23508 = ( n_n522  &  wire16  &  n_n509 ) | ( wire16  &  n_n509  &  n_n520 ) ;
 assign _23538 = ( wire283 ) | ( wire67 ) | ( wire364 ) | ( wire53 ) ;
 assign _23540 = ( n_n4323 ) | ( wire12569 ) | ( wire12578 ) | ( wire12579 ) ;
 assign _23541 = ( n_n3533 ) | ( wire12453 ) | ( wire12456 ) | ( _23490 ) ;
 assign _23543 = ( wire15  &  n_n455  &  n_n509 ) | ( n_n455  &  wire24  &  n_n509 ) ;
 assign _23548 = ( n_n4476 ) | ( n_n4471 ) | ( n_n4472 ) | ( _23543 ) ;
 assign _23567 = ( n_n4504 ) | ( n_n4503 ) | ( wire12510 ) ;
 assign _23568 = ( n_n4489 ) | ( wire66 ) | ( n_n4490 ) | ( wire12490 ) ;
 assign _23569 = ( wire12493 ) | ( wire12514 ) | ( _23548 ) | ( _23567 ) ;
 assign _23648 = ( wire15  &  n_n390  &  n_n509 ) | ( wire24  &  n_n390  &  n_n509 ) ;
 assign _23670 = ( wire256 ) | ( wire12561 ) | ( wire12564 ) ;
 assign _23708 = ( wire213 ) | ( wire276 ) | ( wire12521 ) | ( _1394 ) ;
 assign _23747 = ( wire12566 ) | ( _23568 ) | ( _23569 ) | ( _23670 ) ;
 assign _23753 = ( n_n4701 ) | ( wire14  &  n_n528  &  n_n535 ) ;
 assign _23780 = ( n_n4689 ) | ( n_n4684 ) | ( wire444 ) | ( wire12428 ) ;
 assign _23821 = ( n_n4755 ) | ( wire12435 ) | ( wire12436 ) | ( _1366 ) ;
 assign _23822 = ( wire12432 ) | ( n_n4693 ) | ( wire12422 ) | ( _23780 ) ;
 assign _23853 = ( n_n4491 ) | ( n_n4438 ) | ( wire184 ) | ( wire12054 ) ;
 assign _23965 = ( n_n473  &  n_n522  &  wire16 ) | ( n_n482  &  n_n522  &  wire16 ) ;
 assign _23986 = ( wire12147 ) | ( wire12146 ) ;
 assign _23987 = ( wire12108 ) | ( wire12109 ) | ( wire12111 ) ;
 assign _24115 = ( n_n4848 ) | ( n_n535  &  n_n260  &  wire23 ) ;
 assign _24138 = ( n_n4825 ) | ( wire186 ) | ( n_n4826 ) ;
 assign _24139 = ( n_n4827 ) | ( n_n4828 ) | ( wire12231 ) | ( wire12226 ) ;
 assign _24226 = ( wire12319 ) | ( wire12318 ) ;
 assign _24227 = ( n_n5054 ) | ( wire97 ) | ( n_n5042 ) | ( wire12316 ) ;
 assign _24250 = ( n_n518  &  wire21  &  n_n130 ) | ( n_n518  &  wire20  &  n_n130 ) ;
 assign _24258 = ( n_n5100 ) | ( n_n518  &  wire11  &  n_n130 ) ;
 assign _24270 = ( wire12256 ) | ( wire12255 ) ;
 assign _24285 = ( n_n5034 ) | ( n_n5027 ) | ( wire253 ) ;
 assign _24286 = ( wire296 ) | ( n_n5019 ) | ( n_n5020 ) | ( wire12253 ) ;
 assign _24317 = ( wire358 ) | ( wire406 ) | ( wire211 ) | ( wire288 ) ;
 assign _24320 = ( n_n5127 ) | ( wire12300 ) | ( wire12301 ) | ( _1240 ) ;
 assign _24373 = ( wire114 ) | ( wire113 ) | ( wire168 ) | ( wire437 ) ;
 assign _24405 = ( n_n5305 ) | ( n_n3019 ) | ( wire204 ) | ( _1204 ) ;
 assign _24444 = ( n_n65  &  n_n482  &  wire22 ) | ( n_n65  &  n_n482  &  wire24 ) ;
 assign _24445 = ( n_n482  &  wire19  &  n_n524 ) | ( n_n482  &  wire19  &  n_n530 ) ;
 assign _24448 = ( n_n482  &  wire19  &  n_n532 ) | ( n_n482  &  wire19  &  n_n534 ) ;
 assign _24456 = ( wire218 ) | ( _1190 ) | ( _24444 ) | ( _24445 ) ;
 assign _24460 = ( n_n1402 ) | ( wire12304 ) | ( _24320 ) | ( _24405 ) ;
 assign _24477 = ( n_n482  &  n_n526  &  wire14 ) | ( n_n482  &  wire14  &  n_n530 ) ;
 assign _24485 = ( wire380 ) | ( wire292 ) ;
 assign _24486 = ( n_n4783 ) | ( wire12762 ) | ( wire12760 ) | ( _24477 ) ;
 assign _24493 = ( wire12225 ) | ( n_n464  &  wire14  &  n_n528 ) ;
 assign _24526 = ( n_n4887 ) | ( wire12770 ) | ( wire12771 ) | ( _1176 ) ;
 assign _24527 = ( n_n834 ) | ( wire12753 ) | ( wire12749 ) | ( _24493 ) ;
 assign _24555 = ( n_n4663 ) | ( n_n482  &  wire10  &  n_n530 ) ;
 assign _24594 = ( wire12393 ) | ( n_n4204 ) | ( wire456 ) | ( _1160 ) ;
 assign _24595 = ( wire12814 ) | ( wire12810 ) | ( wire12811 ) | ( _24555 ) ;
 assign _24602 = ( n_n4921 ) | ( n_n473  &  n_n522  &  wire17 ) ;
 assign _24620 = ( n_n4920 ) | ( n_n4919 ) | ( wire340 ) ;
 assign _24621 = ( wire154 ) | ( n_n4896 ) | ( wire12722 ) | ( wire12724 ) ;
 assign _24749 = ( n_n5074 ) | ( n_n5082 ) | ( wire12909 ) ;
 assign _24750 = ( n_n5050 ) | ( n_n5049 ) | ( wire12908 ) | ( wire12904 ) ;
 assign _24759 = ( wire88 ) | ( wire12917 ) | ( wire12924 ) ;
 assign _24803 = ( wire297 ) | ( wire394 ) | ( wire265 ) | ( wire12935 ) ;
 assign _24805 = ( n_n5039 ) | ( wire231 ) | ( wire12941 ) | ( wire12943 ) ;
 assign _24806 = ( wire28 ) | ( wire12930 ) | ( _24759 ) ;
 assign _24831 = ( wire12949 ) | ( wire333 ) ;
 assign _24874 = ( wire22  &  n_n464  &  n_n130 ) | ( n_n464  &  wire20  &  n_n130 ) ;
 assign _24885 = ( n_n5181 ) | ( n_n5184 ) | ( wire107 ) | ( wire12996 ) ;
 assign _24886 = ( wire12952 ) | ( wire12960 ) | ( wire12961 ) | ( _24831 ) ;
 assign _24893 = ( wire13028 ) | ( n_n491  &  wire13  &  n_n530 ) ;
 assign _24946 = ( n_n518  &  wire21  &  n_n455 ) | ( n_n518  &  n_n455  &  wire11 ) ;
 assign _24947 = ( n_n522  &  n_n518  &  wire13 ) | ( n_n524  &  n_n518  &  wire13 ) ;
 assign _24948 = ( n_n4469 ) | ( n_n518  &  wire13  &  n_n528 ) ;
 assign _24968 = ( n_n482  &  wire22  &  n_n536 ) | ( n_n482  &  n_n536  &  wire20 ) ;
 assign _24971 = ( n_n482  &  wire16  &  n_n528 ) | ( n_n482  &  wire16  &  n_n520 ) ;
 assign _24973 = ( n_n4400 ) | ( n_n4407 ) | ( n_n4402 ) | ( _24968 ) ;
 assign _24974 = ( wire328 ) | ( wire79 ) | ( wire13070 ) ;
 assign _24978 = ( wire22  &  n_n536  &  n_n500 ) | ( n_n536  &  wire11  &  n_n500 ) ;
 assign _24983 = ( n_n4365 ) | ( n_n4368 ) | ( wire13055 ) | ( _24978 ) ;
 assign _25017 = ( n_n4345 ) | ( wire124 ) | ( wire675 ) | ( wire13085 ) ;
 assign _25018 = ( wire13066 ) | ( wire13063 ) | ( _24983 ) ;
 assign _25047 = ( n_n522  &  wire10  &  n_n509 ) | ( n_n524  &  wire10  &  n_n509 ) ;
 assign _25048 = ( wire15  &  n_n390  &  n_n509 ) | ( n_n390  &  n_n509  &  wire20 ) ;
 assign _25076 = ( n_n473  &  wire22  &  n_n455 ) | ( n_n473  &  n_n455  &  wire23 ) ;
 assign _25084 = ( wire455 ) | ( wire82 ) | ( wire13128 ) | ( _1018 ) ;
 assign _25085 = ( n_n3861 ) | ( wire13124 ) | ( wire13117 ) | ( wire13120 ) ;
 assign _25094 = ( wire25  &  n_n535  &  n_n260 ) | ( wire15  &  n_n535  &  n_n260 ) ;
 assign _25187 = ( wire12601 ) | ( wire139 ) | ( wire310 ) ;
 assign _25250 = ( n_n518  &  wire21  &  n_n390 ) | ( n_n518  &  wire11  &  n_n390 ) ;
 assign _25251 = ( n_n526  &  n_n518  &  wire10 ) | ( n_n522  &  n_n518  &  wire10 ) ;
 assign _25252 = ( n_n4593 ) | ( n_n524  &  n_n518  &  wire10 ) ;
 assign _25280 = ( n_n4635 ) | ( n_n4620 ) | ( wire13461 ) ;
 assign _25314 = ( n_n4533 ) | ( n_n4536 ) | ( wire379 ) | ( wire13479 ) ;
 assign _25315 = ( wire13468 ) | ( wire13465 ) | ( _25280 ) ;
 assign _25322 = ( n_n4389 ) | ( n_n526  &  n_n491  &  wire16 ) ;
 assign _25336 = ( n_n4397 ) | ( n_n4398 ) | ( wire13534 ) ;
 assign _25337 = ( n_n4411 ) | ( n_n4412 ) | ( wire79 ) | ( wire13529 ) ;
 assign _25342 = ( wire16  &  n_n518  &  n_n532 ) | ( wire16  &  n_n518  &  n_n534 ) ;
 assign _25369 = ( n_n522  &  wire16  &  n_n500 ) | ( wire16  &  n_n520  &  n_n500 ) ;
 assign _25381 = ( n_n4365 ) | ( wire13055 ) | ( wire13542 ) | ( wire13543 ) ;
 assign _25382 = ( n_n2446 ) | ( n_n4279 ) | ( wire13520 ) | ( wire13516 ) ;
 assign _25401 = ( wire15  &  n_n455  &  n_n509 ) | ( n_n455  &  wire24  &  n_n509 ) ;
 assign _25431 = ( wire22  &  n_n455  &  n_n500 ) | ( n_n455  &  wire24  &  n_n500 ) ;
 assign _25432 = ( n_n522  &  wire13  &  n_n500 ) | ( wire13  &  n_n500  &  n_n530 ) ;
 assign _25436 = ( n_n491  &  wire13  &  n_n532 ) | ( n_n491  &  wire13  &  n_n530 ) ;
 assign _25438 = ( n_n4505 ) | ( _25431 ) | ( _25432 ) | ( _25436 ) ;
 assign _25451 = ( n_n4982 ) | ( n_n4981 ) | ( wire57 ) | ( wire13417 ) ;
 assign _25538 = ( wire13163 ) | ( wire13162 ) ;
 assign _25555 = ( wire102 ) | ( wire245 ) | ( wire277 ) | ( wire176 ) ;
 assign _25558 = ( n_n4843 ) | ( wire13177 ) | ( wire13178 ) | ( _904 ) ;
 assign _25595 = ( wire131 ) | ( wire13182 ) | ( wire13185 ) ;
 assign _25596 = ( n_n4065 ) | ( wire13166 ) | ( n_n3996 ) | ( _25538 ) ;
 assign _25597 = ( wire13181 ) | ( wire13187 ) | ( _25558 ) | ( _25595 ) ;
 assign _25598 = ( wire134 ) | ( n_n4980 ) | ( wire13422 ) | ( _25451 ) ;
 assign _25613 = ( wire24  &  n_n535  &  n_n195 ) | ( n_n535  &  n_n195  &  wire20 ) ;
 assign _25616 = ( wire228 ) | ( wire13217 ) | ( wire13218 ) ;
 assign _25630 = ( n_n4869 ) | ( wire17  &  n_n500  &  n_n530 ) ;
 assign _25638 = ( wire25  &  n_n464  &  n_n260 ) | ( n_n464  &  wire11  &  n_n260 ) ;
 assign _25639 = ( n_n464  &  n_n532  &  wire17 ) | ( n_n464  &  n_n534  &  wire17 ) ;
 assign _25642 = ( n_n4926 ) | ( n_n473  &  wire15  &  n_n260 ) ;
 assign _25663 = ( n_n526  &  n_n518  &  wire14 ) | ( n_n518  &  wire14  &  n_n528 ) ;
 assign _25671 = ( wire13246 ) | ( n_n534  &  n_n509  &  wire14 ) ;
 assign _25724 = ( wire109 ) | ( n_n4752 ) | ( wire13272 ) | ( wire13274 ) ;
 assign _25725 = ( wire13270 ) | ( wire445 ) | ( wire13265 ) | ( wire13268 ) ;
 assign _25791 = ( n_n518  &  wire21  &  n_n130 ) | ( n_n518  &  wire20  &  n_n130 ) ;
 assign _25808 = ( wire19  &  n_n534  &  n_n500 ) | ( wire19  &  n_n528  &  n_n500 ) ;
 assign _25813 = ( n_n5252 ) | ( n_n5261 ) | ( n_n5259 ) | ( _25808 ) ;
 assign _25815 = ( wire25  &  n_n65  &  n_n509 ) | ( n_n65  &  wire22  &  n_n509 ) ;
 assign _25818 = ( n_n5239 ) | ( n_n5245 ) | ( n_n5242 ) | ( _25815 ) ;
 assign _25825 = ( wire13347 ) | ( wire203 ) | ( wire205 ) ;
 assign _25826 = ( wire13338 ) | ( wire13342 ) | ( _25813 ) | ( _25818 ) ;
 assign _25832 = ( wire13350 ) | ( n_n65  &  wire11  &  n_n535 ) ;
 assign _25847 = ( n_n5303 ) | ( n_n5309 ) | ( n_n5304 ) | ( _22502 ) ;
 assign _25860 = ( n_n5279 ) | ( n_n5280 ) | ( wire333 ) | ( wire13334 ) ;
 assign _25862 = ( wire13365 ) | ( n_n1530 ) | ( wire13361 ) | ( _25832 ) ;
 assign _25892 = ( n_n4540 ) | ( n_n524  &  wire13  &  n_n500 ) ;
 assign _25931 = ( n_n5112 ) | ( n_n5123 ) | ( wire13576 ) ;
 assign _25940 = ( wire25  &  n_n65  &  n_n482 ) | ( n_n65  &  n_n482  &  wire22 ) ;
 assign _25945 = ( n_n5333 ) | ( n_n5312 ) | ( n_n5298 ) | ( _25940 ) ;
 assign _25967 = ( n_n4362 ) | ( n_n4312 ) | ( wire13674 ) ;
 assign _25970 = ( wire25  &  n_n518  &  n_n455 ) | ( wire25  &  n_n455  &  n_n509 ) ;
 assign _25975 = ( n_n4413 ) | ( n_n4470 ) | ( wire13673 ) | ( _25970 ) ;
 assign _25978 = ( wire13662 ) | ( wire13663 ) | ( wire13666 ) | ( _25892 ) ;
 assign _25980 = ( wire13572 ) | ( n_n3920 ) | ( wire13683 ) | ( _25978 ) ;
 assign _26007 = ( n_n5171 ) | ( n_n5174 ) | ( wire14036 ) ;
 assign _26036 = ( wire22  &  n_n464  &  n_n130 ) | ( n_n464  &  n_n130  &  wire23 ) ;
 assign _26043 = ( wire14040 ) | ( wire14055 ) | ( wire14056 ) | ( _26007 ) ;
 assign _26064 = ( n_n5288 ) | ( wire13971 ) | ( wire13972 ) | ( _778 ) ;
 assign _26108 = ( n_n65  &  wire11  &  n_n509 ) | ( n_n65  &  n_n509  &  wire23 ) ;
 assign _26110 = ( wire384 ) | ( wire446 ) | ( wire181 ) | ( wire434 ) ;
 assign _26122 = ( n_n526  &  n_n491  &  wire18 ) | ( n_n491  &  n_n534  &  wire18 ) ;
 assign _26133 = ( n_n5005 ) | ( n_n5010 ) | ( wire14018 ) | ( wire14021 ) ;
 assign _26177 = ( wire13975 ) | ( wire14023 ) | ( _26064 ) | ( _26133 ) ;
 assign _26195 = ( wire118 ) | ( wire309 ) | ( wire14078 ) ;
 assign _26246 = ( n_n482  &  wire21  &  n_n536 ) | ( n_n482  &  n_n536  &  wire11 ) ;
 assign _26247 = ( n_n482  &  n_n526  &  wire16 ) | ( n_n482  &  wire16  &  n_n530 ) ;
 assign _26248 = ( n_n4404 ) | ( n_n482  &  n_n536  &  wire23 ) ;
 assign _26253 = ( n_n4408 ) | ( n_n473  &  n_n536  &  wire11 ) ;
 assign _26270 = ( wire15  &  n_n536  &  n_n500 ) | ( n_n536  &  wire23  &  n_n500 ) ;
 assign _26291 = ( n_n4335 ) | ( n_n4324 ) | ( n_n4329 ) | ( _25342 ) ;
 assign _26294 = ( n_n4319 ) | ( n_n526  &  wire16  &  n_n535 ) ;
 assign _26299 = ( n_n4338 ) | ( n_n4337 ) | ( wire156 ) | ( wire14192 ) ;
 assign _26304 = ( n_n4460 ) | ( wire25  &  n_n518  &  n_n455 ) ;
 assign _26306 = ( n_n455  &  wire24  &  n_n509 ) | ( n_n455  &  wire24  &  n_n500 ) ;
 assign _26307 = ( wire13  &  n_n509  &  n_n530 ) | ( wire13  &  n_n500  &  n_n530 ) ;
 assign _26324 = ( wire14133 ) | ( wire22  &  n_n455  &  n_n535 ) ;
 assign _26339 = ( n_n522  &  wire13  &  n_n500 ) | ( n_n524  &  wire13  &  n_n500 ) ;
 assign _26353 = ( n_n4247 ) | ( wire170 ) | ( wire14205 ) | ( _932 ) ;
 assign _26354 = ( wire470 ) | ( wire14144 ) | ( wire14148 ) | ( _26324 ) ;
 assign _26367 = ( n_n522  &  wire17  &  n_n500 ) | ( n_n524  &  wire17  &  n_n500 ) ;
 assign _26379 = ( wire13215 ) | ( n_n535  &  n_n195  &  wire20 ) ;
 assign _26416 = ( n_n4919 ) | ( wire13870 ) | ( wire13874 ) | ( _690 ) ;
 assign _26417 = ( wire13844 ) | ( wire13836 ) | ( wire13841 ) | ( _26379 ) ;
 assign _26451 = ( n_n4711 ) | ( n_n4721 ) | ( _670 ) | ( _22059 ) ;
 assign _26476 = ( wire25  &  n_n491  &  n_n325 ) | ( wire15  &  n_n491  &  n_n325 ) ;
 assign _26486 = ( wire11769 ) | ( n_n522  &  wire17  &  n_n535 ) ;
 assign _26498 = ( wire102 ) | ( n_n522  &  n_n518  &  wire17 ) ;
 assign _26499 = ( n_n4856 ) | ( n_n4850 ) | ( wire13815 ) | ( wire13816 ) ;
 assign _26500 = ( wire40 ) | ( wire245 ) | ( wire13813 ) ;
 assign _26515 = ( n_n4795 ) | ( wire158 ) | ( wire13798 ) | ( wire13800 ) ;
 assign _26519 = ( wire13796 ) | ( wire13797 ) | ( wire14213 ) ;
 assign _26573 = ( wire25  &  n_n491  &  n_n390 ) | ( n_n491  &  wire24  &  n_n390 ) ;
 assign _26577 = ( n_n4629 ) | ( n_n4583 ) | ( n_n4630 ) | ( _26573 ) ;
 assign _26585 = ( wire13760 ) | ( n_n4662 ) | ( n_n4683 ) | ( wire13756 ) ;
 assign _26606 = ( n_n4908 ) | ( n_n491  &  wire24  &  n_n260 ) ;
 assign _26631 = ( wire14222 ) | ( wire14065 ) | ( wire14066 ) | ( wire14068 ) ;
 assign _26646 = ( n_n491  &  n_n524  &  wire10 ) | ( n_n491  &  wire10  &  n_n532 ) ;
 assign _26648 = ( wire140 ) | ( wire14398 ) | ( wire431 ) ;
 assign _26776 = ( wire11520 ) | ( wire13  &  n_n535  &  n_n520 ) ;
 assign _26794 = ( wire14523 ) | ( wire13  &  n_n528  &  n_n535 ) ;
 assign _26795 = ( n_n4442 ) | ( n_n4437 ) | ( wire14524 ) | ( wire14526 ) ;
 assign _26796 = ( wire98 ) | ( wire215 ) | ( wire14522 ) ;
 assign _26834 = ( n_n482  &  wire21  &  n_n195 ) | ( n_n482  &  wire11  &  n_n195 ) ;
 assign _26840 = ( n_n5063 ) | ( n_n473  &  n_n524  &  wire18 ) ;
 assign _26875 = ( wire14655 ) | ( n_n4152 ) | ( wire14652 ) | ( _26840 ) ;
 assign _26878 = ( n_n524  &  wire17  &  n_n535 ) | ( n_n528  &  wire17  &  n_n535 ) ;
 assign _26879 = ( wire15  &  n_n535  &  n_n260 ) | ( wire22  &  n_n535  &  n_n260 ) ;
 assign _26880 = ( n_n4832 ) | ( n_n535  &  n_n260  &  wire20 ) ;
 assign _26883 = ( n_n526  &  n_n464  &  wire14 ) | ( n_n464  &  wire14  &  n_n530 ) ;
 assign _26907 = ( n_n4786 ) | ( n_n4204 ) | ( wire447 ) | ( _564 ) ;
 assign _26926 = ( wire295 ) | ( wire375 ) | ( wire324 ) | ( wire14691 ) ;
 assign _26929 = ( n_n4853 ) | ( n_n2727 ) | ( wire14726 ) | ( _560 ) ;
 assign _26931 = ( n_n3645 ) | ( wire14723 ) | ( wire14730 ) | ( _26907 ) ;
 assign _26964 = ( n_n4885 ) | ( n_n491  &  n_n532  &  wire17 ) ;
 assign _27049 = ( n_n4579 ) | ( n_n526  &  wire10  &  n_n509 ) ;
 assign _27085 = ( n_n4408 ) | ( n_n4406 ) | ( wire14334 ) | ( wire14338 ) ;
 assign _27086 = ( wire14307 ) | ( wire14308 ) | ( wire14311 ) | ( _27049 ) ;
 assign _27110 = ( wire12883 ) | ( wire15  &  n_n130  &  n_n500 ) ;
 assign _27137 = ( wire33 ) | ( wire14631 ) | ( wire14635 ) ;
 assign _27138 = ( wire14614 ) | ( n_n3772 ) | ( wire14610 ) | ( _27110 ) ;
 assign _27142 = ( n_n5278 ) | ( n_n65  &  n_n491  &  wire24 ) ;
 assign _27156 = ( wire409 ) | ( wire205 ) | ( wire14550 ) ;
 assign _27192 = ( n_n522  &  n_n518  &  wire14 ) | ( n_n524  &  n_n518  &  wire14 ) ;
 assign _27197 = ( n_n4715 ) | ( n_n4716 ) | ( n_n4723 ) | ( _27192 ) ;
 assign _27206 = ( wire14347 ) | ( wire14355 ) | ( wire14356 ) | ( _27197 ) ;
 assign _27223 = ( wire72 ) | ( n_n482  &  wire22  &  n_n390 ) ;
 assign _27224 = ( n_n4664 ) | ( n_n4669 ) | ( wire14365 ) | ( wire14367 ) ;
 assign _27225 = ( n_n4674 ) | ( n_n4673 ) | ( wire14362 ) | ( wire80 ) ;
 assign _27243 = ( n_n4754 ) | ( n_n4749 ) | ( wire109 ) | ( wire14385 ) ;
 assign _27245 = ( wire14350 ) | ( wire14351 ) | ( wire14774 ) | ( _27206 ) ;
 assign _27260 = ( n_n4439 ) | ( n_n455  &  wire24  &  n_n535 ) ;
 assign _27356 = ( wire25  &  n_n536  &  n_n500 ) | ( n_n536  &  wire24  &  n_n500 ) ;
 assign _27364 = ( wire25  &  n_n482  &  n_n536 ) | ( n_n482  &  n_n536  &  wire24 ) ;
 assign _27368 = ( n_n4388 ) | ( n_n4392 ) | ( n_n4394 ) | ( _27364 ) ;
 assign _27369 = ( wire15029 ) | ( wire15028 ) ;
 assign _27388 = ( wire14519 ) | ( n_n464  &  n_n536  &  wire24 ) ;
 assign _27389 = ( n_n4432 ) | ( n_n4431 ) | ( wire37 ) | ( wire15052 ) ;
 assign _27390 = ( wire15044 ) | ( n_n4421 ) | ( wire215 ) | ( wire15043 ) ;
 assign _27424 = ( wire335 ) | ( n_n5115 ) | ( wire11914 ) ;
 assign _27425 = ( n_n5100 ) | ( n_n5103 ) | ( wire15245 ) | ( wire15243 ) ;
 assign _27427 = ( n_n5065 ) | ( n_n524  &  n_n535  &  wire12 ) ;
 assign _27452 = ( wire297 ) | ( wire394 ) | ( wire15261 ) ;
 assign _27453 = ( n_n4152 ) | ( wire90 ) | ( wire15235 ) | ( _27427 ) ;
 assign _27469 = ( n_n5288 ) | ( n_n5286 ) | ( wire218 ) ;
 assign _27470 = ( wire115 ) | ( n_n5315 ) | ( wire13557 ) | ( wire15188 ) ;
 assign _27472 = ( n_n65  &  n_n482  &  wire22 ) | ( n_n65  &  n_n482  &  wire11 ) ;
 assign _27475 = ( n_n5305 ) | ( n_n5302 ) | ( n_n5298 ) | ( _27472 ) ;
 assign _27476 = ( n_n65  &  n_n491  &  wire22 ) | ( n_n65  &  n_n491  &  wire11 ) ;
 assign _27478 = ( n_n5274 ) | ( n_n5271 ) | ( n_n5280 ) | ( _27476 ) ;
 assign _27489 = ( n_n5262 ) | ( n_n5259 ) | ( wire334 ) | ( wire15180 ) ;
 assign _27498 = ( wire15195 ) | ( wire15198 ) | ( _27475 ) | ( _27478 ) ;
 assign _27515 = ( wire254 ) | ( wire288 ) | ( wire407 ) | ( wire15280 ) ;
 assign _27519 = ( n_n65  &  wire21  &  n_n535 ) | ( n_n65  &  wire11  &  n_n535 ) ;
 assign _27547 = ( wire211 ) | ( wire15289 ) | ( wire15292 ) | ( wire15294 ) ;
 assign _27548 = ( wire15206 ) | ( wire15184 ) | ( wire15185 ) | ( _27498 ) ;
 assign _27572 = ( n_n4797 ) | ( n_n473  &  n_n524  &  wire14 ) ;
 assign _27574 = ( n_n482  &  n_n526  &  wire14 ) | ( n_n526  &  n_n464  &  wire14 ) ;
 assign _27575 = ( n_n482  &  wire11  &  n_n325 ) | ( n_n464  &  wire11  &  n_n325 ) ;
 assign _27581 = ( wire131 ) | ( wire313 ) | ( _27574 ) | ( _27575 ) ;
 assign _27582 = ( wire14917 ) | ( wire14918 ) | ( _27572 ) | ( _27581 ) ;
 assign _27584 = ( wire12179 ) | ( wire25  &  n_n491  &  n_n260 ) ;
 assign _27589 = ( n_n522  &  wire17  &  n_n500 ) | ( n_n524  &  wire17  &  n_n500 ) ;
 assign _27591 = ( n_n509  &  n_n528  &  wire17 ) | ( n_n509  &  wire17  &  n_n520 ) ;
 assign _27623 = ( n_n4918 ) | ( n_n4917 ) | ( wire14956 ) | ( wire14957 ) ;
 assign _27671 = ( n_n4717 ) | ( n_n4716 ) | ( _362 ) | ( _25663 ) ;
 assign _27702 = ( n_n4778 ) | ( wire15020 ) | ( wire15021 ) | ( _356 ) ;
 assign _27703 = ( wire15006 ) | ( n_n4222 ) | ( wire14999 ) | ( wire15002 ) ;
 assign _27731 = ( n_n4886 ) | ( wire22  &  n_n509  &  n_n260 ) ;
 assign _27741 = ( n_n526  &  n_n518  &  wire12 ) | ( n_n518  &  n_n532  &  wire12 ) ;
 assign _27832 = ( n_n491  &  n_n524  &  wire14 ) | ( n_n491  &  wire14  &  n_n530 ) ;
 assign _27833 = ( wire15  &  n_n491  &  n_n325 ) | ( n_n491  &  wire24  &  n_n325 ) ;
 assign _27835 = ( wire15763 ) | ( _27832 ) | ( _27833 ) ;
 assign _27854 = ( n_n4721 ) | ( n_n4716 ) | ( n_n4713 ) | ( _22059 ) ;
 assign _27859 = ( n_n4749 ) | ( n_n509  &  n_n325  &  wire23 ) ;
 assign _27861 = ( wire244 ) | ( n_n4725 ) | ( n_n4726 ) | ( wire15747 ) ;
 assign _27868 = ( n_n473  &  n_n534  &  wire17 ) | ( n_n473  &  n_n528  &  wire17 ) ;
 assign _27885 = ( n_n4996 ) | ( n_n4999 ) | ( wire15707 ) ;
 assign _27896 = ( wire13217 ) | ( wire228 ) ;
 assign _27897 = ( n_n4956 ) | ( n_n4965 ) | ( wire13218 ) | ( wire15723 ) ;
 assign _27906 = ( wire15712 ) | ( _27885 ) | ( _27896 ) | ( _27897 ) ;
 assign _27910 = ( n_n4884 ) | ( wire11  &  n_n260  &  n_n500 ) ;
 assign _27917 = ( wire25  &  n_n491  &  n_n260 ) | ( n_n491  &  n_n260  &  wire23 ) ;
 assign _27951 = ( n_n3450 ) | ( wire15802 ) | ( wire15805 ) | ( _27910 ) ;
 assign _27952 = ( wire15743 ) | ( wire15738 ) | ( wire15739 ) | ( wire15741 ) ;
 assign _27996 = ( n_n5230 ) | ( n_n5168 ) | ( wire107 ) | ( wire15375 ) ;
 assign _28000 = ( n_n4515 ) | ( n_n482  &  wire13  &  n_n534 ) ;
 assign _28058 = ( wire15328 ) | ( n_n4609 ) | ( wire401 ) | ( wire15326 ) ;
 assign _28071 = ( wire25  &  n_n509  &  n_n325 ) | ( wire24  &  n_n509  &  n_n325 ) ;
 assign _28106 = ( n_n390  &  n_n535  &  wire20 ) | ( n_n390  &  n_n535  &  wire23 ) ;
 assign _28114 = ( n_n4663 ) | ( wire225 ) | ( wire11856 ) ;
 assign _28116 = ( wire309 ) | ( wire140 ) | ( wire391 ) | ( wire157 ) ;
 assign _28124 = ( wire15490 ) | ( wire190 ) ;
 assign _28137 = ( wire15469 ) | ( wire15493 ) | ( _28114 ) | ( _28124 ) ;
 assign _28144 = ( n_n526  &  wire16  &  n_n509 ) | ( wire16  &  n_n509  &  n_n528 ) ;
 assign _28151 = ( wire67 ) | ( n_n4349 ) | ( wire15517 ) | ( _28144 ) ;
 assign _28172 = ( wire25  &  n_n482  &  n_n536 ) | ( n_n482  &  n_n536  &  wire11 ) ;
 assign _28175 = ( n_n4388 ) | ( n_n4392 ) | ( n_n4396 ) | ( _28172 ) ;
 assign _28185 = ( n_n4374 ) | ( n_n4369 ) | ( n_n4373 ) | ( wire15546 ) ;
 assign _28238 = ( n_n5032 ) | ( n_n5028 ) | ( wire265 ) ;
 assign _28239 = ( n_n5039 ) | ( wire97 ) | ( wire13983 ) | ( wire15597 ) ;
 assign _28262 = ( n_n5179 ) | ( n_n5173 ) | ( wire44 ) | ( wire15591 ) ;
 assign _28268 = ( n_n5183 ) | ( n_n5188 ) | ( wire15557 ) ;
 assign _28280 = ( n_n65  &  wire21  &  n_n509 ) | ( n_n65  &  n_n509  &  wire23 ) ;
 assign _28289 = ( wire15562 ) | ( wire15575 ) | ( wire15576 ) | ( _28268 ) ;
 assign _28301 = ( n_n5295 ) | ( wire15666 ) | ( wire15667 ) | ( _230 ) ;
 assign _28305 = ( n_n5281 ) | ( wire19  &  n_n491  &  n_n534 ) ;
 assign _28312 = ( wire25  &  n_n65  &  n_n464 ) | ( n_n65  &  n_n464  &  wire24 ) ;
 assign _28313 = ( wire19  &  n_n464  &  n_n528 ) | ( wire19  &  n_n464  &  n_n530 ) ;
 assign _28320 = ( n_n2937 ) | ( wire15593 ) | ( _28262 ) | ( _28301 ) ;
 assign _28341 = ( n_n4975 ) | ( n_n5000 ) | ( wire299 ) ;
 assign _28352 = ( wire24  &  n_n535  &  n_n195 ) | ( n_n535  &  n_n195  &  wire20 ) ;
 assign _28355 = ( n_n526  &  n_n464  &  wire17 ) | ( n_n522  &  n_n464  &  wire17 ) ;
 assign _28357 = ( wire25  &  n_n518  &  n_n195 ) | ( wire25  &  n_n535  &  n_n195 ) ;
 assign _28359 = ( wire317 ) | ( wire772 ) | ( _220 ) | ( _28357 ) ;
 assign _28361 = ( wire13215 ) | ( wire13216 ) | ( wire16175 ) | ( _28352 ) ;
 assign _28362 = ( wire16158 ) | ( wire16155 ) | ( _28341 ) ;
 assign _28370 = ( n_n526  &  n_n464  &  wire14 ) | ( n_n524  &  n_n464  &  wire14 ) ;
 assign _28382 = ( n_n522  &  wire17  &  n_n535 ) | ( wire17  &  n_n535  &  n_n520 ) ;
 assign _28406 = ( n_n4886 ) | ( n_n491  &  wire24  &  n_n260 ) ;
 assign _28412 = ( wire25  &  n_n491  &  n_n325 ) | ( wire15  &  n_n491  &  n_n325 ) ;
 assign _28413 = ( n_n325  &  wire20  &  n_n500 ) | ( n_n325  &  wire23  &  n_n500 ) ;
 assign _28416 = ( n_n4764 ) | ( n_n4763 ) | ( n_n4762 ) | ( _28412 ) ;
 assign _28422 = ( n_n4791 ) | ( n_n4792 ) | ( wire380 ) | ( wire16229 ) ;
 assign _28424 = ( n_n522  &  n_n518  &  wire14 ) | ( n_n524  &  n_n518  &  wire14 ) ;
 assign _28427 = ( n_n4718 ) | ( n_n4717 ) | ( n_n4723 ) | ( _28424 ) ;
 assign _28441 = ( n_n4709 ) | ( n_n4708 ) | ( _204 ) | ( _206 ) ;
 assign _28496 = ( n_n5131 ) | ( n_n5127 ) | ( wire15875 ) ;
 assign _28538 = ( wire15830 ) | ( wire15829 ) ;
 assign _28546 = ( n_n4725 ) | ( wire14  &  n_n535  &  n_n530 ) ;
 assign _28573 = ( n_n482  &  wire19  &  n_n532 ) | ( n_n482  &  wire19  &  n_n530 ) ;
 assign _28574 = ( n_n65  &  wire15  &  n_n482 ) | ( n_n65  &  n_n482  &  wire22 ) ;
 assign _28575 = ( n_n482  &  wire19  &  n_n524 ) | ( n_n482  &  wire19  &  n_n528 ) ;
 assign _28577 = ( n_n5296 ) | ( n_n5299 ) | ( n_n5289 ) | ( _28573 ) ;
 assign _28581 = ( wire203 ) | ( wire334 ) ;
 assign _28589 = ( wire218 ) | ( wire11946 ) | ( wire16293 ) | ( _172 ) ;
 assign _28605 = ( wire16300 ) | ( wire16305 ) | ( _28577 ) | ( _28581 ) ;
 assign _28607 = ( n_n5082 ) | ( n_n464  &  n_n195  &  wire23 ) ;
 assign _28618 = ( n_n5067 ) | ( n_n464  &  n_n534  &  wire18 ) ;
 assign _28636 = ( n_n5130 ) | ( n_n5129 ) | ( wire422 ) ;
 assign _28637 = ( n_n5112 ) | ( n_n5110 ) | ( wire15968 ) | ( wire15964 ) ;
 assign _28642 = ( n_n5045 ) | ( n_n473  &  wire15  &  n_n195 ) ;
 assign _28665 = ( wire347 ) | ( wire65 ) ;
 assign _28666 = ( wire15  &  n_n455  &  n_n509 ) | ( n_n455  &  wire24  &  n_n509 ) ;
 assign _28668 = ( wire14438 ) | ( n_n522  &  wire13  &  n_n509 ) ;
 assign _28669 = ( n_n4476 ) | ( wire184 ) | ( _144 ) | ( _28666 ) ;
 assign _28677 = ( wire22  &  n_n518  &  n_n455 ) | ( wire22  &  n_n455  &  n_n535 ) ;
 assign _28704 = ( wire15995 ) | ( _28665 ) | ( _28668 ) | ( _28669 ) ;
 assign _28709 = ( n_n526  &  wire10  &  n_n509 ) | ( n_n522  &  wire10  &  n_n509 ) ;
 assign _28710 = ( wire15  &  n_n390  &  n_n509 ) | ( n_n390  &  n_n509  &  wire20 ) ;
 assign _28731 = ( n_n491  &  wire11  &  n_n390 ) | ( n_n491  &  wire24  &  n_n390 ) ;
 assign _28734 = ( n_n4634 ) | ( wire26 ) | ( n_n4633 ) ;
 assign _28735 = ( wire309 ) | ( n_n4642 ) | ( wire16059 ) | ( wire16057 ) ;
 assign _28741 = ( n_n4574 ) | ( wire15  &  n_n390  &  n_n535 ) ;
 assign _28749 = ( n_n4557 ) | ( wire430 ) | ( n_n4558 ) ;
 assign _28750 = ( n_n4582 ) | ( n_n4581 ) | ( wire276 ) | ( wire16031 ) ;
 assign _28753 = ( wire15  &  n_n482  &  n_n536 ) | ( n_n482  &  n_n536  &  wire11 ) ;
 assign _28757 = ( n_n4391 ) | ( n_n4398 ) | ( n_n4396 ) | ( _28753 ) ;
 assign _28767 = ( n_n4421 ) | ( wire215 ) | ( wire16094 ) | ( wire16093 ) ;
 assign _28771 = ( wire12569 ) | ( wire21  &  n_n536  &  n_n535 ) ;
 assign _28786 = ( wire13055 ) | ( wire15  &  n_n536  &  n_n500 ) ;
 assign _28787 = ( n_n4368 ) | ( wire16088 ) | ( _120 ) | ( _24978 ) ;
 assign _28790 = ( wire25  &  n_n536  &  n_n500 ) | ( n_n536  &  wire24  &  n_n500 ) ;
 assign _28794 = ( n_n4386 ) | ( wire12447 ) | ( wire14460 ) | ( wire16091 ) ;
 assign _28812 = ( wire385 ) | ( n_n5215 ) | ( wire16272 ) | ( wire16270 ) ;
 assign _28817 = ( wire453 ) | ( n_n464  &  n_n532  &  wire12 ) ;
 assign _28838 = ( wire288 ) | ( wire16282 ) | ( wire16286 ) ;
 assign _28839 = ( wire16263 ) | ( n_n2291 ) | ( wire16259 ) | ( _28817 ) ;
 assign _28844 = ( wire25  &  n_n65  &  n_n509 ) | ( n_n65  &  wire15  &  n_n509 ) ;
 assign _28847 = ( n_n5238 ) | ( n_n5244 ) | ( n_n5242 ) | ( _28844 ) ;
 assign _28857 = ( wire16686 ) | ( wire16691 ) | ( wire16692 ) | ( _28847 ) ;
 assign _28879 = ( wire358 ) | ( wire125 ) | ( wire44 ) | ( wire332 ) ;
 assign _28882 = ( wire168 ) | ( wire16698 ) | ( wire16702 ) ;
 assign _28884 = ( wire16696 ) | ( wire16704 ) | ( _28857 ) | ( _28882 ) ;
 assign _28885 = ( n_n473  &  wire22  &  n_n195 ) | ( n_n473  &  wire21  &  n_n195 ) ;
 assign _28888 = ( n_n5060 ) | ( n_n5055 ) | ( n_n5058 ) | ( _28885 ) ;
 assign _28895 = ( n_n5024 ) | ( wire14661 ) | ( wire253 ) | ( wire13400 ) ;
 assign _28900 = ( wire25  &  n_n535  &  n_n130 ) | ( wire11  &  n_n535  &  n_n130 ) ;
 assign _28912 = ( n_n518  &  wire21  &  n_n130 ) | ( n_n518  &  wire20  &  n_n130 ) ;
 assign _28923 = ( n_n65  &  n_n482  &  wire11 ) | ( n_n65  &  n_n482  &  wire24 ) ;
 assign _28927 = ( n_n5294 ) | ( n_n5299 ) | ( n_n5292 ) | ( _28923 ) ;
 assign _28931 = ( wire14542 ) | ( n_n65  &  n_n491  &  wire20 ) ;
 assign _28934 = ( wire16753 ) | ( wire16754 ) | ( wire16749 ) | ( _28927 ) ;
 assign _28935 = ( n_n5302 ) | ( n_n473  &  wire19  &  n_n532 ) ;
 assign _28949 = ( wire117 ) | ( wire12969 ) | ( wire16761 ) | ( _28935 ) ;
 assign _28951 = ( wire16745 ) | ( n_n2214 ) | ( wire16742 ) | ( _28895 ) ;
 assign _28952 = ( wire16763 ) | ( wire16682 ) | ( wire16683 ) | ( _28884 ) ;
 assign _29002 = ( n_n482  &  wire22  &  n_n536 ) | ( n_n482  &  n_n536  &  wire24 ) ;
 assign _29003 = ( n_n482  &  wire21  &  n_n536 ) | ( n_n482  &  n_n536  &  wire11 ) ;
 assign _29004 = ( n_n482  &  wire16  &  n_n534 ) | ( n_n482  &  wire16  &  n_n530 ) ;
 assign _29006 = ( n_n4393 ) | ( n_n4398 ) | ( n_n4402 ) | ( _29002 ) ;
 assign _29007 = ( n_n4440 ) | ( n_n4434 ) | ( wire16527 ) | ( wire215 ) ;
 assign _29028 = ( n_n2435 ) | ( wire54 ) | ( wire282 ) ;
 assign _29029 = ( wire16545 ) | ( wire16537 ) | ( wire16538 ) | ( wire16544 ) ;
 assign _29041 = ( wire15  &  n_n509  &  n_n130 ) | ( wire22  &  n_n509  &  n_n130 ) ;
 assign _29050 = ( n_n4981 ) | ( n_n5005 ) | ( wire16799 ) ;
 assign _29051 = ( n_n5122 ) | ( wire16790 ) | ( wire16788 ) | ( _29041 ) ;
 assign _29082 = ( n_n518  &  n_n536  &  wire20 ) | ( n_n536  &  n_n509  &  wire20 ) ;
 assign _29086 = ( n_n4367 ) | ( n_n4374 ) | ( n_n4358 ) | ( _29082 ) ;
 assign _29091 = ( wire16770 ) | ( wire16769 ) ;
 assign _29098 = ( n_n4883 ) | ( n_n4895 ) | ( n_n4890 ) | ( _26367 ) ;
 assign _29100 = ( n_n4859 ) | ( n_n526  &  n_n509  &  wire17 ) ;
 assign _29196 = ( n_n4937 ) | ( n_n473  &  n_n260  &  wire20 ) ;
 assign _29216 = ( n_n509  &  n_n528  &  wire18 ) | ( n_n509  &  wire18  &  n_n530 ) ;
 assign _29219 = ( n_n4987 ) | ( n_n4979 ) | ( wire16438 ) | ( _29216 ) ;
 assign _29241 = ( wire16462 ) | ( wire250 ) ;
 assign _29242 = ( wire341 ) | ( wire362 ) | ( wire16461 ) ;
 assign _29247 = ( n_n4487 ) | ( n_n4478 ) | ( n_n4476 ) | ( _28666 ) ;
 assign _29258 = ( wire65 ) | ( wire66 ) | ( wire16574 ) ;
 assign _29270 = ( n_n518  &  wire21  &  n_n455 ) | ( n_n518  &  n_n455  &  wire23 ) ;
 assign _29306 = ( wire365 ) | ( n_n4591 ) | ( n_n4592 ) ;
 assign _29324 = ( n_n491  &  wire11  &  n_n390 ) | ( n_n491  &  wire24  &  n_n390 ) ;
 assign _29335 = ( wire16621 ) | ( wire16635 ) | ( wire16636 ) | ( _29306 ) ;


endmodule

