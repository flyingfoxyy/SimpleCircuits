module dalu (
	Psh2, Psh1, Psh0, Popsel3, Popsel2, Popsel1, Popsel0, Pmusel4, 
	Pmusel3, Pmusel2, Pmusel1, PinD15, PinD14, PinD13, PinD12, PinD11, PinD10, PinD9, 
	PinD8, PinD7, PinD6, PinD5, PinD4, PinD3, PinD2, PinD1, PinD0, PinC15, 
	PinC14, PinC13, PinC12, PinC11, PinC10, PinC9, PinC8, PinC7, PinC6, PinC5, 
	PinC4, PinC3, PinC2, PinC1, PinC0, PinB15, PinB14, PinB13, PinB12, PinB11, 
	PinB10, PinB9, PinB8, PinB7, PinB6, PinB5, PinB4, PinB3, PinB2, PinB1, 
	PinB0, PinA15, PinA14, PinA13, PinA12, PinA11, PinA10, PinA9, PinA8, PinA7, 
	PinA6, PinA5, PinA4, PinA3, PinA2, PinA1, PinA0, PO15, PO14, PO13, 
	PO12, PO11, PO10, PO9, PO8, PO7, PO6, PO5, PO4, PO3, 
	PO2, PO1, PO0);

input Psh2, Psh1, Psh0, Popsel3, Popsel2, Popsel1, Popsel0, Pmusel4, Pmusel3, Pmusel2, Pmusel1, PinD15, PinD14, PinD13, PinD12, PinD11, PinD10, PinD9, PinD8, PinD7, PinD6, PinD5, PinD4, PinD3, PinD2, PinD1, PinD0, PinC15, PinC14, PinC13, PinC12, PinC11, PinC10, PinC9, PinC8, PinC7, PinC6, PinC5, PinC4, PinC3, PinC2, PinC1, PinC0, PinB15, PinB14, PinB13, PinB12, PinB11, PinB10, PinB9, PinB8, PinB7, PinB6, PinB5, PinB4, PinB3, PinB2, PinB1, PinB0, PinA15, PinA14, PinA13, PinA12, PinA11, PinA10, PinA9, PinA8, PinA7, PinA6, PinA5, PinA4, PinA3, PinA2, PinA1, PinA0;

output PO15, PO14, PO13, PO12, PO11, PO10, PO9, PO8, PO7, PO6, PO5, PO4, PO3, PO2, PO1, PO0;

wire n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n18, n20, n17, n22, n25, n28, n31, n34, n35, n36, n40, n39, n41, n46, n47, n45, n44, n49, n48, n54, n53, n57, n56, n60, n59, n63, n62, n66, n65, n69, n68, n72, n71, n77, n76, n74, n79, n78, n82, n83, n84, n81, n86, n87, n88, n94, n95, n92, n93, n91, n97, n96, n98, n103, n104, n102, n101, n106, n107, n105, n110, n108, n109, n111, n116, n117, n115, n114, n119, n118, n121, n120, n122, n127, n128, n126, n125, n130, n129, n131, n132, n137, n138, n136, n135, n139, n140, n145, n146, n144, n143, n148, n149, n147, n151, n150, n152, n153, n158, n159, n157, n156, n160, n162, n161, n164, n168, n167, n171, n170, n174, n173, n177, n176, n180, n179, n183, n182, n184, n185, n187, n186, n189, n190, n188, n192, n193, n191, n194, n195, n202, n200, n199, n204, n203, n205, n208, n207, n206, n210, n211, n209, n212, n214, n215, n213, n218, n217, n220, n221, n219, n223, n222, n224, n225, n226, n231, n232, n230, n229, n233, n234, n239, n240, n237, n241, n244, n242, n245, n247, n246, n249, n248, n251, n250, n253, n254, n252, n256, n255, n257, n261, n263, n262, n265, n264, n266, n268, n267, n273, n270, n274, n277, n279, n278, n282, n283, n288, n285, n289, n293, n294, n298, n295, n300, n299, n302, n301, n303, n306, n307, n312, n309, n313, n316, n318, n317, n322, n319, n326, n323, n329, n333, n330, n335, n334, n339, n336, n340, n341, n343, n344, n345, n348, n349, n351, n353, n354, n359, n360, n363, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n389, n390, n392, n393, n394, n395, n396, n397, n399, n400, n401, n403, n406, n407, n408, n409, n410, n411, n413, n414, n415;

assign PO15 = ( (~ n1) ) ;
 assign PO14 = ( (~ n2) ) ;
 assign PO13 = ( (~ n3) ) ;
 assign PO12 = ( (~ n4) ) ;
 assign PO11 = ( (~ n5) ) ;
 assign PO10 = ( (~ n6) ) ;
 assign PO9 = ( (~ n7) ) ;
 assign PO8 = ( (~ n8) ) ;
 assign PO7 = ( (~ n9) ) ;
 assign PO6 = ( (~ n10) ) ;
 assign PO5 = ( (~ n11) ) ;
 assign PO4 = ( (~ n12) ) ;
 assign PO3 = ( (~ n13) ) ;
 assign PO2 = ( (~ n14) ) ;
 assign PO1 = ( (~ n15) ) ;
 assign PO0 = ( (~ n16) ) ;
 assign n1 = ( n184  &  n185  &  n36 ) | ( n184  &  n185  &  n120 ) ;
 assign n2 = ( n194  &  n193 ) | ( n194  &  n120 ) ;
 assign n3 = ( n205  &  n199 ) | ( n205  &  n120 ) ;
 assign n4 = ( n212  &  n96 ) | ( n212  &  n209 ) ;
 assign n5 = ( n109  &  n218 ) | ( n218  &  n217 ) | ( n218  &  (~ n344) ) ;
 assign n6 = ( n222  &  n224  &  n225 ) | ( n224  &  n225  &  (~ n354) ) ;
 assign n7 = ( n81  &  n86  &  n87 ) | ( n86  &  n87  &  (~ n354) ) ;
 assign n8 = ( n97  &  n91 ) | ( n97  &  n96 ) ;
 assign n9 = ( n110  &  n108 ) | ( n110  &  n109 ) ;
 assign n10 = ( n121  &  n114 ) | ( n121  &  n120 ) ;
 assign n11 = ( n131  &  n125 ) | ( n131  &  n120 ) ;
 assign n12 = ( n139  &  n96 ) | ( n139  &  n135 ) ;
 assign n13 = ( n152  &  n143 ) | ( n152  &  n120 ) ;
 assign n14 = ( n160  &  n96 ) | ( n160  &  n156 ) ;
 assign n15 = ( n233  &  n229 ) | ( n233  &  n96 ) ;
 assign n16 = ( n241  &  n237 ) | ( n241  &  n96 ) ;
 assign n18 = ( n164  &  n309 ) ;
 assign n20 = ( n34 ) | ( n35 ) ;
 assign n17 = ( (~ PinD12)  &  (~ PinB12) ) | ( (~ PinB12)  &  n18 ) | ( (~ PinD12)  &  n20 ) | ( n18  &  n20 ) ;
 assign n22 = ( (~ PinD9)  &  (~ PinB9) ) | ( (~ PinB9)  &  n18 ) | ( (~ PinD9)  &  n20 ) | ( n18  &  n20 ) ;
 assign n25 = ( (~ PinD14)  &  (~ PinB14) ) | ( (~ PinB14)  &  n18 ) | ( (~ PinD14)  &  n20 ) | ( n18  &  n20 ) ;
 assign n28 = ( (~ PinD10)  &  (~ PinB10) ) | ( (~ PinB10)  &  n18 ) | ( (~ PinD10)  &  n20 ) | ( n18  &  n20 ) ;
 assign n31 = ( (~ PinD11)  &  (~ PinB11) ) | ( (~ PinB11)  &  n18 ) | ( (~ PinD11)  &  n20 ) | ( n18  &  n20 ) ;
 assign n34 = ( Pmusel2  &  Pmusel1 ) | ( (~ Pmusel2)  &  (~ Pmusel1) ) ;
 assign n35 = ( Pmusel4 ) | ( (~ Pmusel3) ) ;
 assign n36 = ( (~ PinD15)  &  (~ PinB15) ) | ( (~ PinB15)  &  n18 ) | ( (~ PinD15)  &  n20 ) | ( n18  &  n20 ) ;
 assign n40 = ( (~ Psh2) ) | ( n36 ) ;
 assign n39 = ( n40  &  Psh2 ) | ( n40  &  n31 ) ;
 assign n41 = ( (~ PinD13)  &  (~ PinB13) ) | ( (~ PinB13)  &  n18 ) | ( (~ PinD13)  &  n20 ) | ( n18  &  n20 ) ;
 assign n46 = ( n22  &  n92 ) | ( n208  &  n92 ) | ( n22  &  n207 ) | ( n208  &  n207 ) ;
 assign n47 = ( n378  &  n39 ) | ( n93  &  n39 ) | ( n378  &  n353 ) | ( n93  &  n353 ) ;
 assign n45 = ( Psh2 ) | ( n351 ) ;
 assign n44 = ( n46  &  n47  &  n17 ) | ( n46  &  n47  &  n45 ) ;
 assign n49 = ( Pmusel2  &  PinC7 ) | ( (~ Pmusel2)  &  PinA7 ) | ( PinC7  &  PinA7 ) ;
 assign n48 = ( (~ Pmusel4)  &  (~ n384) ) | ( (~ Pmusel4)  &  n49  &  (~ n76) ) ;
 assign n54 = ( Pmusel2  &  PinC6 ) | ( (~ Pmusel2)  &  PinA6 ) | ( PinC6  &  PinA6 ) ;
 assign n53 = ( (~ Pmusel4)  &  (~ n386) ) | ( (~ Pmusel4)  &  n54  &  (~ n76) ) ;
 assign n57 = ( Pmusel2  &  PinC5 ) | ( (~ Pmusel2)  &  PinA5 ) | ( PinC5  &  PinA5 ) ;
 assign n56 = ( (~ Pmusel4)  &  (~ n389) ) | ( (~ Pmusel4)  &  n57  &  (~ n76) ) ;
 assign n60 = ( Pmusel2  &  PinC3 ) | ( (~ Pmusel2)  &  PinA3 ) | ( PinC3  &  PinA3 ) ;
 assign n59 = ( (~ Pmusel4)  &  (~ n394) ) | ( (~ Pmusel4)  &  n60  &  (~ n76) ) ;
 assign n63 = ( Pmusel2  &  PinC2 ) | ( (~ Pmusel2)  &  PinA2 ) | ( PinC2  &  PinA2 ) ;
 assign n62 = ( (~ Pmusel4)  &  (~ n396) ) | ( (~ Pmusel4)  &  n63  &  (~ n76) ) ;
 assign n66 = ( Pmusel2  &  PinC1 ) | ( (~ Pmusel2)  &  PinA1 ) | ( PinC1  &  PinA1 ) ;
 assign n65 = ( (~ Pmusel4)  &  (~ n409) ) | ( (~ Pmusel4)  &  n66  &  (~ n76) ) ;
 assign n69 = ( Pmusel2  &  PinC0 ) | ( (~ Pmusel2)  &  PinA0 ) | ( PinC0  &  PinA0 ) ;
 assign n68 = ( (~ Pmusel4)  &  (~ n413) ) | ( (~ Pmusel4)  &  n69  &  (~ n76) ) ;
 assign n72 = ( Pmusel2  &  PinC4 ) | ( (~ Pmusel2)  &  PinA4 ) | ( PinC4  &  PinA4 ) ;
 assign n71 = ( (~ Pmusel4)  &  (~ n392) ) | ( (~ Pmusel4)  &  n72  &  (~ n76) ) ;
 assign n77 = ( (~ PinD8)  &  (~ PinB8) ) | ( (~ PinB8)  &  n348 ) | ( (~ PinD8)  &  n349 ) | ( n348  &  n349 ) ;
 assign n76 = ( Pmusel3 ) | ( (~ Pmusel1) ) ;
 assign n74 = ( n77  &  n76 ) | ( n77  &  (~ n376) ) ;
 assign n79 = ( Pmusel2  &  PinC9 ) | ( (~ Pmusel2)  &  PinA9 ) | ( PinC9  &  PinA9 ) ;
 assign n78 = ( (~ Pmusel4)  &  (~ n377) ) | ( (~ Pmusel4)  &  (~ n76)  &  n79 ) ;
 assign n82 = ( Popsel1  &  Popsel0 ) | ( (~ Popsel1)  &  (~ Popsel0) ) ;
 assign n83 = ( (~ PinA9)  &  (~ n78)  &  n261 ) | ( n20  &  (~ n78)  &  n261 ) ;
 assign n84 = ( Popsel0 ) | ( Popsel1 ) ;
 assign n81 = ( n82  &  n44 ) | ( n83  &  n44 ) | ( n82  &  n84 ) | ( n83  &  n84 ) ;
 assign n86 = ( n109 ) | ( n242 ) | ( (~ n344) ) ;
 assign n87 = ( n44 ) | ( n120 ) ;
 assign n88 = ( (~ PinD8)  &  (~ PinB8) ) | ( (~ PinB8)  &  n18 ) | ( (~ PinD8)  &  n20 ) | ( n18  &  n20 ) ;
 assign n94 = ( n102  &  n31 ) | ( n207  &  n31 ) | ( n102  &  n45 ) | ( n207  &  n45 ) ;
 assign n95 = ( n381  &  n382  &  n28 ) | ( n381  &  n382  &  n360 ) ;
 assign n92 = ( (~ Psh2)  &  n22 ) | ( Psh2  &  n41 ) | ( n22  &  n41 ) ;
 assign n93 = ( Psh1 ) | ( (~ Psh0) ) ;
 assign n91 = ( n94  &  n95  &  n92 ) | ( n94  &  n95  &  n93 ) ;
 assign n97 = ( n383  &  n359 ) | ( n383  &  n380  &  n379 ) ;
 assign n96 = ( n84  &  n120 ) | ( n120  &  (~ n354) ) ;
 assign n98 = ( (~ PinD7)  &  (~ PinB7) ) | ( (~ PinB7)  &  n18 ) | ( (~ PinD7)  &  n20 ) | ( n18  &  n20 ) ;
 assign n103 = ( n115  &  n28 ) | ( n207  &  n28 ) | ( n115  &  n45 ) | ( n207  &  n45 ) ;
 assign n104 = ( n385  &  n382  &  n22 ) | ( n385  &  n382  &  n360 ) ;
 assign n102 = ( Psh2  &  n17 ) | ( (~ Psh2)  &  n88 ) | ( n17  &  n88 ) ;
 assign n101 = ( n103  &  n104  &  n102 ) | ( n103  &  n104  &  n93 ) ;
 assign n106 = ( n264 ) | ( n279 ) ;
 assign n107 = ( n253  &  n266 ) | ( (~ n253)  &  (~ n266) ) ;
 assign n105 = ( n106 ) | ( n107 ) ;
 assign n110 = ( n270  &  n101 ) | ( n359  &  n101 ) | ( n270  &  n96 ) | ( n359  &  n96 ) ;
 assign n108 = ( n105  &  n267 ) | ( (~ n105)  &  (~ n267) ) ;
 assign n109 = ( Popsel3 ) | ( n345 ) ;
 assign n111 = ( (~ PinD6)  &  (~ PinB6) ) | ( (~ PinB6)  &  n18 ) | ( (~ PinD6)  &  n20 ) | ( n18  &  n20 ) ;
 assign n116 = ( n126  &  n22 ) | ( n207  &  n22 ) | ( n126  &  n45 ) | ( n207  &  n45 ) ;
 assign n117 = ( n387  &  n88 ) | ( n387  &  n360 ) ;
 assign n115 = ( Psh2  &  n31 ) | ( (~ Psh2)  &  n98 ) | ( n31  &  n98 ) ;
 assign n114 = ( n116  &  n117  &  n115 ) | ( n116  &  n117  &  n93 ) ;
 assign n119 = ( (~ PinA6)  &  (~ n53)  &  n277 ) | ( n20  &  (~ n53)  &  n277 ) ;
 assign n118 = ( n82  &  n114 ) | ( n119  &  n114 ) | ( n82  &  n84 ) | ( n119  &  n84 ) ;
 assign n121 = ( n109  &  n118 ) | ( n118  &  (~ n274) ) | ( n109  &  (~ n354) ) | ( (~ n274)  &  (~ n354) ) ;
 assign n120 = ( Popsel3 ) | ( (~ Popsel2) ) | ( (~ n84) ) ;
 assign n122 = ( (~ PinD5)  &  (~ PinB5) ) | ( (~ PinB5)  &  n18 ) | ( (~ PinD5)  &  n20 ) | ( n18  &  n20 ) ;
 assign n127 = ( n136  &  n88 ) | ( n207  &  n88 ) | ( n136  &  n45 ) | ( n207  &  n45 ) ;
 assign n128 = ( n390  &  n98 ) | ( n390  &  n360 ) ;
 assign n126 = ( Psh2  &  n28 ) | ( (~ Psh2)  &  n111 ) | ( n28  &  n111 ) ;
 assign n125 = ( n127  &  n128  &  n126 ) | ( n127  &  n128  &  n93 ) ;
 assign n130 = ( (~ PinA5)  &  (~ n56)  &  n282 ) | ( n20  &  (~ n56)  &  n282 ) ;
 assign n129 = ( n82  &  n125 ) | ( n130  &  n125 ) | ( n82  &  n84 ) | ( n130  &  n84 ) ;
 assign n131 = ( n109  &  n129 ) | ( n129  &  (~ n278) ) | ( n109  &  (~ n354) ) | ( (~ n278)  &  (~ n354) ) ;
 assign n132 = ( (~ PinD4)  &  (~ PinB4) ) | ( (~ PinB4)  &  n18 ) | ( (~ PinD4)  &  n20 ) | ( n18  &  n20 ) ;
 assign n137 = ( n144  &  n98 ) | ( n207  &  n98 ) | ( n144  &  n45 ) | ( n207  &  n45 ) ;
 assign n138 = ( n393  &  n111 ) | ( n393  &  n360 ) ;
 assign n136 = ( Psh2  &  n22 ) | ( (~ Psh2)  &  n122 ) | ( n22  &  n122 ) ;
 assign n135 = ( n137  &  n138  &  n136 ) | ( n137  &  n138  &  n93 ) ;
 assign n139 = ( n283  &  n285 ) | ( n109  &  n285 ) | ( n283  &  n359 ) | ( n109  &  n359 ) ;
 assign n140 = ( (~ PinD3)  &  (~ PinB3) ) | ( (~ PinB3)  &  n18 ) | ( (~ PinD3)  &  n20 ) | ( n18  &  n20 ) ;
 assign n145 = ( n157  &  n111 ) | ( n207  &  n111 ) | ( n157  &  n45 ) | ( n207  &  n45 ) ;
 assign n146 = ( n395  &  n122 ) | ( n395  &  n360 ) ;
 assign n144 = ( Psh2  &  n88 ) | ( (~ Psh2)  &  n132 ) | ( n88  &  n132 ) ;
 assign n143 = ( n145  &  n146  &  n144 ) | ( n145  &  n146  &  n93 ) ;
 assign n148 = ( n248 ) | ( n335 ) ;
 assign n149 = ( n245  &  n253 ) | ( (~ n245)  &  (~ n253) ) ;
 assign n147 = ( n148 ) | ( n149 ) ;
 assign n151 = ( (~ PinA3)  &  (~ n59)  &  n293 ) | ( n20  &  (~ n59)  &  n293 ) ;
 assign n150 = ( n82  &  n143 ) | ( n151  &  n143 ) | ( n82  &  n84 ) | ( n151  &  n84 ) ;
 assign n152 = ( n109  &  n150 ) | ( n150  &  n289 ) | ( n109  &  (~ n354) ) | ( n289  &  (~ n354) ) ;
 assign n153 = ( (~ PinD2)  &  (~ PinB2) ) | ( (~ PinB2)  &  n18 ) | ( (~ PinD2)  &  n20 ) | ( n18  &  n20 ) ;
 assign n158 = ( n230  &  n122 ) | ( n207  &  n122 ) | ( n230  &  n45 ) | ( n207  &  n45 ) ;
 assign n159 = ( n397  &  n132 ) | ( n397  &  n360 ) ;
 assign n157 = ( Psh2  &  n98 ) | ( (~ Psh2)  &  n140 ) | ( n98  &  n140 ) ;
 assign n156 = ( n158  &  n159  &  n157 ) | ( n158  &  n159  &  n93 ) ;
 assign n160 = ( n109  &  n295 ) | ( (~ n294)  &  n295 ) | ( n109  &  n359 ) | ( (~ n294)  &  n359 ) ;
 assign n162 = ( Pmusel2  &  PinC15 ) | ( (~ Pmusel2)  &  PinA15 ) | ( PinC15  &  PinA15 ) ;
 assign n161 = ( (~ Pmusel4)  &  (~ n399) ) | ( (~ Pmusel4)  &  (~ n76)  &  n162 ) ;
 assign n164 = ( (~ Pmusel2) ) | ( (~ Pmusel1) ) | ( n35 ) ;
 assign n168 = ( Pmusel2  &  PinC14 ) | ( (~ Pmusel2)  &  PinA14 ) | ( PinC14  &  PinA14 ) ;
 assign n167 = ( (~ Pmusel4)  &  (~ n400) ) | ( (~ Pmusel4)  &  (~ n76)  &  n168 ) ;
 assign n171 = ( Pmusel2  &  PinC13 ) | ( (~ Pmusel2)  &  PinA13 ) | ( PinC13  &  PinA13 ) ;
 assign n170 = ( (~ Pmusel4)  &  (~ n401) ) | ( (~ Pmusel4)  &  (~ n76)  &  n171 ) ;
 assign n174 = ( Pmusel2  &  PinC12 ) | ( (~ Pmusel2)  &  PinA12 ) | ( PinC12  &  PinA12 ) ;
 assign n173 = ( (~ Pmusel4)  &  (~ n403) ) | ( (~ Pmusel4)  &  (~ n76)  &  n174 ) ;
 assign n177 = ( Pmusel2  &  PinC11 ) | ( (~ Pmusel2)  &  PinA11 ) | ( PinC11  &  PinA11 ) ;
 assign n176 = ( (~ Pmusel4)  &  (~ n406) ) | ( (~ Pmusel4)  &  (~ n76)  &  n177 ) ;
 assign n180 = ( Pmusel2  &  PinC10 ) | ( (~ Pmusel2)  &  PinA10 ) | ( PinC10  &  PinA10 ) ;
 assign n179 = ( (~ Pmusel4)  &  (~ n407) ) | ( (~ Pmusel4)  &  (~ n76)  &  n180 ) ;
 assign n183 = ( (~ PinA15)  &  (~ n161)  &  n306 ) | ( n20  &  (~ n161)  &  n306 ) ;
 assign n182 = ( n82  &  n36 ) | ( n183  &  n36 ) | ( n82  &  n84 ) | ( n183  &  n84 ) ;
 assign n184 = ( n182 ) | ( (~ n354) ) ;
 assign n185 = ( n109 ) | ( n189 ) | ( n301 ) | ( n190 ) ;
 assign n187 = ( (~ Psh2)  &  (~ Psh1) ) | ( Psh2  &  Psh0 ) | ( (~ Psh1)  &  Psh0 ) ;
 assign n186 = ( n187  &  n93 ) ;
 assign n189 = ( n299 ) | ( n318 ) ;
 assign n190 = ( n253  &  n303 ) | ( (~ n253)  &  (~ n303) ) ;
 assign n188 = ( n189 ) | ( n190 ) ;
 assign n192 = ( (~ PinC14)  &  (~ n167)  &  n312 ) | ( (~ n167)  &  n312  &  n309 ) ;
 assign n193 = ( n25  &  n36 ) | ( n25  &  n186 ) | ( n36  &  (~ n186) ) ;
 assign n191 = ( n82  &  n193 ) | ( n192  &  n193 ) | ( n82  &  n84 ) | ( n192  &  n84 ) ;
 assign n194 = ( n109  &  n191 ) | ( n191  &  n307 ) | ( n109  &  (~ n354) ) | ( n307  &  (~ n354) ) ;
 assign n195 = ( (~ n36)  &  (~ n353) ) | ( (~ Psh2)  &  Psh1  &  (~ n36) ) ;
 assign n202 = ( Psh1  &  n41 ) | ( n40  &  n41 ) | ( Psh1  &  (~ n186) ) | ( n40  &  (~ n186) ) ;
 assign n200 = ( Psh2 ) | ( n93 ) ;
 assign n199 = ( n25  &  (~ n195)  &  n202 ) | ( (~ n195)  &  n202  &  n200 ) ;
 assign n204 = ( (~ PinC13)  &  (~ n170)  &  n316 ) | ( (~ n170)  &  n309  &  n316 ) ;
 assign n203 = ( n82  &  n199 ) | ( n204  &  n199 ) | ( n82  &  n84 ) | ( n204  &  n84 ) ;
 assign n205 = ( n109  &  n203 ) | ( n203  &  (~ n313) ) | ( n109  &  (~ n354) ) | ( (~ n313)  &  (~ n354) ) ;
 assign n208 = ( (~ Psh2) ) | ( n351 ) ;
 assign n207 = ( Psh0 ) | ( Psh1 ) ;
 assign n206 = ( n208  &  Psh2 ) | ( n208  &  n207 ) ;
 assign n210 = ( n41  &  n25 ) | ( n200  &  n25 ) | ( n41  &  n360 ) | ( n200  &  n360 ) ;
 assign n211 = ( n36  &  n40 ) | ( n40  &  n45 ) | ( n36  &  (~ n351) ) | ( n45  &  (~ n351) ) ;
 assign n209 = ( n210  &  n211  &  n17 ) | ( n210  &  n211  &  n206 ) ;
 assign n212 = ( n109  &  n319 ) | ( (~ n317)  &  n319 ) | ( n109  &  n359 ) | ( (~ n317)  &  n359 ) ;
 assign n214 = ( n17  &  n41 ) | ( n200  &  n41 ) | ( n17  &  n360 ) | ( n200  &  n360 ) ;
 assign n215 = ( n25  &  n40 ) | ( n40  &  n45 ) | ( n25  &  (~ n351) ) | ( n45  &  (~ n351) ) ;
 assign n213 = ( n214  &  n215  &  n31 ) | ( n214  &  n215  &  n206 ) ;
 assign n218 = ( n323  &  n213 ) | ( n359  &  n213 ) | ( n323  &  n96 ) | ( n359  &  n96 ) ;
 assign n217 = ( n253  &  n257 ) | ( (~ n253)  &  (~ n257) ) ;
 assign n220 = ( n378  &  n41 ) | ( n207  &  n41 ) | ( n378  &  n45 ) | ( n207  &  n45 ) ;
 assign n221 = ( n408  &  n382  &  n17 ) | ( n408  &  n382  &  n360 ) ;
 assign n219 = ( n220  &  n221  &  n39 ) | ( n220  &  n221  &  n93 ) ;
 assign n223 = ( (~ PinA10)  &  (~ n179)  &  n329 ) | ( n20  &  (~ n179)  &  n329 ) ;
 assign n222 = ( n82  &  n219 ) | ( n223  &  n219 ) | ( n82  &  n84 ) | ( n223  &  n84 ) ;
 assign n224 = ( n109 ) | ( n255 ) | ( (~ n344) ) ;
 assign n225 = ( n219 ) | ( n120 ) ;
 assign n226 = ( (~ PinD1)  &  (~ PinB1) ) | ( (~ PinB1)  &  n18 ) | ( (~ PinD1)  &  n20 ) | ( n18  &  n20 ) ;
 assign n231 = ( n411  &  n132 ) | ( n207  &  n132 ) | ( n411  &  n45 ) | ( n207  &  n45 ) ;
 assign n232 = ( n410  &  n140 ) | ( n410  &  n360 ) ;
 assign n230 = ( Psh2  &  n111 ) | ( (~ Psh2)  &  n153 ) | ( n111  &  n153 ) ;
 assign n229 = ( n231  &  n232  &  n230 ) | ( n231  &  n232  &  n93 ) ;
 assign n233 = ( n109  &  n330 ) | ( n330  &  (~ n334) ) | ( n109  &  n359 ) | ( (~ n334)  &  n359 ) ;
 assign n234 = ( (~ PinD0)  &  (~ PinB0) ) | ( (~ PinB0)  &  n18 ) | ( (~ PinD0)  &  n20 ) | ( n18  &  n20 ) ;
 assign n239 = ( n140  &  n411 ) | ( n45  &  n411 ) | ( n140  &  n93 ) | ( n45  &  n93 ) ;
 assign n240 = ( n414  &  n415  &  n153 ) | ( n414  &  n415  &  n360 ) ;
 assign n237 = ( (~ n186)  &  n239  &  n240 ) | ( n234  &  n239  &  n240 ) ;
 assign n241 = ( n336  &  n340 ) | ( n359  &  n340 ) | ( n336  &  n109 ) | ( n359  &  n109 ) ;
 assign n244 = ( n79  &  (~ n341) ) ;
 assign n242 = ( n244  &  n253 ) | ( (~ n244)  &  (~ n253) ) ;
 assign n245 = ( n63  &  (~ n341) ) ;
 assign n247 = ( n60  &  (~ n341) ) ;
 assign n246 = ( n247  &  n253 ) | ( (~ n247)  &  (~ n253) ) ;
 assign n249 = ( n66  &  (~ n341) ) ;
 assign n248 = ( n249  &  n253 ) | ( (~ n249)  &  (~ n253) ) ;
 assign n251 = ( n69  &  (~ n341) ) ;
 assign n250 = ( n251  &  n253 ) | ( (~ n251)  &  (~ n253) ) ;
 assign n253 = ( n162  &  (~ n341) ) ;
 assign n254 = ( n341 ) | ( (~ n376) ) ;
 assign n252 = ( (~ n253)  &  n254 ) | ( n253  &  (~ n254) ) ;
 assign n256 = ( n180  &  (~ n341) ) ;
 assign n255 = ( n253  &  n256 ) | ( (~ n253)  &  (~ n256) ) ;
 assign n257 = ( n177  &  (~ n341) ) ;
 assign n261 = ( (~ PinC9) ) | ( n164  &  n309 ) ;
 assign n263 = ( n72  &  (~ n341) ) ;
 assign n262 = ( n253  &  n263 ) | ( (~ n253)  &  (~ n263) ) ;
 assign n265 = ( n57  &  (~ n341) ) ;
 assign n264 = ( n253  &  n265 ) | ( (~ n253)  &  (~ n265) ) ;
 assign n266 = ( n54  &  (~ n341) ) ;
 assign n268 = ( n49  &  (~ n341) ) ;
 assign n267 = ( n253  &  n268 ) | ( (~ n253)  &  (~ n268) ) ;
 assign n273 = ( (~ PinC7) ) | ( n164  &  n309 ) ;
 assign n270 = ( (~ PinA7)  &  (~ n48)  &  n273 ) | ( n20  &  (~ n48)  &  n273 ) ;
 assign n274 = ( (~ n106)  &  n107 ) | ( n106  &  (~ n107) ) ;
 assign n277 = ( (~ PinC6) ) | ( n164  &  n309 ) ;
 assign n279 = ( n262 ) | ( n343 ) ;
 assign n278 = ( (~ n279)  &  n264 ) | ( n279  &  (~ n264) ) ;
 assign n282 = ( (~ PinC5) ) | ( n164  &  n309 ) ;
 assign n283 = ( n262  &  n343 ) | ( (~ n262)  &  (~ n343) ) ;
 assign n288 = ( (~ PinC4) ) | ( n164  &  n309 ) ;
 assign n285 = ( (~ PinA4)  &  (~ n71)  &  n288 ) | ( n20  &  (~ n71)  &  n288 ) ;
 assign n289 = ( n147  &  n246 ) | ( (~ n147)  &  (~ n246) ) ;
 assign n293 = ( (~ PinC3) ) | ( n164  &  n309 ) ;
 assign n294 = ( (~ n148)  &  n149 ) | ( n148  &  (~ n149) ) ;
 assign n298 = ( (~ PinC2) ) | ( n164  &  n309 ) ;
 assign n295 = ( (~ PinA2)  &  (~ n62)  &  n298 ) | ( n20  &  (~ n62)  &  n298 ) ;
 assign n300 = ( n174  &  (~ n341) ) ;
 assign n299 = ( n253  &  n300 ) | ( (~ n253)  &  (~ n300) ) ;
 assign n302 = ( n168  &  (~ n341) ) ;
 assign n301 = ( n253  &  n302 ) | ( (~ n253)  &  (~ n302) ) ;
 assign n303 = ( n171  &  (~ n341) ) ;
 assign n306 = ( (~ PinC15) ) | ( n164  &  n309 ) ;
 assign n307 = ( n188  &  n301 ) | ( (~ n188)  &  (~ n301) ) ;
 assign n312 = ( (~ PinC14)  &  (~ PinA14) ) | ( (~ PinC14)  &  n20 ) | ( (~ PinA14)  &  n164 ) | ( n20  &  n164 ) ;
 assign n309 = ( (~ Pmusel4) ) | ( Pmusel3 ) | ( Pmusel2 ) | ( Pmusel1 ) ;
 assign n313 = ( (~ n189)  &  n190 ) | ( n189  &  (~ n190) ) ;
 assign n316 = ( (~ PinC13)  &  (~ PinA13) ) | ( (~ PinC13)  &  n20 ) | ( (~ PinA13)  &  n164 ) | ( n20  &  n164 ) ;
 assign n318 = ( n262 ) | ( n264 ) | ( n107 ) | ( n267 ) | ( n344 ) ;
 assign n317 = ( (~ n318)  &  n299 ) | ( n318  &  (~ n299) ) ;
 assign n322 = ( (~ PinC12)  &  (~ PinA12) ) | ( (~ PinC12)  &  n20 ) | ( (~ PinA12)  &  n164 ) | ( n20  &  n164 ) ;
 assign n319 = ( (~ PinC12)  &  (~ n173)  &  n322 ) | ( (~ n173)  &  n309  &  n322 ) ;
 assign n326 = ( (~ PinC11) ) | ( n164  &  n309 ) ;
 assign n323 = ( (~ PinA11)  &  (~ n176)  &  n326 ) | ( n20  &  (~ n176)  &  n326 ) ;
 assign n329 = ( (~ PinC10) ) | ( n164  &  n309 ) ;
 assign n333 = ( (~ PinC1) ) | ( n164  &  n309 ) ;
 assign n330 = ( (~ PinA1)  &  (~ n65)  &  n333 ) | ( n20  &  (~ n65)  &  n333 ) ;
 assign n335 = ( n250 ) | ( (~ n253) ) ;
 assign n334 = ( (~ n335)  &  n248 ) | ( n335  &  (~ n248) ) ;
 assign n339 = ( (~ PinC0) ) | ( n164  &  n309 ) ;
 assign n336 = ( (~ PinA0)  &  (~ n68)  &  n339 ) | ( n20  &  (~ n68)  &  n339 ) ;
 assign n340 = ( (~ n250)  &  n253 ) | ( n250  &  (~ n253) ) ;
 assign n341 = ( (~ Pmusel4) ) | ( Pmusel3 ) | ( n34 ) ;
 assign n343 = ( n149 ) | ( n246 ) | ( n248 ) | ( n250 ) | ( (~ n253) ) ;
 assign n344 = ( n242 ) | ( n252 ) | ( n255 ) | ( n217 ) | ( n343 ) ;
 assign n345 = ( Popsel2  &  n84 ) | ( (~ Popsel2)  &  (~ n84) ) ;
 assign n348 = ( (~ Pmusel3) ) | ( Pmusel2 ) | ( Pmusel1 ) ;
 assign n349 = ( Pmusel3 ) | ( (~ Pmusel2) ) | ( Pmusel1 ) ;
 assign n351 = ( (~ Psh1) ) | ( (~ Psh0) ) ;
 assign n353 = ( (~ Psh1) ) | ( Psh0 ) ;
 assign n354 = ( Popsel3  &  (~ Popsel2) ) ;
 assign n359 = ( n82 ) | ( (~ n354) ) ;
 assign n360 = ( Psh2 ) | ( n353 ) ;
 assign n363 = ( (~ Psh2) ) | ( n353 ) ;
 assign n376 = ( Pmusel2  &  PinC8 ) | ( (~ Pmusel2)  &  PinA8 ) | ( PinC8  &  PinA8 ) ;
 assign n377 = ( (~ PinD9)  &  (~ PinB9) ) | ( (~ PinB9)  &  n348 ) | ( (~ PinD9)  &  n349 ) | ( n348  &  n349 ) ;
 assign n378 = ( Psh2  &  n25 ) | ( (~ Psh2)  &  n28 ) | ( n25  &  n28 ) ;
 assign n379 = ( Pmusel4  &  (~ PinA8) ) | ( Pmusel4  &  n20 ) | ( (~ PinA8)  &  n74 ) | ( n20  &  n74 ) ;
 assign n380 = ( (~ PinC8) ) | ( n164  &  n309 ) ;
 assign n381 = ( n88 ) | ( n208 ) ;
 assign n382 = ( n353 ) | ( n40 ) ;
 assign n383 = ( n109 ) | ( n252 ) | ( (~ n344) ) ;
 assign n384 = ( (~ PinD7)  &  (~ PinB7) ) | ( (~ PinB7)  &  n348 ) | ( (~ PinD7)  &  n349 ) | ( n348  &  n349 ) ;
 assign n385 = ( n98 ) | ( n208 ) ;
 assign n386 = ( (~ PinD6)  &  (~ PinB6) ) | ( (~ PinB6)  &  n348 ) | ( (~ PinD6)  &  n349 ) | ( n348  &  n349 ) ;
 assign n387 = ( n25  &  n111 ) | ( n363  &  n111 ) | ( n25  &  n208 ) | ( n363  &  n208 ) ;
 assign n389 = ( (~ PinD5)  &  (~ PinB5) ) | ( (~ PinB5)  &  n348 ) | ( (~ PinD5)  &  n349 ) | ( n348  &  n349 ) ;
 assign n390 = ( n41  &  n122 ) | ( n363  &  n122 ) | ( n41  &  n208 ) | ( n363  &  n208 ) ;
 assign n392 = ( (~ PinD4)  &  (~ PinB4) ) | ( (~ PinB4)  &  n348 ) | ( (~ PinD4)  &  n349 ) | ( n348  &  n349 ) ;
 assign n393 = ( n17  &  n132 ) | ( n363  &  n132 ) | ( n17  &  n208 ) | ( n363  &  n208 ) ;
 assign n394 = ( (~ PinD3)  &  (~ PinB3) ) | ( (~ PinB3)  &  n348 ) | ( (~ PinD3)  &  n349 ) | ( n348  &  n349 ) ;
 assign n395 = ( n31  &  n140 ) | ( n363  &  n140 ) | ( n31  &  n208 ) | ( n363  &  n208 ) ;
 assign n396 = ( (~ PinD2)  &  (~ PinB2) ) | ( (~ PinB2)  &  n348 ) | ( (~ PinD2)  &  n349 ) | ( n348  &  n349 ) ;
 assign n397 = ( n28  &  n153 ) | ( n363  &  n153 ) | ( n28  &  n208 ) | ( n363  &  n208 ) ;
 assign n399 = ( (~ PinD15)  &  (~ PinB15) ) | ( (~ PinB15)  &  n348 ) | ( (~ PinD15)  &  n349 ) | ( n348  &  n349 ) ;
 assign n400 = ( (~ PinD14)  &  (~ PinB14) ) | ( (~ PinB14)  &  n348 ) | ( (~ PinD14)  &  n349 ) | ( n348  &  n349 ) ;
 assign n401 = ( (~ PinD13)  &  (~ PinB13) ) | ( (~ PinB13)  &  n348 ) | ( (~ PinD13)  &  n349 ) | ( n348  &  n349 ) ;
 assign n403 = ( (~ PinD12)  &  (~ PinB12) ) | ( (~ PinB12)  &  n348 ) | ( (~ PinD12)  &  n349 ) | ( n348  &  n349 ) ;
 assign n406 = ( (~ PinD11)  &  (~ PinB11) ) | ( (~ PinB11)  &  n348 ) | ( (~ PinD11)  &  n349 ) | ( n348  &  n349 ) ;
 assign n407 = ( (~ PinD10)  &  (~ PinB10) ) | ( (~ PinB10)  &  n348 ) | ( (~ PinD10)  &  n349 ) | ( n348  &  n349 ) ;
 assign n408 = ( n28 ) | ( n208 ) ;
 assign n409 = ( (~ PinD1)  &  (~ PinB1) ) | ( (~ PinB1)  &  n348 ) | ( (~ PinD1)  &  n349 ) | ( n348  &  n349 ) ;
 assign n410 = ( n22  &  n226 ) | ( n363  &  n226 ) | ( n22  &  n208 ) | ( n363  &  n208 ) ;
 assign n411 = ( Psh2  &  n122 ) | ( (~ Psh2)  &  n226 ) | ( n122  &  n226 ) ;
 assign n413 = ( (~ PinD0)  &  (~ PinB0) ) | ( (~ PinB0)  &  n348 ) | ( (~ PinD0)  &  n349 ) | ( n348  &  n349 ) ;
 assign n414 = ( n88 ) | ( n363 ) ;
 assign n415 = ( (~ Psh2) ) | ( n132 ) | ( n207 ) ;


endmodule

