module i8 (
	PV133_10_, PV133_9_, PV133_8_, PV133_7_, PV133_6_, PV133_5_, PV133_4_, PV133_3_, 
	PV133_2_, PV133_1_, PV133_0_, PV122_0_, PV121_17_, PV121_16_, PV119_0_, PV118_1_, PV118_0_, PV116_31_, 
	PV116_30_, PV116_29_, PV116_28_, PV116_27_, PV116_26_, PV116_25_, PV116_24_, PV116_23_, PV116_22_, PV116_21_, 
	PV116_20_, PV116_19_, PV116_18_, PV116_17_, PV116_16_, PV116_15_, PV116_14_, PV116_13_, PV116_12_, PV116_11_, 
	PV116_10_, PV116_9_, PV116_8_, PV116_7_, PV116_6_, PV116_5_, PV116_4_, PV116_3_, PV116_2_, PV116_1_, 
	PV116_0_, PV84_31_, PV84_30_, PV84_29_, PV84_28_, PV84_27_, PV84_26_, PV84_25_, PV84_24_, PV84_23_, 
	PV84_22_, PV84_21_, PV84_20_, PV84_19_, PV84_18_, PV84_17_, PV84_16_, PV84_15_, PV84_14_, PV84_13_, 
	PV84_12_, PV84_11_, PV84_10_, PV84_9_, PV84_8_, PV84_7_, PV84_6_, PV84_5_, PV84_4_, PV84_3_, 
	PV84_2_, PV84_1_, PV84_0_, PV52_0_, PV51_0_, PV50_0_, PV49_0_, PV48_0_, PV47_31_, PV47_30_, 
	PV47_29_, PV47_28_, PV47_27_, PV47_26_, PV47_25_, PV47_24_, PV47_23_, PV47_22_, PV47_21_, PV47_20_, 
	PV47_19_, PV47_18_, PV47_17_, PV47_16_, PV47_15_, PV47_14_, PV47_13_, PV47_12_, PV47_11_, PV47_10_, 
	PV47_9_, PV47_8_, PV47_7_, PV47_6_, PV47_5_, PV47_4_, PV47_3_, PV47_2_, PV47_1_, PV47_0_, 
	PV15_14_, PV15_13_, PV15_12_, PV15_11_, PV15_10_, PV15_9_, PV15_8_, PV15_7_, PV15_6_, PV15_5_, 
	PV15_4_, PV15_3_, PV15_2_, PV15_1_, PV15_0_, PV214_0_, PV213_0_, PV212_14_, PV212_13_, PV212_12_, 
	PV212_11_, PV212_10_, PV212_9_, PV212_8_, PV212_7_, PV212_6_, PV212_5_, PV212_4_, PV212_3_, PV212_2_, 
	PV212_1_, PV212_0_, PV197_31_, PV197_30_, PV197_29_, PV197_28_, PV197_27_, PV197_26_, PV197_25_, PV197_24_, 
	PV197_23_, PV197_22_, PV197_21_, PV197_20_, PV197_19_, PV197_18_, PV197_17_, PV197_16_, PV197_15_, PV197_14_, 
	PV197_13_, PV197_12_, PV197_11_, PV197_10_, PV197_9_, PV197_8_, PV197_7_, PV197_6_, PV197_5_, PV197_4_, 
	PV197_3_, PV197_2_, PV197_1_, PV197_0_, PV165_14_, PV165_13_, PV165_12_, PV165_11_, PV165_10_, PV165_9_, 
	PV165_8_, PV165_7_, PV165_6_, PV165_5_, PV165_4_, PV165_3_, PV165_2_, PV165_1_, PV165_0_, PV150_0_, 
	PV149_2_, PV149_1_, PV149_0_, PV146_0_, PV145_1_, PV145_0_, PV143_0_, PV142_5_, PV142_4_, PV142_3_, 
	PV142_2_, PV142_1_, PV142_0_, PV136_1_, PV136_0_, PV134_0_);

input PV133_10_, PV133_9_, PV133_8_, PV133_7_, PV133_6_, PV133_5_, PV133_4_, PV133_3_, PV133_2_, PV133_1_, PV133_0_, PV122_0_, PV121_17_, PV121_16_, PV119_0_, PV118_1_, PV118_0_, PV116_31_, PV116_30_, PV116_29_, PV116_28_, PV116_27_, PV116_26_, PV116_25_, PV116_24_, PV116_23_, PV116_22_, PV116_21_, PV116_20_, PV116_19_, PV116_18_, PV116_17_, PV116_16_, PV116_15_, PV116_14_, PV116_13_, PV116_12_, PV116_11_, PV116_10_, PV116_9_, PV116_8_, PV116_7_, PV116_6_, PV116_5_, PV116_4_, PV116_3_, PV116_2_, PV116_1_, PV116_0_, PV84_31_, PV84_30_, PV84_29_, PV84_28_, PV84_27_, PV84_26_, PV84_25_, PV84_24_, PV84_23_, PV84_22_, PV84_21_, PV84_20_, PV84_19_, PV84_18_, PV84_17_, PV84_16_, PV84_15_, PV84_14_, PV84_13_, PV84_12_, PV84_11_, PV84_10_, PV84_9_, PV84_8_, PV84_7_, PV84_6_, PV84_5_, PV84_4_, PV84_3_, PV84_2_, PV84_1_, PV84_0_, PV52_0_, PV51_0_, PV50_0_, PV49_0_, PV48_0_, PV47_31_, PV47_30_, PV47_29_, PV47_28_, PV47_27_, PV47_26_, PV47_25_, PV47_24_, PV47_23_, PV47_22_, PV47_21_, PV47_20_, PV47_19_, PV47_18_, PV47_17_, PV47_16_, PV47_15_, PV47_14_, PV47_13_, PV47_12_, PV47_11_, PV47_10_, PV47_9_, PV47_8_, PV47_7_, PV47_6_, PV47_5_, PV47_4_, PV47_3_, PV47_2_, PV47_1_, PV47_0_, PV15_14_, PV15_13_, PV15_12_, PV15_11_, PV15_10_, PV15_9_, PV15_8_, PV15_7_, PV15_6_, PV15_5_, PV15_4_, PV15_3_, PV15_2_, PV15_1_, PV15_0_;

output PV214_0_, PV213_0_, PV212_14_, PV212_13_, PV212_12_, PV212_11_, PV212_10_, PV212_9_, PV212_8_, PV212_7_, PV212_6_, PV212_5_, PV212_4_, PV212_3_, PV212_2_, PV212_1_, PV212_0_, PV197_31_, PV197_30_, PV197_29_, PV197_28_, PV197_27_, PV197_26_, PV197_25_, PV197_24_, PV197_23_, PV197_22_, PV197_21_, PV197_20_, PV197_19_, PV197_18_, PV197_17_, PV197_16_, PV197_15_, PV197_14_, PV197_13_, PV197_12_, PV197_11_, PV197_10_, PV197_9_, PV197_8_, PV197_7_, PV197_6_, PV197_5_, PV197_4_, PV197_3_, PV197_2_, PV197_1_, PV197_0_, PV165_14_, PV165_13_, PV165_12_, PV165_11_, PV165_10_, PV165_9_, PV165_8_, PV165_7_, PV165_6_, PV165_5_, PV165_4_, PV165_3_, PV165_2_, PV165_1_, PV165_0_, PV150_0_, PV149_2_, PV149_1_, PV149_0_, PV146_0_, PV145_1_, PV145_0_, PV143_0_, PV142_5_, PV142_4_, PV142_3_, PV142_2_, PV142_1_, PV142_0_, PV136_1_, PV136_0_, PV134_0_;

wire n1, n6, n7, n5, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n73, n71, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n94, n93, n91, n95, n96, n102, n100, n99, n105, n103, n108, n109, n113, n111, n117, n118, n115, n122, n123, n120, n127, n128, n125, n132, n133, n130, n137, n138, n135, n142, n143, n140, n147, n148, n145, n152, n153, n150, n157, n158, n155, n162, n163, n160, n167, n168, n165, n172, n173, n170, n177, n176, n175, n179, n181, n183, n185, n187, n189, n191, n193, n195, n197, n199, n201, n203, n205, n207, n208, n210, n212, n213, n211, n216, n215, n214, n219, n217, n221, n220, n224, n223, n225, n229, n227, n230, n231, n234, n233, n235, n238, n237, n239, n242, n241, n243, n246, n245, n247, n250, n249, n251, n255, n253, n257, n256, n258, n262, n260, n263, n267, n265, n270, n271, n268, n273, n272, n275, n274, n279, n278, n276, n277, n282, n280, n281, n285, n283, n284, n286, n289, n287, n288, n292, n290, n291, n295, n293, n294, n298, n296, n297, n301, n299, n300, n304, n302, n303, n307, n305, n306, n310, n308, n309, n313, n311, n312, n316, n314, n315, n319, n317, n318, n322, n320, n321, n325, n323, n324, n328, n326, n327, n331, n329, n330, n334, n332, n333, n336, n337, n335, n340, n341, n339, n344, n345, n343, n348, n349, n347, n353, n354, n351, n358, n359, n356, n363, n364, n361, n367, n368, n366, n371, n372, n370, n375, n374, n378, n377, n381, n380, n384, n383, n387, n386, n390, n389, n393, n392, n396, n395, n399, n398, n402, n401, n403, n404, n405, n408, n409, n411, n412, n418, n437, n447, n448, n449, n450, n451, n452, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n474, n479, n481, n485, n486;

assign PV214_0_ = ( (~ n449) ) ;
 assign PV213_0_ = ( (~ n448) ) ;
 assign PV212_14_ = ( (~ n74) ) ;
 assign PV212_13_ = ( (~ n75) ) ;
 assign PV212_12_ = ( (~ n76) ) ;
 assign PV212_11_ = ( (~ n77) ) ;
 assign PV212_10_ = ( (~ n78) ) ;
 assign PV212_9_ = ( (~ n79) ) ;
 assign PV212_8_ = ( (~ n80) ) ;
 assign PV212_7_ = ( (~ n81) ) ;
 assign PV212_6_ = ( (~ n82) ) ;
 assign PV212_5_ = ( (~ n83) ) ;
 assign PV212_4_ = ( (~ n84) ) ;
 assign PV212_3_ = ( (~ n85) ) ;
 assign PV212_2_ = ( (~ n86) ) ;
 assign PV212_1_ = ( (~ n87) ) ;
 assign PV212_0_ = ( (~ n88) ) ;
 assign PV197_31_ = ( (~ n39) ) ;
 assign PV197_30_ = ( (~ n40) ) ;
 assign PV197_29_ = ( (~ n41) ) ;
 assign PV197_28_ = ( (~ n42) ) ;
 assign PV197_27_ = ( (~ n43) ) ;
 assign PV197_26_ = ( (~ n44) ) ;
 assign PV197_25_ = ( (~ n45) ) ;
 assign PV197_24_ = ( (~ n46) ) ;
 assign PV197_23_ = ( (~ n47) ) ;
 assign PV197_22_ = ( (~ n48) ) ;
 assign PV197_21_ = ( (~ n49) ) ;
 assign PV197_20_ = ( (~ n50) ) ;
 assign PV197_19_ = ( (~ n51) ) ;
 assign PV197_18_ = ( (~ n52) ) ;
 assign PV197_17_ = ( (~ n53) ) ;
 assign PV197_16_ = ( (~ n54) ) ;
 assign PV197_15_ = ( (~ n55) ) ;
 assign PV197_14_ = ( (~ n56) ) ;
 assign PV197_13_ = ( (~ n57) ) ;
 assign PV197_12_ = ( (~ n58) ) ;
 assign PV197_11_ = ( (~ n59) ) ;
 assign PV197_10_ = ( (~ n60) ) ;
 assign PV197_9_ = ( (~ n61) ) ;
 assign PV197_8_ = ( (~ n62) ) ;
 assign PV197_7_ = ( (~ n63) ) ;
 assign PV197_6_ = ( (~ n64) ) ;
 assign PV197_5_ = ( (~ n65) ) ;
 assign PV197_4_ = ( (~ n66) ) ;
 assign PV197_3_ = ( (~ n67) ) ;
 assign PV197_2_ = ( (~ n68) ) ;
 assign PV197_1_ = ( (~ n69) ) ;
 assign PV197_0_ = ( (~ n70) ) ;
 assign PV165_14_ = ( (~ n24) ) ;
 assign PV165_13_ = ( (~ n25) ) ;
 assign PV165_12_ = ( (~ n26) ) ;
 assign PV165_11_ = ( (~ n27) ) ;
 assign PV165_10_ = ( (~ n28) ) ;
 assign PV165_9_ = ( (~ n29) ) ;
 assign PV165_8_ = ( (~ n30) ) ;
 assign PV165_7_ = ( (~ n31) ) ;
 assign PV165_6_ = ( (~ n32) ) ;
 assign PV165_5_ = ( (~ n33) ) ;
 assign PV165_4_ = ( (~ n34) ) ;
 assign PV165_3_ = ( (~ n35) ) ;
 assign PV165_2_ = ( (~ n36) ) ;
 assign PV165_1_ = ( (~ n37) ) ;
 assign PV165_0_ = ( (~ n38) ) ;
 assign PV150_0_ = ( (~ n23) ) ;
 assign PV149_2_ = ( (~ n20) ) ;
 assign PV149_1_ = ( (~ n21) ) ;
 assign PV149_0_ = ( (~ n22) ) ;
 assign PV146_0_ = ( (~ n19) ) ;
 assign PV145_1_ = ( (~ n17) ) ;
 assign PV145_0_ = ( (~ n18) ) ;
 assign PV143_0_ = ( (~ n16) ) ;
 assign PV142_5_ = ( (~ n10) ) ;
 assign PV142_4_ = ( (~ n11) ) ;
 assign PV142_3_ = ( (~ n12) ) ;
 assign PV142_2_ = ( (~ n13) ) ;
 assign PV142_1_ = ( (~ n14) ) ;
 assign PV142_0_ = ( (~ n15) ) ;
 assign PV136_1_ = ( (~ n8) ) ;
 assign PV136_0_ = ( (~ n9) ) ;
 assign PV134_0_ = ( (~ n450) ) ;
 assign n1 = ( PV133_7_  &  (~ PV133_2_)  &  (~ PV133_1_) ) | ( (~ PV133_2_)  &  (~ PV133_1_)  &  (~ n93) ) ;
 assign n6 = ( (~ PV133_2_) ) | ( (~ PV133_1_) ) ;
 assign n7 = ( PV133_9_ ) | ( PV133_4_ ) ;
 assign n5 = ( n6 ) | ( PV133_8_ ) | ( n7 ) ;
 assign n8 = ( (~ n217)  &  n221 ) | ( n99  &  (~ n217)  &  n220 ) ;
 assign n9 = ( n224  &  n221 ) | ( n224  &  n223  &  n109 ) ;
 assign n10 = ( (~ PV116_8_)  &  n227 ) | ( (~ PV116_8_)  &  n230 ) | ( n227  &  (~ n404) ) | ( n230  &  (~ n404) ) ;
 assign n11 = ( n234  &  n230 ) | ( n234  &  n233  &  n231 ) ;
 assign n12 = ( n238  &  n230 ) | ( n238  &  n237  &  n235 ) ;
 assign n13 = ( n242  &  n230 ) | ( n242  &  n241  &  n239 ) ;
 assign n14 = ( n246  &  n230 ) | ( n246  &  n245  &  n243 ) ;
 assign n15 = ( n250  &  n230 ) | ( n250  &  n249  &  n247 ) ;
 assign n16 = ( (~ PV116_9_)  &  n253 ) | ( (~ PV116_9_)  &  n256 ) | ( n253  &  (~ n404) ) | ( n256  &  (~ n404) ) ;
 assign n17 = ( (~ PV116_11_)  &  n230 ) | ( (~ PV116_11_)  &  n260 ) | ( n230  &  (~ n404) ) | ( n260  &  (~ n404) ) ;
 assign n18 = ( (~ PV116_10_)  &  n230 ) | ( (~ PV116_10_)  &  n265 ) | ( n230  &  (~ n404) ) | ( n265  &  (~ n404) ) ;
 assign n19 = ( n275  &  n268 ) | ( n275  &  n272  &  n274 ) ;
 assign n20 = ( n279  &  n278 ) | ( n279  &  n276  &  n277 ) ;
 assign n21 = ( n282  &  n278 ) | ( n282  &  n280  &  n281 ) ;
 assign n22 = ( n285  &  n278 ) | ( n285  &  n283  &  n284 ) ;
 assign n23 = ( n289  &  n286 ) | ( n289  &  n287  &  n288 ) ;
 assign n24 = ( n292  &  n278 ) | ( n292  &  n290  &  n291 ) ;
 assign n25 = ( n295  &  n278 ) | ( n295  &  n293  &  n294 ) ;
 assign n26 = ( n298  &  n278 ) | ( n298  &  n296  &  n297 ) ;
 assign n27 = ( n301  &  n278 ) | ( n301  &  n299  &  n300 ) ;
 assign n28 = ( n304  &  n278 ) | ( n304  &  n302  &  n303 ) ;
 assign n29 = ( n307  &  n278 ) | ( n307  &  n305  &  n306 ) ;
 assign n30 = ( n310  &  n278 ) | ( n310  &  n308  &  n309 ) ;
 assign n31 = ( n313  &  n278 ) | ( n313  &  n311  &  n312 ) ;
 assign n32 = ( n316  &  n278 ) | ( n316  &  n314  &  n315 ) ;
 assign n33 = ( n319  &  n278 ) | ( n319  &  n317  &  n318 ) ;
 assign n34 = ( n322  &  n278 ) | ( n322  &  n320  &  n321 ) ;
 assign n35 = ( n325  &  n278 ) | ( n325  &  n323  &  n324 ) ;
 assign n36 = ( n328  &  n278 ) | ( n328  &  n326  &  n327 ) ;
 assign n37 = ( n331  &  n278 ) | ( n331  &  n329  &  n330 ) ;
 assign n38 = ( n334  &  n278 ) | ( n334  &  n332  &  n333 ) ;
 assign n39 = ( (~ PV116_31_)  &  n108 ) | ( (~ PV116_31_)  &  n335 ) | ( n108  &  (~ n404) ) | ( n335  &  (~ n404) ) ;
 assign n40 = ( (~ PV116_30_)  &  n108 ) | ( (~ PV116_30_)  &  n339 ) | ( n108  &  (~ n404) ) | ( n339  &  (~ n404) ) ;
 assign n41 = ( (~ PV116_29_)  &  n108 ) | ( (~ PV116_29_)  &  n343 ) | ( n108  &  (~ n404) ) | ( n343  &  (~ n404) ) ;
 assign n42 = ( (~ PV116_28_)  &  n108 ) | ( (~ PV116_28_)  &  n347 ) | ( n108  &  (~ n404) ) | ( n347  &  (~ n404) ) ;
 assign n43 = ( (~ PV116_27_)  &  n108 ) | ( (~ PV116_27_)  &  n351 ) | ( n108  &  (~ n404) ) | ( n351  &  (~ n404) ) ;
 assign n44 = ( (~ PV116_26_)  &  n108 ) | ( (~ PV116_26_)  &  n356 ) | ( n108  &  (~ n404) ) | ( n356  &  (~ n404) ) ;
 assign n45 = ( (~ PV116_25_)  &  n108 ) | ( (~ PV116_25_)  &  n361 ) | ( n108  &  (~ n404) ) | ( n361  &  (~ n404) ) ;
 assign n46 = ( (~ PV116_24_)  &  n108 ) | ( (~ PV116_24_)  &  n366 ) | ( n108  &  (~ n404) ) | ( n366  &  (~ n404) ) ;
 assign n47 = ( (~ PV116_23_)  &  n108 ) | ( (~ PV116_23_)  &  n370 ) | ( n108  &  (~ n404) ) | ( n370  &  (~ n404) ) ;
 assign n48 = ( (~ PV116_22_)  &  n108 ) | ( (~ PV116_22_)  &  n374 ) | ( n108  &  (~ n404) ) | ( n374  &  (~ n404) ) ;
 assign n49 = ( (~ PV116_21_)  &  n108 ) | ( (~ PV116_21_)  &  n377 ) | ( n108  &  (~ n404) ) | ( n377  &  (~ n404) ) ;
 assign n50 = ( (~ PV116_20_)  &  n108 ) | ( (~ PV116_20_)  &  n380 ) | ( n108  &  (~ n404) ) | ( n380  &  (~ n404) ) ;
 assign n51 = ( (~ PV116_19_)  &  n108 ) | ( (~ PV116_19_)  &  n383 ) | ( n108  &  (~ n404) ) | ( n383  &  (~ n404) ) ;
 assign n52 = ( (~ PV116_18_)  &  n108 ) | ( (~ PV116_18_)  &  n386 ) | ( n108  &  (~ n404) ) | ( n386  &  (~ n404) ) ;
 assign n53 = ( (~ PV116_17_)  &  n108 ) | ( (~ PV116_17_)  &  n389 ) | ( n108  &  (~ n404) ) | ( n389  &  (~ n404) ) ;
 assign n54 = ( (~ PV116_16_)  &  n108 ) | ( (~ PV116_16_)  &  n392 ) | ( n108  &  (~ n404) ) | ( n392  &  (~ n404) ) ;
 assign n55 = ( (~ PV116_15_)  &  n108 ) | ( (~ PV116_15_)  &  n395 ) | ( n108  &  (~ n404) ) | ( n395  &  (~ n404) ) ;
 assign n56 = ( (~ PV116_14_)  &  n108 ) | ( (~ PV116_14_)  &  n398 ) | ( n108  &  (~ n404) ) | ( n398  &  (~ n404) ) ;
 assign n57 = ( (~ PV116_13_)  &  n103 ) | ( (~ PV116_13_)  &  n108 ) | ( n103  &  (~ n404) ) | ( n108  &  (~ n404) ) ;
 assign n58 = ( (~ PV116_12_)  &  n108 ) | ( (~ PV116_12_)  &  n111 ) | ( n108  &  (~ n404) ) | ( n111  &  (~ n404) ) ;
 assign n59 = ( (~ PV116_11_)  &  n108 ) | ( (~ PV116_11_)  &  n115 ) | ( n108  &  (~ n404) ) | ( n115  &  (~ n404) ) ;
 assign n60 = ( (~ PV116_10_)  &  n108 ) | ( (~ PV116_10_)  &  n120 ) | ( n108  &  (~ n404) ) | ( n120  &  (~ n404) ) ;
 assign n61 = ( (~ PV116_9_)  &  n108 ) | ( (~ PV116_9_)  &  n125 ) | ( n108  &  (~ n404) ) | ( n125  &  (~ n404) ) ;
 assign n62 = ( (~ PV116_8_)  &  n108 ) | ( (~ PV116_8_)  &  n130 ) | ( n108  &  (~ n404) ) | ( n130  &  (~ n404) ) ;
 assign n63 = ( (~ PV116_7_)  &  n108 ) | ( (~ PV116_7_)  &  n135 ) | ( n108  &  (~ n404) ) | ( n135  &  (~ n404) ) ;
 assign n64 = ( (~ PV116_6_)  &  n108 ) | ( (~ PV116_6_)  &  n140 ) | ( n108  &  (~ n404) ) | ( n140  &  (~ n404) ) ;
 assign n65 = ( (~ PV116_5_)  &  n108 ) | ( (~ PV116_5_)  &  n145 ) | ( n108  &  (~ n404) ) | ( n145  &  (~ n404) ) ;
 assign n66 = ( (~ PV116_4_)  &  n108 ) | ( (~ PV116_4_)  &  n150 ) | ( n108  &  (~ n404) ) | ( n150  &  (~ n404) ) ;
 assign n67 = ( (~ PV116_3_)  &  n108 ) | ( (~ PV116_3_)  &  n155 ) | ( n108  &  (~ n404) ) | ( n155  &  (~ n404) ) ;
 assign n68 = ( (~ PV116_2_)  &  n108 ) | ( (~ PV116_2_)  &  n160 ) | ( n108  &  (~ n404) ) | ( n160  &  (~ n404) ) ;
 assign n69 = ( (~ PV116_1_)  &  n108 ) | ( (~ PV116_1_)  &  n165 ) | ( n108  &  (~ n404) ) | ( n165  &  (~ n404) ) ;
 assign n70 = ( (~ PV116_0_)  &  n108 ) | ( (~ PV116_0_)  &  n170 ) | ( n108  &  (~ n404) ) | ( n170  &  (~ n404) ) ;
 assign n73 = ( PV133_6_ ) | ( n7 ) ;
 assign n71 = ( (~ PV133_3_) ) | ( n6 ) | ( n73 ) ;
 assign n74 = ( (~ PV84_31_)  &  n179 ) | ( n175  &  n179 ) ;
 assign n75 = ( (~ PV84_30_)  &  n181 ) | ( n175  &  n181 ) ;
 assign n76 = ( (~ PV84_29_)  &  n183 ) | ( n175  &  n183 ) ;
 assign n77 = ( (~ PV84_28_)  &  n185 ) | ( n175  &  n185 ) ;
 assign n78 = ( (~ PV84_27_)  &  n187 ) | ( n175  &  n187 ) ;
 assign n79 = ( (~ PV84_26_)  &  n189 ) | ( n175  &  n189 ) ;
 assign n80 = ( (~ PV84_25_)  &  n191 ) | ( n175  &  n191 ) ;
 assign n81 = ( (~ PV84_24_)  &  n193 ) | ( n175  &  n193 ) ;
 assign n82 = ( (~ PV84_23_)  &  n195 ) | ( n175  &  n195 ) ;
 assign n83 = ( (~ PV84_22_)  &  n197 ) | ( n175  &  n197 ) ;
 assign n84 = ( (~ PV84_21_)  &  n199 ) | ( n175  &  n199 ) ;
 assign n85 = ( (~ PV84_20_)  &  n201 ) | ( n175  &  n201 ) ;
 assign n86 = ( (~ PV84_19_)  &  n203 ) | ( n175  &  n203 ) ;
 assign n87 = ( (~ PV84_18_)  &  n205 ) | ( n175  &  n205 ) ;
 assign n88 = ( (~ PV84_17_)  &  n207 ) | ( n175  &  n207 ) ;
 assign n89 = ( (~ PV133_10_)  &  (~ PV133_3_) ) | ( (~ PV133_10_)  &  n6 ) ;
 assign n94 = ( PV133_10_ ) | ( n6 ) ;
 assign n93 = ( PV133_5_ ) | ( PV133_6_ ) ;
 assign n91 = ( (~ PV133_2_)  &  n94 ) | ( (~ PV133_8_)  &  n94  &  n93 ) ;
 assign n95 = ( PV133_8_  &  PV133_1_ ) | ( (~ PV133_2_)  &  PV133_1_  &  (~ n93) ) ;
 assign n96 = ( PV133_0_  &  (~ n95) ) | ( (~ PV133_7_)  &  PV133_5_  &  (~ n95) ) ;
 assign n102 = ( n1 ) | ( (~ n91) ) | ( n405 ) ;
 assign n100 = ( n91 ) | ( n405 ) ;
 assign n99 = ( (~ PV84_2_)  &  n102 ) | ( n102  &  n100 ) ;
 assign n105 = ( (~ PV84_5_)  &  (~ PV47_30_) ) | ( (~ PV47_30_)  &  n408 ) | ( (~ PV84_5_)  &  n409 ) | ( n408  &  n409 ) ;
 assign n103 = ( (~ PV84_13_)  &  n99  &  n105 ) | ( n89  &  n99  &  n105 ) ;
 assign n108 = ( (~ PV133_10_)  &  n71  &  n176  &  n213  &  n401  &  n403 ) ;
 assign n109 = ( (~ PV84_1_)  &  n102 ) | ( n102  &  n100 ) ;
 assign n113 = ( (~ PV84_4_)  &  (~ PV47_29_) ) | ( (~ PV47_29_)  &  n408 ) | ( (~ PV84_4_)  &  n409 ) | ( n408  &  n409 ) ;
 assign n111 = ( (~ PV84_12_)  &  n109  &  n113 ) | ( n89  &  n109  &  n113 ) ;
 assign n117 = ( (~ PV84_3_)  &  n102 ) | ( n102  &  n408 ) ;
 assign n118 = ( (~ PV84_11_)  &  (~ PV47_28_) ) | ( (~ PV47_28_)  &  n89 ) | ( (~ PV84_11_)  &  n409 ) | ( n89  &  n409 ) ;
 assign n115 = ( (~ PV84_0_)  &  n117  &  n118 ) | ( n100  &  n117  &  n118 ) ;
 assign n122 = ( (~ PV84_2_)  &  n102 ) | ( n102  &  n408 ) ;
 assign n123 = ( (~ PV84_10_)  &  (~ PV47_27_) ) | ( (~ PV47_27_)  &  n89 ) | ( (~ PV84_10_)  &  n409 ) | ( n89  &  n409 ) ;
 assign n120 = ( (~ PV47_31_)  &  n122  &  n123 ) | ( n100  &  n122  &  n123 ) ;
 assign n127 = ( (~ PV84_1_)  &  n102 ) | ( n102  &  n408 ) ;
 assign n128 = ( (~ PV84_9_)  &  (~ PV47_26_) ) | ( (~ PV47_26_)  &  n89 ) | ( (~ PV84_9_)  &  n409 ) | ( n89  &  n409 ) ;
 assign n125 = ( (~ PV47_30_)  &  n127  &  n128 ) | ( n100  &  n127  &  n128 ) ;
 assign n132 = ( (~ PV84_0_)  &  n102 ) | ( n102  &  n408 ) ;
 assign n133 = ( (~ PV84_8_)  &  (~ PV47_25_) ) | ( (~ PV47_25_)  &  n89 ) | ( (~ PV84_8_)  &  n409 ) | ( n89  &  n409 ) ;
 assign n130 = ( (~ PV47_29_)  &  n132  &  n133 ) | ( n100  &  n132  &  n133 ) ;
 assign n137 = ( (~ PV47_31_)  &  n102 ) | ( n102  &  n408 ) ;
 assign n138 = ( (~ PV84_7_)  &  (~ PV47_24_) ) | ( (~ PV47_24_)  &  n89 ) | ( (~ PV84_7_)  &  n409 ) | ( n89  &  n409 ) ;
 assign n135 = ( (~ PV47_28_)  &  n137  &  n138 ) | ( n100  &  n137  &  n138 ) ;
 assign n142 = ( (~ PV47_30_)  &  n102 ) | ( n102  &  n408 ) ;
 assign n143 = ( (~ PV84_6_)  &  (~ PV47_23_) ) | ( (~ PV47_23_)  &  n89 ) | ( (~ PV84_6_)  &  n409 ) | ( n89  &  n409 ) ;
 assign n140 = ( (~ PV47_27_)  &  n142  &  n143 ) | ( n100  &  n142  &  n143 ) ;
 assign n147 = ( (~ PV47_29_)  &  n102 ) | ( n102  &  n408 ) ;
 assign n148 = ( (~ PV84_5_)  &  (~ PV47_22_) ) | ( (~ PV47_22_)  &  n89 ) | ( (~ PV84_5_)  &  n409 ) | ( n89  &  n409 ) ;
 assign n145 = ( (~ PV47_26_)  &  n147  &  n148 ) | ( n100  &  n147  &  n148 ) ;
 assign n152 = ( (~ PV47_28_)  &  n102 ) | ( n102  &  n408 ) ;
 assign n153 = ( (~ PV84_4_)  &  (~ PV47_21_) ) | ( (~ PV47_21_)  &  n89 ) | ( (~ PV84_4_)  &  n409 ) | ( n89  &  n409 ) ;
 assign n150 = ( (~ PV47_25_)  &  n152  &  n153 ) | ( n100  &  n152  &  n153 ) ;
 assign n157 = ( (~ PV47_27_)  &  n102 ) | ( n102  &  n408 ) ;
 assign n158 = ( (~ PV84_3_)  &  (~ PV47_20_) ) | ( (~ PV47_20_)  &  n89 ) | ( (~ PV84_3_)  &  n409 ) | ( n89  &  n409 ) ;
 assign n155 = ( (~ PV47_24_)  &  n157  &  n158 ) | ( n100  &  n157  &  n158 ) ;
 assign n162 = ( (~ PV47_26_)  &  n102 ) | ( n102  &  n408 ) ;
 assign n163 = ( (~ PV84_2_)  &  (~ PV47_19_) ) | ( (~ PV47_19_)  &  n89 ) | ( (~ PV84_2_)  &  n409 ) | ( n89  &  n409 ) ;
 assign n160 = ( (~ PV47_23_)  &  n162  &  n163 ) | ( n100  &  n162  &  n163 ) ;
 assign n167 = ( (~ PV47_25_)  &  n102 ) | ( n102  &  n408 ) ;
 assign n168 = ( (~ PV84_1_)  &  (~ PV47_18_) ) | ( (~ PV47_18_)  &  n89 ) | ( (~ PV84_1_)  &  n409 ) | ( n89  &  n409 ) ;
 assign n165 = ( (~ PV47_22_)  &  n167  &  n168 ) | ( n100  &  n167  &  n168 ) ;
 assign n172 = ( (~ PV47_24_)  &  n102 ) | ( n102  &  n408 ) ;
 assign n173 = ( (~ PV84_0_)  &  (~ PV47_17_) ) | ( (~ PV47_17_)  &  n89 ) | ( (~ PV84_0_)  &  n409 ) | ( n89  &  n409 ) ;
 assign n170 = ( (~ PV47_21_)  &  n172  &  n173 ) | ( n100  &  n172  &  n173 ) ;
 assign n177 = ( PV133_2_ ) | ( n213 ) ;
 assign n176 = ( PV133_5_ ) | ( n411 ) ;
 assign n175 = ( (~ PV133_10_)  &  PV133_2_  &  n177 ) | ( (~ PV133_10_)  &  n177  &  n176 ) ;
 assign n179 = ( (~ PV116_14_)  &  n451 ) | ( (~ n404)  &  n451 ) ;
 assign n181 = ( (~ PV116_13_)  &  n451 ) | ( (~ n404)  &  n451 ) ;
 assign n183 = ( (~ PV116_12_)  &  n451 ) | ( (~ n404)  &  n451 ) ;
 assign n185 = ( (~ PV116_11_)  &  n451 ) | ( (~ n404)  &  n451 ) ;
 assign n187 = ( (~ PV116_10_)  &  n451 ) | ( (~ n404)  &  n451 ) ;
 assign n189 = ( (~ PV116_9_)  &  n451 ) | ( (~ n404)  &  n451 ) ;
 assign n191 = ( (~ PV116_8_)  &  n451 ) | ( (~ n404)  &  n451 ) ;
 assign n193 = ( (~ PV116_7_)  &  n451 ) | ( (~ n404)  &  n451 ) ;
 assign n195 = ( (~ PV116_6_)  &  n451 ) | ( (~ n404)  &  n451 ) ;
 assign n197 = ( (~ PV116_5_)  &  n451 ) | ( (~ n404)  &  n451 ) ;
 assign n199 = ( (~ PV116_4_)  &  n451 ) | ( (~ n404)  &  n451 ) ;
 assign n201 = ( (~ PV116_3_)  &  n451 ) | ( (~ n404)  &  n451 ) ;
 assign n203 = ( (~ PV116_2_)  &  n451 ) | ( (~ n404)  &  n451 ) ;
 assign n205 = ( (~ PV116_1_)  &  n451 ) | ( (~ n404)  &  n451 ) ;
 assign n207 = ( (~ PV116_0_)  &  n451 ) | ( (~ n404)  &  n451 ) ;
 assign n208 = ( (~ PV133_10_)  &  PV133_9_ ) | ( PV133_9_  &  (~ PV122_0_) ) | ( (~ PV133_10_)  &  n94 ) | ( (~ PV122_0_)  &  n94 ) ;
 assign n210 = ( PV133_10_  &  (~ PV84_0_) ) ;
 assign n212 = ( PV133_10_ ) | ( n412 ) ;
 assign n213 = ( PV133_1_ ) | ( n412 ) ;
 assign n211 = ( PV133_2_  &  PV133_10_ ) | ( n212  &  PV133_10_ ) | ( PV133_2_  &  n213 ) | ( n212  &  n213 ) ;
 assign n216 = ( PV133_1_ ) | ( n215 ) ;
 assign n215 = ( PV133_7_ ) | ( PV133_10_ ) | ( PV133_9_ ) ;
 assign n214 = ( n216  &  PV133_2_ ) | ( n216  &  n215 ) ;
 assign n219 = ( PV133_10_ ) | ( PV133_9_ ) | ( (~ PV133_8_) ) ;
 assign n217 = ( PV52_0_  &  n219  &  (~ n485) ) | ( n214  &  n219  &  (~ n485) ) ;
 assign n221 = ( (~ PV133_10_)  &  n5  &  n418 ) ;
 assign n220 = ( (~ PV47_2_)  &  (~ PV15_1_) ) | ( (~ PV15_1_)  &  n89 ) | ( (~ PV47_2_)  &  n409 ) | ( n89  &  n409 ) ;
 assign n224 = ( (~ PV116_1_)  &  n452  &  (~ n486) ) | ( (~ n404)  &  n452  &  (~ n486) ) ;
 assign n223 = ( (~ PV47_1_)  &  (~ PV15_0_) ) | ( (~ PV15_0_)  &  n89 ) | ( (~ PV47_1_)  &  n409 ) | ( n89  &  n409 ) ;
 assign n225 = ( (~ PV84_8_)  &  n102 ) | ( n102  &  n100 ) ;
 assign n229 = ( (~ PV47_0_)  &  (~ PV15_7_) ) | ( (~ PV15_7_)  &  n408 ) | ( (~ PV47_0_)  &  n409 ) | ( n408  &  n409 ) ;
 assign n227 = ( (~ PV47_8_)  &  n225  &  n229 ) | ( n89  &  n225  &  n229 ) ;
 assign n230 = ( n73  &  n257 ) ;
 assign n231 = ( (~ PV84_7_)  &  n102 ) | ( n102  &  n100 ) ;
 assign n234 = ( (~ PV116_7_) ) | ( (~ n404) ) ;
 assign n233 = ( (~ PV47_7_)  &  (~ PV15_6_) ) | ( (~ PV15_6_)  &  n89 ) | ( (~ PV47_7_)  &  n409 ) | ( n89  &  n409 ) ;
 assign n235 = ( (~ PV84_6_)  &  n102 ) | ( n102  &  n100 ) ;
 assign n238 = ( (~ PV116_6_) ) | ( (~ n404) ) ;
 assign n237 = ( (~ PV47_6_)  &  (~ PV15_5_) ) | ( (~ PV15_5_)  &  n89 ) | ( (~ PV47_6_)  &  n409 ) | ( n89  &  n409 ) ;
 assign n239 = ( (~ PV84_5_)  &  n102 ) | ( n102  &  n100 ) ;
 assign n242 = ( (~ PV116_5_) ) | ( (~ n404) ) ;
 assign n241 = ( (~ PV47_5_)  &  (~ PV15_4_) ) | ( (~ PV15_4_)  &  n89 ) | ( (~ PV47_5_)  &  n409 ) | ( n89  &  n409 ) ;
 assign n243 = ( (~ PV84_4_)  &  n102 ) | ( n102  &  n100 ) ;
 assign n246 = ( (~ PV116_4_) ) | ( (~ n404) ) ;
 assign n245 = ( (~ PV47_4_)  &  (~ PV15_3_) ) | ( (~ PV15_3_)  &  n89 ) | ( (~ PV47_4_)  &  n409 ) | ( n89  &  n409 ) ;
 assign n247 = ( (~ PV84_3_)  &  n102 ) | ( n102  &  n100 ) ;
 assign n250 = ( (~ PV116_3_) ) | ( (~ n404) ) ;
 assign n249 = ( (~ PV47_3_)  &  (~ PV15_2_) ) | ( (~ PV15_2_)  &  n89 ) | ( (~ PV47_3_)  &  n409 ) | ( n89  &  n409 ) ;
 assign n251 = ( (~ PV84_9_)  &  n102 ) | ( n102  &  n100 ) ;
 assign n255 = ( (~ PV47_1_)  &  (~ PV15_8_) ) | ( (~ PV15_8_)  &  n408 ) | ( (~ PV47_1_)  &  n409 ) | ( n408  &  n409 ) ;
 assign n253 = ( (~ PV47_9_)  &  n251  &  n255 ) | ( n89  &  n251  &  n255 ) ;
 assign n257 = ( (~ PV133_10_)  &  n412 ) ;
 assign n256 = ( n257  &  n7 ) ;
 assign n258 = ( (~ PV84_11_)  &  n102 ) | ( n102  &  n100 ) ;
 assign n262 = ( (~ PV47_3_)  &  (~ PV15_10_) ) | ( (~ PV15_10_)  &  n408 ) | ( (~ PV47_3_)  &  n409 ) | ( n408  &  n409 ) ;
 assign n260 = ( (~ PV47_11_)  &  n258  &  n262 ) | ( n89  &  n258  &  n262 ) ;
 assign n263 = ( (~ PV84_10_)  &  n102 ) | ( n102  &  n100 ) ;
 assign n267 = ( (~ PV47_2_)  &  (~ PV15_9_) ) | ( (~ PV15_9_)  &  n408 ) | ( (~ PV47_2_)  &  n409 ) | ( n408  &  n409 ) ;
 assign n265 = ( (~ PV47_10_)  &  n263  &  n267 ) | ( n89  &  n263  &  n267 ) ;
 assign n270 = ( (~ PV47_4_)  &  n102 ) | ( n102  &  n408 ) ;
 assign n271 = ( (~ PV47_12_)  &  (~ PV15_11_) ) | ( (~ PV15_11_)  &  n89 ) | ( (~ PV47_12_)  &  n409 ) | ( n89  &  n409 ) ;
 assign n268 = ( (~ PV47_1_)  &  n270  &  n271 ) | ( n100  &  n270  &  n271 ) ;
 assign n273 = ( (~ PV133_3_) ) | ( n7 ) ;
 assign n272 = ( n273  &  n257  &  PV133_2_ ) | ( n273  &  n257  &  n73 ) ;
 assign n275 = ( (~ PV116_12_)  &  (~ PV84_12_) ) | ( (~ PV84_12_)  &  (~ n404) ) | ( (~ PV116_12_)  &  n437 ) | ( (~ n404)  &  n437 ) ;
 assign n274 = ( PV133_1_ ) | ( n7 ) ;
 assign n279 = ( (~ PV116_15_)  &  (~ PV84_15_) ) | ( (~ PV84_15_)  &  (~ n404) ) | ( (~ PV116_15_)  &  n437 ) | ( (~ n404)  &  n437 ) ;
 assign n278 = ( n411  &  n272 ) ;
 assign n276 = ( (~ PV47_15_)  &  (~ PV15_14_) ) | ( (~ PV15_14_)  &  n89 ) | ( (~ PV47_15_)  &  n409 ) | ( n89  &  n409 ) ;
 assign n277 = ( (~ PV47_4_)  &  n102  &  n454 ) | ( n102  &  n100  &  n454 ) ;
 assign n282 = ( (~ PV116_14_)  &  (~ PV84_14_) ) | ( (~ PV84_14_)  &  (~ n404) ) | ( (~ PV116_14_)  &  n437 ) | ( (~ n404)  &  n437 ) ;
 assign n280 = ( (~ PV47_14_)  &  (~ PV15_13_) ) | ( (~ PV15_13_)  &  n89 ) | ( (~ PV47_14_)  &  n409 ) | ( n89  &  n409 ) ;
 assign n281 = ( (~ PV47_3_)  &  n102  &  n455 ) | ( n102  &  n100  &  n455 ) ;
 assign n285 = ( (~ PV116_13_)  &  (~ PV84_13_) ) | ( (~ PV84_13_)  &  (~ n404) ) | ( (~ PV116_13_)  &  n437 ) | ( (~ n404)  &  n437 ) ;
 assign n283 = ( (~ PV47_13_)  &  (~ PV15_12_) ) | ( (~ PV15_12_)  &  n89 ) | ( (~ PV47_13_)  &  n409 ) | ( n89  &  n409 ) ;
 assign n284 = ( (~ PV47_2_)  &  n102  &  n456 ) | ( n102  &  n100  &  n456 ) ;
 assign n286 = ( n278  &  PV133_2_ ) | ( n278  &  n274 ) ;
 assign n289 = ( (~ PV116_16_)  &  (~ PV84_16_) ) | ( (~ PV84_16_)  &  (~ n404) ) | ( (~ PV116_16_)  &  n437 ) | ( (~ n404)  &  n437 ) ;
 assign n287 = ( (~ PV47_16_)  &  (~ PV47_1_) ) | ( (~ PV47_1_)  &  n89 ) | ( (~ PV47_16_)  &  n409 ) | ( n89  &  n409 ) ;
 assign n288 = ( (~ PV47_5_)  &  n102  &  n457 ) | ( n102  &  n100  &  n457 ) ;
 assign n292 = ( (~ PV116_31_)  &  (~ PV84_31_) ) | ( (~ PV84_31_)  &  (~ n404) ) | ( (~ PV116_31_)  &  n437 ) | ( (~ n404)  &  n437 ) ;
 assign n290 = ( (~ PV47_31_)  &  (~ PV47_16_) ) | ( (~ PV47_16_)  &  n89 ) | ( (~ PV47_31_)  &  n409 ) | ( n89  &  n409 ) ;
 assign n291 = ( (~ PV47_20_)  &  n102  &  n458 ) | ( n102  &  n100  &  n458 ) ;
 assign n295 = ( (~ PV116_30_)  &  (~ PV84_30_) ) | ( (~ PV84_30_)  &  (~ n404) ) | ( (~ PV116_30_)  &  n437 ) | ( (~ n404)  &  n437 ) ;
 assign n293 = ( (~ PV47_30_)  &  (~ PV47_15_) ) | ( (~ PV47_15_)  &  n89 ) | ( (~ PV47_30_)  &  n409 ) | ( n89  &  n409 ) ;
 assign n294 = ( (~ PV47_19_)  &  n102  &  n459 ) | ( n102  &  n100  &  n459 ) ;
 assign n298 = ( (~ PV116_29_)  &  (~ PV84_29_) ) | ( (~ PV84_29_)  &  (~ n404) ) | ( (~ PV116_29_)  &  n437 ) | ( (~ n404)  &  n437 ) ;
 assign n296 = ( (~ PV47_29_)  &  (~ PV47_14_) ) | ( (~ PV47_14_)  &  n89 ) | ( (~ PV47_29_)  &  n409 ) | ( n89  &  n409 ) ;
 assign n297 = ( (~ PV47_18_)  &  n102  &  n460 ) | ( n102  &  n100  &  n460 ) ;
 assign n301 = ( (~ PV116_28_)  &  (~ PV84_28_) ) | ( (~ PV84_28_)  &  (~ n404) ) | ( (~ PV116_28_)  &  n437 ) | ( (~ n404)  &  n437 ) ;
 assign n299 = ( (~ PV47_28_)  &  (~ PV47_13_) ) | ( (~ PV47_13_)  &  n89 ) | ( (~ PV47_28_)  &  n409 ) | ( n89  &  n409 ) ;
 assign n300 = ( (~ PV47_17_)  &  n102  &  n461 ) | ( n102  &  n100  &  n461 ) ;
 assign n304 = ( (~ PV116_27_)  &  (~ PV84_27_) ) | ( (~ PV84_27_)  &  (~ n404) ) | ( (~ PV116_27_)  &  n437 ) | ( (~ n404)  &  n437 ) ;
 assign n302 = ( (~ PV47_27_)  &  (~ PV47_12_) ) | ( (~ PV47_12_)  &  n89 ) | ( (~ PV47_27_)  &  n409 ) | ( n89  &  n409 ) ;
 assign n303 = ( (~ PV47_16_)  &  n102  &  n462 ) | ( n102  &  n100  &  n462 ) ;
 assign n307 = ( (~ PV116_26_)  &  (~ PV84_26_) ) | ( (~ PV84_26_)  &  (~ n404) ) | ( (~ PV116_26_)  &  n437 ) | ( (~ n404)  &  n437 ) ;
 assign n305 = ( (~ PV47_26_)  &  (~ PV47_11_) ) | ( (~ PV47_11_)  &  n89 ) | ( (~ PV47_26_)  &  n409 ) | ( n89  &  n409 ) ;
 assign n306 = ( (~ PV47_15_)  &  n102  &  n463 ) | ( n102  &  n100  &  n463 ) ;
 assign n310 = ( (~ PV116_25_)  &  (~ PV84_25_) ) | ( (~ PV84_25_)  &  (~ n404) ) | ( (~ PV116_25_)  &  n437 ) | ( (~ n404)  &  n437 ) ;
 assign n308 = ( (~ PV47_25_)  &  (~ PV47_10_) ) | ( (~ PV47_10_)  &  n89 ) | ( (~ PV47_25_)  &  n409 ) | ( n89  &  n409 ) ;
 assign n309 = ( (~ PV47_14_)  &  n102  &  n464 ) | ( n102  &  n100  &  n464 ) ;
 assign n313 = ( (~ PV116_24_)  &  (~ PV84_24_) ) | ( (~ PV84_24_)  &  (~ n404) ) | ( (~ PV116_24_)  &  n437 ) | ( (~ n404)  &  n437 ) ;
 assign n311 = ( (~ PV47_24_)  &  (~ PV47_9_) ) | ( (~ PV47_9_)  &  n89 ) | ( (~ PV47_24_)  &  n409 ) | ( n89  &  n409 ) ;
 assign n312 = ( (~ PV47_13_)  &  n102  &  n465 ) | ( n102  &  n100  &  n465 ) ;
 assign n316 = ( (~ PV116_23_)  &  (~ PV84_23_) ) | ( (~ PV84_23_)  &  (~ n404) ) | ( (~ PV116_23_)  &  n437 ) | ( (~ n404)  &  n437 ) ;
 assign n314 = ( (~ PV47_23_)  &  (~ PV47_8_) ) | ( (~ PV47_8_)  &  n89 ) | ( (~ PV47_23_)  &  n409 ) | ( n89  &  n409 ) ;
 assign n315 = ( (~ PV47_12_)  &  n102  &  n466 ) | ( n102  &  n100  &  n466 ) ;
 assign n319 = ( (~ PV116_22_)  &  (~ PV84_22_) ) | ( (~ PV84_22_)  &  (~ n404) ) | ( (~ PV116_22_)  &  n437 ) | ( (~ n404)  &  n437 ) ;
 assign n317 = ( (~ PV47_22_)  &  (~ PV47_7_) ) | ( (~ PV47_7_)  &  n89 ) | ( (~ PV47_22_)  &  n409 ) | ( n89  &  n409 ) ;
 assign n318 = ( (~ PV47_11_)  &  n102  &  n467 ) | ( n102  &  n100  &  n467 ) ;
 assign n322 = ( (~ PV116_21_)  &  (~ PV84_21_) ) | ( (~ PV84_21_)  &  (~ n404) ) | ( (~ PV116_21_)  &  n437 ) | ( (~ n404)  &  n437 ) ;
 assign n320 = ( (~ PV47_21_)  &  (~ PV47_6_) ) | ( (~ PV47_6_)  &  n89 ) | ( (~ PV47_21_)  &  n409 ) | ( n89  &  n409 ) ;
 assign n321 = ( (~ PV47_10_)  &  n102  &  n468 ) | ( n102  &  n100  &  n468 ) ;
 assign n325 = ( (~ PV116_20_)  &  (~ PV84_20_) ) | ( (~ PV84_20_)  &  (~ n404) ) | ( (~ PV116_20_)  &  n437 ) | ( (~ n404)  &  n437 ) ;
 assign n323 = ( (~ PV47_20_)  &  (~ PV47_5_) ) | ( (~ PV47_5_)  &  n89 ) | ( (~ PV47_20_)  &  n409 ) | ( n89  &  n409 ) ;
 assign n324 = ( (~ PV47_9_)  &  n102  &  n469 ) | ( n102  &  n100  &  n469 ) ;
 assign n328 = ( (~ PV116_19_)  &  (~ PV84_19_) ) | ( (~ PV84_19_)  &  (~ n404) ) | ( (~ PV116_19_)  &  n437 ) | ( (~ n404)  &  n437 ) ;
 assign n326 = ( (~ PV47_19_)  &  (~ PV47_4_) ) | ( (~ PV47_4_)  &  n89 ) | ( (~ PV47_19_)  &  n409 ) | ( n89  &  n409 ) ;
 assign n327 = ( (~ PV47_8_)  &  n102  &  n470 ) | ( n102  &  n100  &  n470 ) ;
 assign n331 = ( (~ PV116_18_)  &  (~ PV84_18_) ) | ( (~ PV84_18_)  &  (~ n404) ) | ( (~ PV116_18_)  &  n437 ) | ( (~ n404)  &  n437 ) ;
 assign n329 = ( (~ PV47_18_)  &  (~ PV47_3_) ) | ( (~ PV47_3_)  &  n89 ) | ( (~ PV47_18_)  &  n409 ) | ( n89  &  n409 ) ;
 assign n330 = ( (~ PV47_7_)  &  n102  &  n471 ) | ( n102  &  n100  &  n471 ) ;
 assign n334 = ( (~ PV116_17_)  &  (~ PV84_17_) ) | ( (~ PV84_17_)  &  (~ n404) ) | ( (~ PV116_17_)  &  n437 ) | ( (~ n404)  &  n437 ) ;
 assign n332 = ( (~ PV47_17_)  &  (~ PV47_2_) ) | ( (~ PV47_2_)  &  n89 ) | ( (~ PV47_17_)  &  n409 ) | ( n89  &  n409 ) ;
 assign n333 = ( (~ PV47_6_)  &  n102  &  n472 ) | ( n102  &  n100  &  n472 ) ;
 assign n336 = ( (~ PV84_23_)  &  n102 ) | ( n102  &  n408 ) ;
 assign n337 = ( (~ PV84_31_)  &  (~ PV84_16_) ) | ( (~ PV84_16_)  &  n89 ) | ( (~ PV84_31_)  &  n409 ) | ( n89  &  n409 ) ;
 assign n335 = ( (~ PV84_20_)  &  n336  &  n337 ) | ( n100  &  n336  &  n337 ) ;
 assign n340 = ( (~ PV84_22_)  &  n102 ) | ( n102  &  n408 ) ;
 assign n341 = ( (~ PV84_30_)  &  (~ PV84_15_) ) | ( (~ PV84_15_)  &  n89 ) | ( (~ PV84_30_)  &  n409 ) | ( n89  &  n409 ) ;
 assign n339 = ( (~ PV84_19_)  &  n340  &  n341 ) | ( n100  &  n340  &  n341 ) ;
 assign n344 = ( (~ PV84_21_)  &  n102 ) | ( n102  &  n408 ) ;
 assign n345 = ( (~ PV84_29_)  &  (~ PV84_14_) ) | ( (~ PV84_14_)  &  n89 ) | ( (~ PV84_29_)  &  n409 ) | ( n89  &  n409 ) ;
 assign n343 = ( (~ PV84_18_)  &  n344  &  n345 ) | ( n100  &  n344  &  n345 ) ;
 assign n348 = ( (~ PV84_20_)  &  n102 ) | ( n102  &  n408 ) ;
 assign n349 = ( (~ PV84_28_)  &  (~ PV84_13_) ) | ( (~ PV84_13_)  &  n89 ) | ( (~ PV84_28_)  &  n409 ) | ( n89  &  n409 ) ;
 assign n347 = ( (~ PV84_17_)  &  n348  &  n349 ) | ( n100  &  n348  &  n349 ) ;
 assign n353 = ( (~ PV84_19_)  &  n102 ) | ( n102  &  n408 ) ;
 assign n354 = ( (~ PV84_27_)  &  (~ PV84_12_) ) | ( (~ PV84_12_)  &  n89 ) | ( (~ PV84_27_)  &  n409 ) | ( n89  &  n409 ) ;
 assign n351 = ( (~ PV84_16_)  &  n353  &  n354 ) | ( n100  &  n353  &  n354 ) ;
 assign n358 = ( (~ PV84_18_)  &  n102 ) | ( n102  &  n408 ) ;
 assign n359 = ( (~ PV84_26_)  &  (~ PV84_11_) ) | ( (~ PV84_11_)  &  n89 ) | ( (~ PV84_26_)  &  n409 ) | ( n89  &  n409 ) ;
 assign n356 = ( (~ PV84_15_)  &  n358  &  n359 ) | ( n100  &  n358  &  n359 ) ;
 assign n363 = ( (~ PV84_17_)  &  n102 ) | ( n102  &  n408 ) ;
 assign n364 = ( (~ PV84_25_)  &  (~ PV84_10_) ) | ( (~ PV84_10_)  &  n89 ) | ( (~ PV84_25_)  &  n409 ) | ( n89  &  n409 ) ;
 assign n361 = ( (~ PV84_14_)  &  n363  &  n364 ) | ( n100  &  n363  &  n364 ) ;
 assign n367 = ( (~ PV84_16_)  &  n102 ) | ( n102  &  n408 ) ;
 assign n368 = ( (~ PV84_24_)  &  (~ PV84_9_) ) | ( (~ PV84_9_)  &  n89 ) | ( (~ PV84_24_)  &  n409 ) | ( n89  &  n409 ) ;
 assign n366 = ( (~ PV84_13_)  &  n367  &  n368 ) | ( n100  &  n367  &  n368 ) ;
 assign n371 = ( (~ PV84_15_)  &  n102 ) | ( n102  &  n408 ) ;
 assign n372 = ( (~ PV84_23_)  &  (~ PV84_8_) ) | ( (~ PV84_8_)  &  n89 ) | ( (~ PV84_23_)  &  n409 ) | ( n89  &  n409 ) ;
 assign n370 = ( (~ PV84_12_)  &  n371  &  n372 ) | ( n100  &  n371  &  n372 ) ;
 assign n375 = ( (~ PV84_14_)  &  (~ PV84_7_) ) | ( (~ PV84_7_)  &  n408 ) | ( (~ PV84_14_)  &  n409 ) | ( n408  &  n409 ) ;
 assign n374 = ( (~ PV84_22_)  &  n258  &  n375 ) | ( n89  &  n258  &  n375 ) ;
 assign n378 = ( (~ PV84_13_)  &  (~ PV84_6_) ) | ( (~ PV84_6_)  &  n408 ) | ( (~ PV84_13_)  &  n409 ) | ( n408  &  n409 ) ;
 assign n377 = ( (~ PV84_21_)  &  n263  &  n378 ) | ( n89  &  n263  &  n378 ) ;
 assign n381 = ( (~ PV84_12_)  &  (~ PV84_5_) ) | ( (~ PV84_5_)  &  n408 ) | ( (~ PV84_12_)  &  n409 ) | ( n408  &  n409 ) ;
 assign n380 = ( (~ PV84_20_)  &  n251  &  n381 ) | ( n89  &  n251  &  n381 ) ;
 assign n384 = ( (~ PV84_11_)  &  (~ PV84_4_) ) | ( (~ PV84_4_)  &  n408 ) | ( (~ PV84_11_)  &  n409 ) | ( n408  &  n409 ) ;
 assign n383 = ( (~ PV84_19_)  &  n225  &  n384 ) | ( n89  &  n225  &  n384 ) ;
 assign n387 = ( (~ PV84_10_)  &  (~ PV84_3_) ) | ( (~ PV84_3_)  &  n408 ) | ( (~ PV84_10_)  &  n409 ) | ( n408  &  n409 ) ;
 assign n386 = ( (~ PV84_18_)  &  n231  &  n387 ) | ( n89  &  n231  &  n387 ) ;
 assign n390 = ( (~ PV84_9_)  &  (~ PV84_2_) ) | ( (~ PV84_2_)  &  n408 ) | ( (~ PV84_9_)  &  n409 ) | ( n408  &  n409 ) ;
 assign n389 = ( (~ PV84_17_)  &  n235  &  n390 ) | ( n89  &  n235  &  n390 ) ;
 assign n393 = ( (~ PV84_8_)  &  (~ PV84_1_) ) | ( (~ PV84_1_)  &  n408 ) | ( (~ PV84_8_)  &  n409 ) | ( n408  &  n409 ) ;
 assign n392 = ( (~ PV84_16_)  &  n239  &  n393 ) | ( n89  &  n239  &  n393 ) ;
 assign n396 = ( (~ PV84_7_)  &  (~ PV84_0_) ) | ( (~ PV84_0_)  &  n408 ) | ( (~ PV84_7_)  &  n409 ) | ( n408  &  n409 ) ;
 assign n395 = ( (~ PV84_15_)  &  n243  &  n396 ) | ( n89  &  n243  &  n396 ) ;
 assign n399 = ( (~ PV84_6_)  &  (~ PV47_31_) ) | ( (~ PV47_31_)  &  n408 ) | ( (~ PV84_6_)  &  n409 ) | ( n408  &  n409 ) ;
 assign n398 = ( (~ PV84_14_)  &  n247  &  n399 ) | ( n89  &  n247  &  n399 ) ;
 assign n402 = ( PV133_9_ ) | ( (~ PV133_5_) ) | ( PV133_1_ ) ;
 assign n401 = ( n402 ) | ( PV118_0_ ) ;
 assign n403 = ( n402 ) | ( PV133_0_ ) ;
 assign n404 = ( (~ PV133_10_)  &  PV133_9_ ) ;
 assign n405 = ( (~ n89) ) | ( (~ n96) ) ;
 assign n408 = ( (~ n89) ) | ( n96 ) ;
 assign n409 = ( (~ n91) ) | ( n405 ) ;
 assign n411 = ( PV133_1_ ) | ( n73 ) ;
 assign n412 = ( PV133_9_ ) | ( (~ PV133_7_) ) ;
 assign n418 = ( PV133_8_ ) | ( n412 ) ;
 assign n437 = ( n6 ) | ( n215 ) | ( PV133_3_ ) | ( PV133_4_ ) ;
 assign n447 = ( (~ PV133_10_)  &  n94  &  (~ n404) ) | ( PV119_0_  &  n94  &  (~ n404) ) ;
 assign n448 = ( (~ PV121_16_)  &  (~ n447) ) | ( (~ n447)  &  n474 ) | ( (~ PV121_16_)  &  (~ n474) ) ;
 assign n449 = ( (~ PV121_17_)  &  n208 ) | ( n208  &  n212 ) | ( (~ PV121_17_)  &  (~ n212) ) ;
 assign n450 = ( (~ PV48_0_)  &  (~ n211) ) | ( (~ PV48_0_)  &  n481 ) | ( n211  &  n481 ) ;
 assign n451 = ( (~ PV133_5_) ) | ( PV133_2_ ) | ( PV118_1_ ) | ( PV118_0_ ) | ( n216 ) ;
 assign n452 = ( (~ PV51_0_) ) | ( n214 ) | ( (~ n219) ) ;
 assign n454 = ( (~ PV47_7_) ) | ( n408 ) ;
 assign n455 = ( (~ PV47_6_) ) | ( n408 ) ;
 assign n456 = ( (~ PV47_5_) ) | ( n408 ) ;
 assign n457 = ( (~ PV47_8_) ) | ( n408 ) ;
 assign n458 = ( (~ PV47_23_) ) | ( n408 ) ;
 assign n459 = ( (~ PV47_22_) ) | ( n408 ) ;
 assign n460 = ( (~ PV47_21_) ) | ( n408 ) ;
 assign n461 = ( (~ PV47_20_) ) | ( n408 ) ;
 assign n462 = ( (~ PV47_19_) ) | ( n408 ) ;
 assign n463 = ( (~ PV47_18_) ) | ( n408 ) ;
 assign n464 = ( (~ PV47_17_) ) | ( n408 ) ;
 assign n465 = ( (~ PV47_16_) ) | ( n408 ) ;
 assign n466 = ( (~ PV47_15_) ) | ( n408 ) ;
 assign n467 = ( (~ PV47_14_) ) | ( n408 ) ;
 assign n468 = ( (~ PV47_13_) ) | ( n408 ) ;
 assign n469 = ( (~ PV47_12_) ) | ( n408 ) ;
 assign n470 = ( (~ PV47_11_) ) | ( n408 ) ;
 assign n471 = ( (~ PV47_10_) ) | ( n408 ) ;
 assign n472 = ( (~ PV47_9_) ) | ( n408 ) ;
 assign n474 = ( PV133_10_ ) | ( n418 ) ;
 assign n479 = ( (~ PV116_0_)  &  n210 ) | ( (~ PV116_0_)  &  n404 ) | ( n210  &  (~ n404) ) ;
 assign n481 = ( (~ PV49_0_)  &  (~ n215) ) | ( (~ PV49_0_)  &  n479 ) | ( n215  &  n479 ) ;
 assign n485 = ( (~ PV116_2_)  &  n214 ) | ( n214  &  (~ n404) ) ;
 assign n486 = ( PV50_0_  &  (~ n219) ) ;


endmodule

