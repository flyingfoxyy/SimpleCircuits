module alu4_mapped (
	i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, 
	i_4_, i_12_, i_1_, i_11_, i_2_, i_0_, o_1_, o_2_, o_0_, o_7_, 
	o_5_, o_6_, o_3_, o_4_);

input i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_, i_1_, i_11_, i_2_, i_0_;

output o_1_, o_2_, o_0_, o_7_, o_5_, o_6_, o_3_, o_4_;

wire n_n860, n_n861, wire1852, wire6485, n_n874, wire1789, wire6528, wire6530, wire6536, wire6537, wire6538, n_n1221, n_n1222, wire6827, wire6828, wire6937, wire6938, wire6949, wire6950, n_n1185, wire6975, wire7001, wire7076, n_n955, wire7337, wire7339, n_n637, wire1867, wire1869, wire6474, wire6475, wire747, wire1861, wire6479, wire8, wire21, wire23, wire414, wire648, wire1841, wire6491, n_n877, wire1832, wire1833, wire6495, wire6496, n_n876, wire1823, wire1825, wire6500, wire6501, n_n878, n_n879, n_n881, wire6520, wire18, wire55, wire126, wire278, wire283, wire327, wire343, wire348, wire386, wire284, wire483, wire6615, wire6616, n_n1240, wire344, wire502, wire6594, wire6627, n_n1241, n_n1248, n_n1229, wire1547, wire6704, wire1535, wire1537, wire6715, n_n1236, n_n1261, n_n1231, n_n1233, wire6791, wire1375, wire1376, wire6834, n_n1121, wire1362, wire1363, wire1366, wire6840, n_n1120, wire1186, wire1195, wire6941, wire6946, n_n1108, wire14, wire6956, n_n1189, wire1096, wire1097, wire6997, n_n1187, n_n658, n_n741, n_n566, n_n764, n_n701, wire323, wire325, wire326, wire947, wire7088, n_n970, wire937, wire20, wire578, wire925, wire7102, wire881, wire882, wire884, n_n984, n_n983, wire7167, wire7168, n_n965, wire7232, wire40, wire50, wire52, wire7329, n_n957, n_n816, n_n853, n_n779, n_n795, wire17, wire33, wire35, wire37, n_n835, wire68, wire288, wire313, wire322, wire336, wire420, n_n833, n_n538, n_n850, n_n498, n_n838, n_n748, n_n725, wire341, n_n665, wire427, wire1756, wire6555, wire425, wire6557, n_n609, wire1746, wire1744, n_n623, n_n619, wire376, wire436, wire435, n_n830, n_n633, n_n631, wire434, n_n716, n_n849, n_n36, n_n685, wire309, wire439, wire438, n_n545, n_n675, wire29, wire289, n_n792, wire295, wire6837, wire443, wire269, wire442, n_n570, n_n787, n_n769, n_n819, n_n273, wire381, wire12, wire377, n_n847, wire27, n_n581, wire264, n_n638, wire15, n_n814, n_n541, wire28, n_n746, wire333, n_n453, n_n761, n_n421, n_n415, n_n369, wire25, n_n358, n_n412, wire279, n_n773, n_n844, wire13, n_n639, wire286, n_n185, n_n432, n_n826, n_n183, wire96, n_n818, n_n153, n_n316, n_n197, n_n843, n_n699, wire293, n_n678, n_n671, wire26, n_n176, n_n712, n_n751, wire265, n_n719, wire31, n_n687, wire34, n_n827, wire267, n_n683, n_n275, n_n35, wire69, wire370, wire70, n_n791, wire106, wire6735, wire1652, wire1656, wire6633, wire454, n_n635, wire453, wire1647, wire1648, n_n752, wire307, n_n592, n_n832, n_n852, wire6587, n_n1243, wire388, wire42, wire6591, wire465, n_n598, n_n575, wire19, wire9, n_n672, n_n810, wire371, wire301, wire346, wire11, n_n653, n_n526, n_n534, n_n242, n_n656, n_n194, n_n346, n_n842, wire281, n_n755, n_n846, wire1503, wire1504, wire6745, n_n1258, n_n670, wire6669, wire113, n_n756, n_n550, n_n732, wire484, wire1679, wire1681, n_n729, wire482, wire487, wire486, wire485, wire6871, wire6872, wire6873, n_n1126, wire22, wire38, wire297, wire1293, wire1294, wire1295, wire1296, n_n1127, wire493, wire342, wire393, wire491, wire1283, wire6890, n_n1112, wire268, n_n274, n_n837, n_n240, wire330, n_n771, n_n606, n_n813, wire290, wire308, wire318, n_n768, wire6748, wire494, wire360, wire1637, wire1643, wire6640, wire497, wire1634, wire1635, n_n1250, wire294, wire296, wire503, wire1669, wire6624, wire277, wire501, wire272, wire298, wire311, wire363, wire1274, wire6893, wire6896, wire104, wire270, wire379, wire507, wire1263, wire6902, wire6905, wire181, wire364, wire512, wire516, wire513, n_n822, n_n840, n_n710, wire520, wire1629, wire1630, wire519, wire6644, wire518, n_n735, wire6642, wire517, wire1624, wire6651, n_n1256, wire525, wire524, wire523, wire6756, wire521, wire1490, wire6752, wire6759, wire350, wire529, wire16, wire533, wire536, n_n597, n_n651, wire1610, wire6658, n_n1255, wire405, wire546, wire1603, wire1605, wire545, wire544, wire543, wire571, wire6683, n_n1253, wire120, wire6678, wire6922, wire553, wire6921, wire552, wire1221, wire6926, n_n1128, wire30, wire352, wire7249, wire7250, wire557, wire338, wire562, wire561, wire560, wire558, wire176, wire7255, n_n1000, wire375, wire170, wire171, wire172, wire565, wire36, wire7257, wire564, n_n503, wire73, wire121, wire573, wire572, n_n1264, n_n1265, n_n851, wire574, n_n624, wire24, wire931, wire932, wire579, wire6848, wire584, wire1418, wire1419, wire583, wire410, wire1414, wire115, wire1400, wire1402, wire6814, n_n1234, wire591, wire594, wire593, wire123, wire276, wire291, wire354, wire7287, wire7288, wire596, n_n277, wire6807, wire1214, wire1215, wire1216, wire1217, wire604, wire606, wire1462, wire1463, wire1466, wire6766, wire292, wire340, wire359, wire6777, wire612, wire1132, wire1134, wire6978, wire6979, n_n1191, wire1154, wire6966, wire351, wire369, wire617, wire616, wire314, wire275, wire356, wire619, n_n612, wire626, wire628, wire633, wire632, wire7129, wire7127, wire638, wire7126, wire637, wire41, wire382, wire641, wire324, wire1064, wire7019, wire649, wire1848, wire1849, wire299, wire316, wire395, wire304, wire384, wire385, wire347, wire657, wire777, wire7185, wire655, wire772, wire773, n_n991, wire660, wire1814, wire6506, wire6507, wire287, wire1805, wire1806, wire1808, wire6512, wire668, wire667, wire7066, wire666, wire1074, wire7013, wire669, wire671, wire406, wire677, wire676, wire403, wire334, wire380, wire686, wire685, wire373, wire7191, n_n993, wire1012, wire7046, wire7047, wire1003, wire1005, wire7050, wire7051, wire696, wire397, wire701, wire7269, wire700, wire704, wire366, wire7275, wire703, wire706, wire707, wire7294, wire7295, wire7296, wire705, wire7178, wire708, wire785, wire718, wire717, wire719, wire7194, wire716, wire256, wire7196, wire762, wire857, wire7140, n_n981, wire836, wire7155, wire824, wire825, wire7161, wire726, wire725, wire724, wire7165, wire723, wire374, wire246, wire247, wire249, wire808, wire809, wire735, wire10, wire737, wire263, wire230, wire231, wire7219, wire736, wire7226, wire738, wire746, wire751, wire54, wire80, wire81, wire752, wire763, wire863, wire864, wire7132, wire7133, wire761, wire51, wire317, wire319, wire329, wire335, wire424, wire6549, wire6550, wire423, wire429, wire428, wire426, wire1740, wire1741, wire440, wire447, wire452, wire451, wire459, wire469, wire468, wire479, wire6622, wire6623, wire515, wire531, wire530, wire541, wire551, wire569, wire576, wire6803, wire615, wire622, wire636, wire635, wire644, wire643, wire646, wire653, wire7184, wire673, wire680, wire684, wire1794, wire683, wire7190, wire689, wire698, wire712, wire728, wire734, wire741, wire7136, wire7322, wire57, wire7325, wire59, wire60, wire7327, wire1202, wire1203, wire62, wire63, wire82, wire83, wire7312, wire64, wire84, wire7313, wire65, wire86, wire95, wire89, wire7304, wire103, wire107, wire112, wire7280, wire127, wire7282, wire128, wire136, wire129, wire130, wire144, wire145, wire139, wire141, wire142, wire143, wire7264, wire150, wire156, wire154, wire163, wire166, wire180, wire182, wire190, wire194, wire1408, wire1409, wire192, wire7235, wire198, wire200, wire207, wire201, wire7239, wire208, wire841, wire842, wire7223, wire212, wire213, wire222, wire7229, wire215, wire223, wire224, wire7215, wire225, wire7208, wire235, wire236, wire241, wire237, wire238, wire253, wire7199, wire245, wire7200, wire7203, wire255, wire6976, wire258, wire7188, wire362, wire768, wire769, wire7181, wire779, wire790, wire791, wire798, wire7175, wire800, wire802, wire801, wire814, wire7157, wire834, wire835, wire843, wire844, wire850, wire852, wire7146, wire845, wire7138, wire853, wire854, wire855, wire856, wire859, wire7134, wire7119, wire7121, wire7015, wire887, wire7122, wire891, wire895, wire905, wire7109, wire907, wire912, wire7110, wire7111, wire909, wire917, wire7094, wire934, wire7100, wire927, wire954, wire7084, wire7085, wire7086, wire948, wire957, wire958, wire7078, wire7080, wire961, wire7068, wire972, wire995, wire987, wire988, wire993, wire1009, wire1021, wire1026, wire1027, wire1023, wire1030, wire7042, wire7043, wire1024, wire1040, wire1041, wire7035, wire1033, wire1043, wire1044, wire1042, wire1047, wire7017, wire7018, wire1067, wire1082, wire1089, wire7004, wire7005, wire1083, wire1087, wire1092, wire1093, wire6994, wire1094, wire6996, wire1103, wire1115, wire1116, wire1117, wire1108, wire1119, wire1109, wire1110, wire1130, wire6983, wire1121, wire1122, wire1123, wire1133, wire1135, wire1152, wire6967, wire1139, wire1143, wire1160, wire1156, wire1162, wire1166, wire1171, wire1168, wire1173, wire1175, wire6959, wire1169, wire1180, wire1181, wire1182, wire1183, wire6945, wire1194, wire1348, wire1196, wire1200, wire1204, wire1213, wire6920, wire1218, wire1228, wire6925, wire1229, wire1230, wire1239, wire1234, wire1235, wire1245, wire1249, wire1250, wire1246, wire1252, wire6908, wire1247, wire1248, wire6897, wire1255, wire1266, wire1272, wire1267, wire1277, wire1279, wire1290, wire6887, wire6875, wire6876, wire1301, wire1302, wire6879, wire1297, wire1298, wire1299, wire1300, wire1307, wire1308, wire1314, wire6864, wire1321, wire1338, wire1339, wire1317, wire1324, wire1331, wire1326, wire1328, wire1329, wire1334, wire1336, wire1337, wire6852, wire1340, wire6853, wire1341, wire1346, wire1343, wire1361, wire6842, wire6843, wire1350, wire1351, wire1352, wire1353, wire6846, wire6835, wire1372, wire6838, wire1373, wire1383, wire6831, wire1377, wire1385, wire1393, wire1394, wire1388, wire1390, wire6816, wire1397, wire1406, wire6812, wire1403, wire6794, wire1410, wire6799, wire6785, wire1423, wire1432, wire1433, wire1425, wire6788, wire1436, wire6776, wire1437, wire1440, wire1441, wire1446, wire1447, wire1450, wire6770, wire6771, wire6772, wire6762, wire6763, wire1464, wire6764, wire1472, wire1474, wire1480, wire1481, wire1488, wire1493, wire6749, wire6750, wire1500, wire1501, wire1502, wire6719, wire1524, wire1525, wire1526, wire1527, wire1528, wire6725, wire1529, wire1530, wire1534, wire6714, wire6708, wire1552, wire1553, wire6698, wire1554, wire1562, wire6686, wire1563, wire6687, wire6688, wire1564, wire1565, wire1574, wire1575, wire1569, wire1571, wire1572, wire1587, wire1588, wire6670, wire1582, wire6672, wire1583, wire6674, wire6675, wire1585, wire1596, wire1611, wire1620, wire6647, wire6636, wire1639, wire1640, wire1644, wire6630, wire6631, wire6563, wire6632, wire1661, wire1663, wire1672, wire1673, wire1675, wire6595, wire1684, wire1685, wire6603, wire1686, wire6598, wire1689, wire1691, wire1704, wire1705, wire6588, wire1699, wire6589, wire6578, wire6579, wire1708, wire6582, wire1709, wire6584, wire6585, wire1720, wire1724, wire1725, wire1722, wire1726, wire6573, wire1729, wire1732, wire6558, wire6559, wire1748, wire1750, wire1763, wire1764, wire1767, wire1768, wire1765, wire1770, wire1776, wire1778, wire1779, wire1780, wire1781, wire1792, wire1803, wire1804, wire1796, wire6515, wire6516, wire1797, wire1798, wire6509, wire1810, wire6510, wire1820, wire1821, wire1816, wire1817, wire1829, wire6493, wire6494, wire1838, wire1839, wire1844, wire1845, wire1850, wire1856, wire1857, wire1853, wire1863, wire6478, wire6473, wire6488, wire6499, wire6504, wire6522, wire6523, wire6524, wire6526, wire6527, wire6554, wire6567, wire6593, wire6600, wire6605, wire6618, wire6620, wire6621, wire6628, wire6629, wire6637, wire6638, wire6643, wire6645, wire6653, wire6654, wire6660, wire6661, wire6665, wire6667, wire6673, wire6693, wire6712, wire6713, wire6730, wire6731, wire6757, wire6780, wire6787, wire6789, wire6806, wire6811, wire6850, wire6854, wire6858, wire6860, wire6865, wire6868, wire6869, wire6870, wire6884, wire6885, wire6886, wire6888, wire6894, wire6899, wire6900, wire6901, wire6904, wire6906, wire6911, wire6913, wire6914, wire6915, wire6916, wire6918, wire6919, wire6923, wire6924, wire6929, wire6930, wire6931, wire6934, wire6942, wire6944, wire6952, wire6958, wire6961, wire6964, wire6968, wire6969, wire6970, wire6972, wire6973, wire6982, wire6984, wire6985, wire6987, wire6991, wire6992, wire6995, wire6999, wire7003, wire7007, wire7008, wire7010, wire7011, wire7021, wire7022, wire7023, wire7024, wire7027, wire7028, wire7029, wire7030, wire7032, wire7033, wire7037, wire7040, wire7041, wire7057, wire7058, wire7059, wire7060, wire7062, wire7063, wire7070, wire7071, wire7074, wire7079, wire7082, wire7083, wire7092, wire7104, wire7105, wire7107, wire7108, wire7113, wire7114, wire7115, wire7117, wire7118, wire7130, wire7144, wire7149, wire7151, wire7163, wire7164, wire7174, wire7177, wire7182, wire7183, wire7202, wire7211, wire7214, wire7218, wire7222, wire7227, wire7228, wire7231, wire7237, wire7241, wire7246, wire7248, wire7251, wire7253, wire7254, wire7260, wire7261, wire7262, wire7263, wire7266, wire7267, wire7268, wire7271, wire7272, wire7273, wire7277, wire7278, wire7279, wire7286, wire7289, wire7292, wire7293, wire7297, wire7302, wire7303, wire7307, wire7308, wire7309, wire7310, wire7311, wire7314, wire7317, wire7318, wire7319, wire7321, wire7324, wire7326, wire7335, wire7336, _25, _41, _42, _52, _53, _64, _67, _68, _196, _197, _204, _221, _222, _267, _268, _274, _279, _284, _292, _296, _301, _310, _313, _314, _319, _372, _411, _412, _413, _414, _430, _431, _459, _520, _523, _524, _536, _537, _575, _629, _630, _666, _684, _685, _808, _810, _812, _813, _840, _844, _845, _847, _855, _856, _863, _864, _865, _870, _871, _872, _873, _875, _876, _880, _881, _893, _894, _897, _901, _930, _933, _934, _941, _948, _951, _952, _986, _987, _990, _991, _993, _1018, _1019, _1047, _1050, _1054, _1081, _1084, _1085, _1113, _1114, _1122, _8162, _8227, _8232, _8334, _8369, _8395, _8407, _8421, _8424, _8425, _8427, _8446, _8451, _8457, _8480, _8482, _8489, _8492, _8496, _8509, _8519, _8521, _8562, _8586, _8588, _8597, _8598, _8600, _8610, _8633, _8662, _8664, _8678, _8680, _8681, _8690, _8728, _8746, _8747, _8751, _8758, _8768, _8774, _8793, _8807, _8808, _8812, _8814, _8824, _8833, _8842, _8852, _8853, _8854, _8869, _8904, _8905, _8908, _8989, _9006, _9028, _9029, _9050, _9055, _9087, _9093, _9115, _9128, _9139, _9141, _9151, _9152, _9168, _9176, _9183, _9185, _9186, _9187, _9198, _9200, _9211, _9277, _9279, _9280, _9285, _9288, _9290, _9296, _9297, _9303, _9304, _9309, _9324, _9328, _9347, _9362, _9364, _9376, _9380, _9382, _9386, _9409, _9492, _9494, _9496, _9504, _9512, _9523, _9528, _9529, _9532, _9535, _9536, _9537, _9539, _9541, _9542, _9543, _9544, _9545, _9570, _9589, _9611, _9615, _9628, _9640, _9669, _9672, _9676, _9805, _9809, _9811, _9837, _9846, _9853, _9856, _9867, _9868, _9881, _9885;

assign o_1_ = ( n_n860 ) | ( n_n861 ) | ( wire1852 ) | ( wire6485 ) ;
 assign o_2_ = ( n_n874 ) | ( wire1789 ) | ( wire6528 ) | ( wire6530 ) ;
 assign o_0_ = ( wire6536 ) | ( wire6537 ) | ( wire6538 ) ;
 assign o_7_ = ( n_n1221 ) | ( n_n1222 ) | ( wire6827 ) | ( wire6828 ) ;
 assign o_5_ = ( wire6937 ) | ( wire6938 ) | ( wire6949 ) | ( wire6950 ) ;
 assign o_6_ = ( n_n1185 ) | ( wire6975 ) | ( wire7001 ) ;
 assign o_3_ = ( wire7040 ) | ( wire7063 ) | ( _9362 ) | ( _9386 ) ;
 assign o_4_ = ( n_n955 ) | ( wire7339 ) | ( _9885 ) ;
 assign n_n860 = ( wire1867 ) | ( wire1869 ) | ( wire6474 ) | ( wire6475 ) ;
 assign n_n861 = ( wire1861 ) | ( wire6479 ) | ( (~ i_3_)  &  wire747 ) ;
 assign wire1852 = ( (~ i_4_)  &  n_n609 ) | ( (~ i_4_)  &  wire1856 ) | ( (~ i_4_)  &  wire1857 ) ;
 assign wire6485 = ( wire1850 ) | ( wire1853 ) | ( wire21  &  wire414 ) ;
 assign n_n874 = ( n_n879 ) | ( n_n881 ) | ( wire6520 ) ;
 assign wire1789 = ( i_5_  &  wire1792 ) | ( i_5_  &  i_12_  &  wire683 ) ;
 assign wire6528 = ( wire6526 ) | ( wire6527 ) ;
 assign wire6530 = ( n_n877 ) | ( n_n876 ) | ( n_n878 ) ;
 assign wire6536 = ( wire126 ) | ( wire343 ) | ( wire1776 ) ;
 assign wire6537 = ( wire348 ) | ( wire386 ) | ( wire1778 ) | ( wire1779 ) ;
 assign wire6538 = ( wire1780 ) | ( wire1781 ) | ( wire278  &  wire327 ) ;
 assign n_n1221 = ( n_n1248 ) | ( n_n1229 ) | ( wire1547 ) | ( wire6704 ) ;
 assign n_n1222 = ( n_n1261 ) | ( n_n1231 ) | ( n_n1233 ) | ( wire6791 ) ;
 assign wire6827 = ( n_n1240 ) | ( n_n1241 ) | ( n_n1236 ) | ( _8774 ) ;
 assign wire6828 = ( wire6567 ) | ( wire6806 ) | ( _8905 ) | ( _8908 ) ;
 assign wire6937 = ( n_n1112 ) | ( wire6934 ) | ( n_n369  &  wire604 ) ;
 assign wire6938 = ( n_n1128 ) | ( wire6919 ) | ( _9050 ) ;
 assign wire6949 = ( n_n1108 ) | ( wire1350 ) | ( wire1353 ) | ( wire6850 ) ;
 assign wire6950 = ( n_n1121 ) | ( n_n1120 ) | ( wire6869 ) | ( wire6870 ) ;
 assign n_n1185 = ( _9187 ) | ( i_2_  &  wire6966 ) ;
 assign wire6975 = ( wire1143 ) | ( wire6969 ) | ( wire6972 ) | ( wire6973 ) ;
 assign wire7001 = ( n_n1187 ) | ( wire6991 ) | ( wire6992 ) | ( wire6999 ) ;
 assign wire7076 = ( wire972 ) | ( wire1083 ) | ( wire7008 ) | ( wire7074 ) ;
 assign n_n955 = ( n_n965 ) | ( _9535 ) | ( _9536 ) | ( _9537 ) ;
 assign wire7337 = ( n_n984 ) | ( n_n983 ) | ( _9570 ) | ( _9589 ) ;
 assign wire7339 = ( wire7318 ) | ( wire7319 ) | ( wire7321 ) | ( wire7336 ) ;
 assign n_n637 = ( i_13_  &  (~ i_11_) ) ;
 assign wire1867 = ( i_3_  &  wire319 ) | ( i_3_  &  n_n842  &  wire728 ) ;
 assign wire1869 = ( (~ i_8_)  &  wire369 ) ;
 assign wire6474 = ( wire23  &  wire370 ) | ( wire277  &  wire6473 ) ;
 assign wire6475 = ( (~ i_9_)  &  i_4_  &  wire313 ) | ( (~ i_9_)  &  i_4_  &  _8162 ) ;
 assign wire747 = ( i_13_  &  (~ i_12_)  &  (~ i_11_) ) | ( (~ i_13_)  &  i_4_  &  i_12_  &  i_11_ ) ;
 assign wire1861 = ( i_13_  &  wire1863 ) | ( i_13_  &  wire6478 ) ;
 assign wire6479 = ( n_n453  &  wire308 ) | ( wire19  &  wire746 ) ;
 assign wire8 = ( i_9_  &  i_10_ ) ;
 assign wire21 = ( i_3_  &  (~ i_4_) ) ;
 assign wire23 = ( (~ i_8_)  &  (~ i_3_) ) ;
 assign wire414 = ( i_9_  &  i_10_ ) | ( i_9_  &  i_8_ ) | ( i_10_  &  (~ i_8_) ) ;
 assign wire648 = ( wire1848 ) | ( wire1849 ) | ( wire33  &  wire649 ) ;
 assign wire1841 = ( wire379  &  wire30 ) | ( wire30  &  wire1844 ) | ( wire30  &  wire1845 ) ;
 assign wire6491 = ( n_n35  &  n_n612 ) | ( wire26  &  wire6488 ) ;
 assign n_n877 = ( wire1841 ) | ( wire6491 ) | ( (~ i_5_)  &  wire648 ) ;
 assign wire1832 = ( wire316  &  wire6494 ) | ( wire6493  &  wire6494 ) ;
 assign wire1833 = ( i_7_  &  wire1838 ) | ( i_7_  &  wire1839 ) ;
 assign wire6495 = ( i_1_  &  wire395 ) | ( i_1_  &  wire34  &  n_n35 ) ;
 assign wire6496 = ( n_n633  &  wire299 ) | ( n_n612  &  wire316 ) ;
 assign n_n876 = ( wire1832 ) | ( wire1833 ) | ( wire6495 ) | ( wire6496 ) ;
 assign wire1823 = ( wire36  &  wire1829 ) | ( i_2_  &  wire36  &  wire653 ) ;
 assign wire1825 = ( i_11_  &  wire384 ) ;
 assign wire6500 = ( n_n36  &  wire385 ) | ( n_n358  &  wire6499 ) ;
 assign wire6501 = ( n_n818  &  (~ wire181) ) | ( i_1_  &  wire304 ) ;
 assign n_n878 = ( wire1823 ) | ( wire1825 ) | ( wire6500 ) | ( wire6501 ) ;
 assign n_n879 = ( wire1814 ) | ( wire6506 ) | ( wire6507 ) ;
 assign n_n881 = ( wire1805 ) | ( wire1806 ) | ( wire1808 ) | ( wire6512 ) ;
 assign wire6520 = ( wire1796 ) | ( wire1797 ) | ( _8232 ) ;
 assign wire18 = ( i_9_  &  i_8_ ) ;
 assign wire55 = ( i_3_ ) | ( i_2_ ) ;
 assign wire126 = ( i_10_  &  (~ i_8_)  &  i_3_ ) ;
 assign wire278 = ( i_10_  &  (~ i_8_) ) ;
 assign wire283 = ( i_9_  &  i_1_ ) ;
 assign wire327 = ( (~ i_6_)  &  i_3_  &  i_2_  &  i_0_ ) ;
 assign wire343 = ( i_9_  &  i_5_  &  i_0_ ) ;
 assign wire348 = ( i_10_  &  (~ i_5_)  &  i_0_ ) ;
 assign wire386 = ( i_9_  &  i_7_  &  i_2_ ) ;
 assign wire284 = ( (~ i_9_)  &  (~ i_13_)  &  (~ i_12_)  &  i_11_ ) ;
 assign wire483 = ( wire1679 ) | ( wire1681 ) | ( n_n748  &  wire484 ) ;
 assign wire6615 = ( wire1673 ) | ( wire1675 ) ;
 assign wire6616 = ( wire1672 ) | ( wire341  &  n_n852  &  wire482 ) ;
 assign n_n1240 = ( wire6615 ) | ( wire6616 ) | ( wire284  &  wire483 ) ;
 assign wire344 = ( (~ i_9_)  &  (~ i_10_) ) ;
 assign wire502 = ( wire1669 ) | ( wire6624 ) | ( (~ i_7_)  &  wire503 ) ;
 assign wire6594 = ( (~ i_13_)  &  (~ i_12_)  &  i_11_ ) ;
 assign wire6627 = ( wire1661 ) | ( wire1663 ) | ( wire501  &  wire6618 ) ;
 assign n_n1241 = ( wire6627 ) | ( wire344  &  wire502  &  wire6594 ) ;
 assign n_n1248 = ( wire1647 ) | ( wire1648 ) | ( n_n638  &  wire454 ) ;
 assign n_n1229 = ( n_n1253 ) | ( wire1564 ) | ( wire6693 ) | ( _8407 ) ;
 assign wire1547 = ( _1113 ) | ( _1114 ) ;
 assign wire6704 = ( n_n1250 ) | ( n_n1256 ) | ( n_n1255 ) | ( wire6667 ) ;
 assign wire1535 = ( _901 ) | ( wire569  &  _8747 ) ;
 assign wire1537 = ( _897 ) | ( i_13_  &  (~ i_12_)  &  wire6714 ) ;
 assign wire6715 = ( wire1534 ) | ( _893 ) | ( _894 ) ;
 assign n_n1236 = ( wire1535 ) | ( wire1537 ) | ( wire6715 ) ;
 assign n_n1261 = ( _1054 ) | ( _8521 ) | ( wire451  &  _8509 ) ;
 assign n_n1231 = ( n_n1258 ) | ( wire1490 ) | ( wire6752 ) | ( wire6759 ) ;
 assign n_n1233 = ( n_n1264 ) | ( n_n1265 ) | ( wire6780 ) | ( _8610 ) ;
 assign wire6791 = ( wire1425 ) | ( wire6730 ) | ( wire6731 ) | ( wire6789 ) ;
 assign wire1375 = ( wire1383  &  wire6831 ) | ( n_n792  &  wire31  &  wire6831 ) ;
 assign wire1376 = ( (~ i_8_)  &  i_11_  &  n_n779  &  n_n849 ) ;
 assign wire6834 = ( wire1377 ) | ( n_n853  &  wire438 ) ;
 assign n_n1121 = ( wire1375 ) | ( wire1376 ) | ( wire6834 ) ;
 assign wire1362 = ( (~ i_13_)  &  (~ i_12_)  &  i_11_  &  wire6835 ) ;
 assign wire1363 = ( (~ i_8_)  &  i_6_  &  n_n716  &  n_n675 ) ;
 assign wire1366 = ( (~ i_6_)  &  wire1372 ) | ( wire6838  &  _9115 ) ;
 assign wire6840 = ( i_6_  &  wire443 ) | ( n_n849  &  wire442 ) ;
 assign n_n1120 = ( wire1362 ) | ( wire1363 ) | ( wire1366 ) | ( wire6840 ) ;
 assign wire1186 = ( (~ i_6_)  &  wire6945 ) | ( wire636  &  _9055 ) ;
 assign wire1195 = ( _684 ) | ( _685 ) ;
 assign wire6941 = ( wire1194 ) | ( wire1196 ) | ( wire313  &  wire9 ) ;
 assign wire6946 = ( i_1_  &  wire340 ) | ( (~ i_13_)  &  i_1_  &  wire632 ) ;
 assign n_n1108 = ( wire1186 ) | ( wire1195 ) | ( wire6941 ) | ( wire6946 ) ;
 assign wire14 = ( (~ i_4_)  &  i_2_ ) ;
 assign wire6956 = ( n_n412  &  wire593 ) | ( wire594  &  wire6952 ) ;
 assign n_n1189 = ( wire6956 ) | ( _536 ) | ( _537 ) ;
 assign wire1096 = ( (~ i_7_)  &  wire6996 ) | ( wire301  &  _9198 ) ;
 assign wire1097 = ( i_7_  &  wire1103 ) | ( n_n672  &  _9200 ) ;
 assign wire6997 = ( wire1094 ) | ( i_7_  &  (~ i_2_)  &  wire628 ) ;
 assign n_n1187 = ( wire1096 ) | ( wire1097 ) | ( wire6997 ) ;
 assign n_n658 = ( i_5_  &  i_6_  &  (~ i_3_) ) ;
 assign n_n741 = ( (~ i_9_)  &  (~ i_10_)  &  (~ i_11_) ) ;
 assign n_n566 = ( (~ i_9_)  &  (~ i_10_)  &  (~ i_12_) ) ;
 assign n_n764 = ( (~ i_9_)  &  i_7_  &  i_8_ ) ;
 assign n_n701 = ( (~ i_10_)  &  (~ i_12_)  &  (~ i_11_) ) ;
 assign wire323 = ( (~ i_5_)  &  (~ i_1_) ) ;
 assign wire325 = ( i_6_  &  (~ i_1_) ) ;
 assign wire326 = ( (~ i_6_)  &  (~ i_1_) ) ;
 assign wire947 = ( wire954  &  wire7085 ) | ( wire7084  &  wire7085 ) ;
 assign wire7088 = ( wire948 ) | ( wire533  &  wire7083 ) ;
 assign n_n970 = ( wire947 ) | ( wire7088 ) | ( _196 ) | ( _197 ) ;
 assign wire937 = ( n_n741  &  wire536  &  _9539 ) ;
 assign wire20 = ( i_5_  &  i_0_ ) ;
 assign wire578 = ( n_n752  &  wire24 ) | ( n_n819  &  wire6848 ) ;
 assign wire925 = ( (~ i_7_)  &  i_5_  &  n_n838  &  wire7094 ) ;
 assign wire7102 = ( wire927 ) | ( wire12  &  n_n670  &  wire579 ) ;
 assign wire881 = ( n_n719  &  n_n837  &  wire7119 ) ;
 assign wire882 = ( (~ i_9_)  &  (~ i_13_)  &  (~ i_12_)  &  wire7121 ) ;
 assign wire884 = ( n_n761  &  wire406 ) | ( n_n761  &  wire887 ) | ( n_n761  &  wire7122 ) ;
 assign n_n984 = ( wire836 ) | ( wire7155 ) | ( _267 ) | ( _268 ) ;
 assign n_n983 = ( wire73 ) | ( wire824 ) | ( wire825 ) | ( wire7161 ) ;
 assign wire7167 = ( wire121 ) | ( wire814 ) | ( wire725  &  wire7164 ) ;
 assign wire7168 = ( wire13  &  wire723 ) | ( wire724  &  wire7163 ) ;
 assign n_n965 = ( n_n991 ) | ( n_n993 ) | ( wire256 ) | ( wire7196 ) ;
 assign wire7232 = ( wire237 ) | ( wire238 ) | ( wire7214 ) | ( wire7231 ) ;
 assign wire40 = ( (~ i_10_)  &  (~ i_13_)  &  n_n838  &  wire7322 ) ;
 assign wire50 = ( n_n687  &  wire57 ) | ( n_n687  &  n_n729  &  wire7325 ) ;
 assign wire52 = ( wire16  &  wire59 ) | ( wire16  &  wire60 ) | ( wire16  &  wire7327 ) ;
 assign wire7329 = ( wire313  &  wire9 ) | ( n_n729  &  wire7324 ) ;
 assign n_n957 = ( wire40 ) | ( wire50 ) | ( wire52 ) | ( wire7329 ) ;
 assign n_n816 = ( (~ i_10_)  &  (~ i_13_)  &  i_11_ ) ;
 assign n_n853 = ( (~ i_13_)  &  i_12_  &  i_11_ ) ;
 assign n_n779 = ( i_4_  &  (~ i_1_)  &  (~ i_2_) ) ;
 assign n_n795 = ( (~ i_9_)  &  (~ i_7_)  &  (~ i_8_) ) ;
 assign wire17 = ( (~ i_13_)  &  i_4_  &  i_12_  &  i_11_ ) ;
 assign wire33 = ( i_1_  &  i_2_ ) ;
 assign wire35 = ( (~ i_5_)  &  i_4_ ) ;
 assign wire37 = ( (~ i_10_)  &  (~ i_13_)  &  i_4_  &  i_12_ ) ;
 assign n_n835 = ( (~ i_1_)  &  (~ i_2_)  &  (~ i_0_) ) ;
 assign wire68 = ( (~ i_10_)  &  (~ i_8_)  &  wire17  &  n_n835 ) ;
 assign wire288 = ( (~ i_8_)  &  (~ i_5_) ) ;
 assign wire313 = ( (~ i_10_)  &  (~ i_13_)  &  i_12_  &  i_11_ ) ;
 assign wire322 = ( (~ i_9_)  &  i_8_  &  i_5_  &  i_6_ ) ;
 assign wire336 = ( (~ i_10_)  &  (~ i_8_)  &  (~ i_6_)  &  (~ i_2_) ) ;
 assign wire420 = ( (~ i_6_)  &  (~ i_2_)  &  i_0_ ) | ( (~ i_1_)  &  (~ i_2_)  &  i_0_ ) ;
 assign n_n833 = ( i_1_  &  (~ i_2_)  &  i_0_ ) ;
 assign n_n538 = ( i_5_  &  i_3_  &  (~ i_4_) ) ;
 assign n_n850 = ( (~ i_7_)  &  (~ i_8_)  &  i_6_ ) ;
 assign n_n498 = ( i_10_  &  (~ i_13_)  &  i_12_  &  (~ i_11_) ) ;
 assign n_n838 = ( (~ i_1_)  &  (~ i_2_)  &  i_0_ ) ;
 assign n_n748 = ( (~ i_7_)  &  i_8_  &  i_6_ ) ;
 assign n_n725 = ( (~ i_10_)  &  (~ i_13_)  &  i_12_  &  (~ i_11_) ) ;
 assign wire341 = ( i_9_  &  (~ i_5_)  &  i_3_  &  (~ i_4_) ) ;
 assign n_n665 = ( i_13_  &  (~ i_12_) ) ;
 assign wire427 = ( n_n623  &  wire429 ) | ( n_n619  &  wire428 ) ;
 assign wire1756 = ( i_9_  &  i_10_  &  i_8_  &  wire426 ) ;
 assign wire6555 = ( wire12  &  n_n638 ) | ( n_n623  &  wire6554 ) ;
 assign wire425 = ( wire1756 ) | ( wire6555 ) | ( i_7_  &  wire427 ) ;
 assign wire6557 = ( (~ i_8_)  &  i_13_  &  (~ i_11_) ) ;
 assign n_n609 = ( i_10_  &  (~ i_8_)  &  (~ i_11_) ) ;
 assign wire1746 = ( i_5_  &  i_6_  &  wire6559 ) | ( i_6_  &  i_0_  &  wire6559 ) ;
 assign wire1744 = ( i_9_  &  i_10_  &  wire6557  &  wire6558 ) ;
 assign n_n623 = ( i_9_  &  i_8_  &  (~ i_11_) ) ;
 assign n_n619 = ( i_9_  &  i_10_  &  i_8_ ) ;
 assign wire376 = ( i_7_  &  i_5_  &  i_1_ ) ;
 assign wire436 = ( n_n835 ) | ( n_n624 ) | ( wire1740 ) | ( wire1741 ) ;
 assign wire435 = ( n_n619  &  wire376 ) | ( n_n623  &  wire436 ) ;
 assign n_n830 = ( i_1_  &  (~ i_2_)  &  (~ i_0_) ) ;
 assign n_n633 = ( i_5_  &  i_6_  &  i_3_ ) ;
 assign n_n631 = ( (~ i_5_)  &  i_6_  &  i_3_ ) ;
 assign wire434 = ( n_n833  &  n_n633 ) | ( n_n830  &  n_n631 ) ;
 assign n_n716 = ( (~ i_13_)  &  i_12_  &  (~ i_11_) ) ;
 assign n_n849 = ( (~ i_10_)  &  (~ i_13_)  &  i_12_ ) ;
 assign n_n36 = ( (~ i_8_)  &  i_11_ ) ;
 assign n_n685 = ( (~ i_3_)  &  i_4_  &  (~ i_1_) ) ;
 assign wire309 = ( (~ i_9_)  &  i_8_ ) ;
 assign wire439 = ( (~ i_9_)  &  i_7_ ) | ( (~ i_10_)  &  (~ i_7_) ) ;
 assign wire438 = ( n_n779  &  wire309 ) | ( n_n685  &  wire439 ) ;
 assign n_n545 = ( (~ i_13_)  &  (~ i_12_)  &  i_11_ ) ;
 assign n_n675 = ( (~ i_3_)  &  (~ i_1_)  &  (~ i_2_) ) ;
 assign wire29 = ( i_7_  &  (~ i_2_) ) ;
 assign wire289 = ( (~ i_8_)  &  i_6_ ) ;
 assign n_n792 = ( (~ i_10_)  &  (~ i_7_)  &  (~ i_8_) ) ;
 assign wire295 = ( (~ i_13_)  &  i_4_  &  i_12_ ) ;
 assign wire6837 = ( (~ i_13_)  &  i_4_  &  i_12_  &  (~ i_1_) ) ;
 assign wire443 = ( n_n675  &  wire295 ) | ( n_n792  &  wire6837 ) ;
 assign wire269 = ( (~ i_7_)  &  i_6_ ) ;
 assign wire442 = ( n_n779  &  wire289 ) | ( n_n685  &  wire269 ) ;
 assign n_n570 = ( (~ i_13_)  &  (~ i_12_) ) ;
 assign n_n787 = ( (~ i_13_)  &  i_11_ ) ;
 assign n_n769 = ( (~ i_9_)  &  i_8_  &  i_6_ ) ;
 assign n_n819 = ( (~ i_9_)  &  i_7_  &  i_6_ ) ;
 assign n_n273 = ( (~ i_3_)  &  i_1_  &  (~ i_2_) ) ;
 assign wire381 = ( (~ i_13_)  &  (~ i_12_)  &  (~ i_11_) ) ;
 assign wire12 = ( i_5_  &  i_6_ ) ;
 assign wire377 = ( (~ i_1_)  &  (~ i_0_) ) ;
 assign n_n847 = ( (~ i_1_)  &  i_2_  &  (~ i_0_) ) ;
 assign wire27 = ( (~ i_7_)  &  (~ i_8_) ) ;
 assign n_n581 = ( i_9_  &  (~ i_7_)  &  (~ i_8_) ) ;
 assign wire264 = ( i_1_  &  i_0_ ) ;
 assign n_n638 = ( i_9_  &  i_7_  &  i_8_ ) ;
 assign wire15 = ( i_3_  &  i_1_ ) ;
 assign n_n814 = ( i_3_  &  i_1_  &  i_2_ ) ;
 assign n_n541 = ( (~ i_5_)  &  i_3_  &  (~ i_4_) ) ;
 assign wire28 = ( (~ i_7_)  &  (~ i_6_) ) ;
 assign n_n746 = ( (~ i_7_)  &  i_8_  &  (~ i_6_) ) ;
 assign wire333 = ( i_1_  &  (~ i_0_) ) ;
 assign n_n453 = ( i_10_  &  (~ i_11_) ) ;
 assign n_n761 = ( (~ i_13_)  &  i_12_ ) ;
 assign n_n421 = ( i_9_  &  i_10_  &  i_11_ ) ;
 assign n_n415 = ( i_10_  &  i_12_  &  i_11_ ) ;
 assign n_n369 = ( i_3_  &  (~ i_4_)  &  i_1_ ) ;
 assign wire25 = ( i_9_  &  i_7_ ) ;
 assign n_n358 = ( i_9_  &  i_7_  &  i_6_ ) ;
 assign n_n412 = ( i_3_  &  (~ i_4_)  &  i_2_ ) ;
 assign wire279 = ( (~ i_10_)  &  (~ i_6_) ) ;
 assign n_n773 = ( (~ i_10_)  &  (~ i_8_)  &  (~ i_6_) ) ;
 assign n_n844 = ( i_1_  &  i_2_  &  i_0_ ) ;
 assign wire13 = ( i_5_  &  (~ i_6_) ) ;
 assign n_n639 = ( i_5_  &  (~ i_6_)  &  i_3_ ) ;
 assign wire286 = ( i_7_  &  i_8_ ) ;
 assign n_n185 = ( i_7_  &  i_8_  &  (~ i_5_) ) ;
 assign n_n432 = ( i_9_  &  i_10_  &  i_12_ ) ;
 assign n_n826 = ( i_3_  &  i_1_  &  i_0_ ) ;
 assign n_n183 = ( i_9_  &  i_12_ ) ;
 assign wire96 = ( (~ i_3_) ) | ( (~ i_2_) ) ;
 assign n_n818 = ( i_3_  &  i_2_  &  i_0_ ) ;
 assign n_n153 = ( i_3_  &  (~ i_4_)  &  i_0_ ) ;
 assign n_n316 = ( i_12_  &  (~ i_11_) ) ;
 assign n_n197 = ( i_9_  &  i_11_ ) ;
 assign n_n843 = ( (~ i_7_)  &  (~ i_8_)  &  (~ i_6_) ) ;
 assign n_n699 = ( (~ i_10_)  &  (~ i_7_)  &  (~ i_6_) ) ;
 assign wire293 = ( (~ i_3_)  &  i_4_ ) ;
 assign n_n678 = ( (~ i_3_)  &  i_4_  &  (~ i_0_) ) ;
 assign n_n671 = ( (~ i_3_)  &  (~ i_2_)  &  (~ i_0_) ) ;
 assign wire26 = ( (~ i_5_)  &  i_6_ ) ;
 assign n_n176 = ( i_8_  &  (~ i_5_)  &  i_6_ ) ;
 assign n_n712 = ( i_5_  &  (~ i_3_)  &  i_4_ ) ;
 assign n_n751 = ( (~ i_9_)  &  (~ i_13_) ) ;
 assign wire265 = ( (~ i_1_)  &  (~ i_2_) ) ;
 assign n_n719 = ( (~ i_9_)  &  (~ i_13_)  &  (~ i_11_) ) ;
 assign wire31 = ( (~ i_3_)  &  (~ i_1_) ) ;
 assign n_n687 = ( (~ i_3_)  &  (~ i_1_)  &  i_0_ ) ;
 assign wire34 = ( i_7_  &  i_5_ ) ;
 assign n_n827 = ( (~ i_9_)  &  i_7_  &  i_5_ ) ;
 assign wire267 = ( (~ i_9_)  &  i_7_ ) ;
 assign n_n683 = ( (~ i_3_)  &  (~ i_1_)  &  (~ i_0_) ) ;
 assign n_n275 = ( (~ i_9_)  &  i_7_  &  (~ i_8_) ) ;
 assign n_n35 = ( i_8_  &  i_12_ ) ;
 assign wire69 = ( (~ i_6_)  &  (~ i_0_)  &  wire17  &  n_n792 ) ;
 assign wire370 = ( (~ i_13_)  &  i_4_  &  i_11_ ) ;
 assign wire70 = ( (~ i_5_)  &  (~ i_6_)  &  n_n792  &  wire370 ) ;
 assign n_n791 = ( i_4_  &  (~ i_1_)  &  (~ i_0_) ) ;
 assign wire106 = ( n_n853  &  n_n792  &  n_n791 ) ;
 assign wire6735 = ( (~ i_9_)  &  i_4_  &  i_1_ ) ;
 assign wire1652 = ( i_5_  &  i_6_  &  i_3_  &  wire6632 ) ;
 assign wire1656 = ( (~ i_5_)  &  (~ i_6_)  &  i_3_  &  _8334 ) ;
 assign wire6633 = ( n_n639  &  n_n852 ) | ( n_n631  &  n_n840 ) ;
 assign wire454 = ( wire1652 ) | ( n_n637  &  wire1656 ) | ( n_n637  &  wire6633 ) ;
 assign n_n635 = ( (~ i_5_)  &  (~ i_6_)  &  i_3_ ) ;
 assign wire453 = ( i_0_  &  n_n639  &  wire265 ) | ( (~ i_0_)  &  wire265  &  n_n635 ) ;
 assign wire1647 = ( wire6630  &  wire6631 ) | ( n_n844  &  wire317  &  wire6631 ) ;
 assign wire1648 = ( i_9_  &  i_8_  &  wire453  &  wire6563 ) ;
 assign n_n752 = ( i_7_  &  i_8_  &  i_6_ ) ;
 assign wire307 = ( i_9_  &  i_5_  &  i_3_  &  (~ i_4_) ) ;
 assign n_n592 = ( i_10_  &  (~ i_7_)  &  (~ i_8_) ) ;
 assign n_n832 = ( i_7_  &  (~ i_8_)  &  (~ i_6_) ) ;
 assign n_n852 = ( (~ i_1_)  &  i_2_  &  i_0_ ) ;
 assign wire6587 = ( wire1708 ) | ( wire1709 ) | ( n_n453  &  wire308 ) ;
 assign n_n1243 = ( wire6587 ) | ( _951 ) | ( _952 ) ;
 assign wire388 = ( (~ i_7_)  &  (~ i_6_)  &  i_0_ ) ;
 assign wire42 = ( (~ i_5_)  &  i_1_  &  i_2_ ) | ( i_1_  &  i_2_  &  i_0_ ) ;
 assign wire6591 = ( (~ i_5_)  &  (~ i_6_)  &  i_2_ ) | ( (~ i_6_)  &  i_2_  &  i_0_ ) ;
 assign wire465 = ( wire388 ) | ( wire42 ) | ( wire6591 ) ;
 assign n_n598 = ( (~ i_6_)  &  i_2_  &  i_0_ ) ;
 assign n_n575 = ( (~ i_10_)  &  (~ i_13_)  &  (~ i_12_) ) ;
 assign wire19 = ( i_8_  &  (~ i_3_) ) ;
 assign wire9 = ( (~ i_9_)  &  i_4_ ) ;
 assign n_n672 = ( (~ i_3_)  &  i_4_  &  (~ i_2_) ) ;
 assign n_n810 = ( (~ i_9_)  &  i_6_  &  i_4_ ) ;
 assign wire371 = ( (~ i_13_)  &  i_4_  &  i_1_ ) ;
 assign wire301 = ( (~ i_13_)  &  (~ i_12_)  &  i_11_  &  (~ i_2_) ) ;
 assign wire346 = ( (~ i_9_)  &  (~ i_3_)  &  i_4_  &  (~ i_2_) ) ;
 assign wire11 = ( (~ i_5_)  &  (~ i_6_) ) ;
 assign n_n653 = ( (~ i_5_)  &  (~ i_6_)  &  (~ i_3_) ) ;
 assign n_n526 = ( (~ i_12_)  &  (~ i_11_) ) ;
 assign n_n534 = ( i_3_  &  (~ i_1_)  &  i_2_ ) ;
 assign n_n242 = ( (~ i_10_)  &  (~ i_7_)  &  (~ i_11_) ) ;
 assign n_n656 = ( i_10_  &  (~ i_7_)  &  (~ i_11_) ) ;
 assign n_n194 = ( i_9_  &  i_7_  &  i_11_ ) ;
 assign n_n346 = ( (~ i_4_)  &  i_1_  &  i_2_ ) ;
 assign n_n842 = ( (~ i_10_)  &  (~ i_13_) ) ;
 assign wire281 = ( i_4_  &  (~ i_1_) ) ;
 assign n_n755 = ( (~ i_9_)  &  (~ i_13_)  &  i_11_ ) ;
 assign n_n846 = ( i_5_  &  i_3_  &  i_4_ ) ;
 assign wire1503 = ( _1047 ) | ( n_n755  &  n_n756  &  wire479 ) ;
 assign wire1504 = ( n_n853  &  wire51 ) | ( n_n853  &  n_n779  &  n_n768 ) ;
 assign wire6745 = ( wire1500 ) | ( wire1501 ) | ( wire1502 ) ;
 assign n_n1258 = ( wire1503 ) | ( wire1504 ) | ( wire6745 ) ;
 assign n_n670 = ( (~ i_3_)  &  (~ i_2_)  &  i_0_ ) ;
 assign wire6669 = ( (~ i_3_)  &  (~ i_1_)  &  (~ i_2_)  &  (~ i_0_) ) ;
 assign wire113 = ( wire17  &  wire6669 ) ;
 assign n_n756 = ( i_7_  &  i_8_  &  (~ i_6_) ) ;
 assign n_n550 = ( (~ i_9_)  &  (~ i_13_)  &  (~ i_12_) ) ;
 assign n_n732 = ( i_5_  &  (~ i_3_)  &  (~ i_4_) ) ;
 assign wire484 = ( i_5_  &  n_n833  &  wire277 ) | ( (~ i_5_)  &  n_n830  &  wire277 ) ;
 assign wire1679 = ( n_n838  &  n_n746  &  n_n732 ) ;
 assign wire1681 = ( n_n752  &  n_n840  &  n_n735 ) ;
 assign n_n729 = ( (~ i_10_)  &  (~ i_13_)  &  (~ i_11_) ) ;
 assign wire482 = ( n_n752  &  n_n575 ) | ( n_n756  &  n_n729 ) ;
 assign wire487 = ( i_9_  &  i_13_  &  (~ i_12_) ) | ( i_9_  &  i_13_  &  i_1_ ) ;
 assign wire486 = ( i_9_  &  i_10_  &  i_13_ ) | ( i_10_  &  (~ i_6_)  &  i_13_ ) ;
 assign wire485 = ( i_10_  &  (~ i_6_) ) | ( (~ i_6_)  &  (~ i_1_) ) ;
 assign wire6871 = ( wire1307 ) | ( i_10_  &  (~ i_11_)  &  wire308 ) ;
 assign wire6872 = ( wire1308 ) | ( i_13_  &  (~ i_11_)  &  wire485 ) ;
 assign wire6873 = ( i_6_  &  wire487 ) | ( i_1_  &  wire486 ) ;
 assign n_n1126 = ( wire6871 ) | ( wire6872 ) | ( wire6873 ) ;
 assign wire22 = ( (~ i_4_)  &  i_1_ ) ;
 assign wire38 = ( i_9_ ) | ( (~ i_1_) ) ;
 assign wire297 = ( (~ i_4_)  &  (~ i_12_)  &  i_11_ ) ;
 assign wire1293 = ( wire6875  &  wire6876 ) ;
 assign wire1294 = ( wire364  &  wire6879 ) | ( wire1301  &  wire6879 ) | ( wire1302  &  wire6879 ) ;
 assign wire1295 = ( wire297  &  wire1297 ) | ( wire297  &  wire1298 ) ;
 assign wire1296 = ( n_n346  &  wire1299 ) | ( n_n346  &  wire1300 ) ;
 assign n_n1127 = ( wire1293 ) | ( wire1294 ) | ( wire1295 ) | ( wire1296 ) ;
 assign wire493 = ( i_10_  &  (~ i_7_)  &  i_6_ ) | ( i_10_  &  (~ i_7_)  &  (~ i_11_) ) ;
 assign wire342 = ( i_9_  &  (~ i_12_)  &  i_11_ ) ;
 assign wire393 = ( i_10_  &  i_7_  &  (~ i_6_)  &  (~ i_11_) ) ;
 assign wire491 = ( n_n748  &  wire342 ) | ( n_n183  &  wire393 ) ;
 assign wire1283 = ( i_3_  &  i_1_  &  wire1290 ) | ( i_3_  &  i_1_  &  wire6887 ) ;
 assign wire6890 = ( wire1279 ) | ( wire6888 ) | ( i_3_  &  wire491 ) ;
 assign n_n1112 = ( n_n1126 ) | ( n_n1127 ) | ( wire1283 ) | ( wire6890 ) ;
 assign wire268 = ( i_7_  &  (~ i_6_) ) ;
 assign n_n274 = ( (~ i_13_)  &  (~ i_11_) ) ;
 assign n_n837 = ( i_7_  &  (~ i_8_)  &  i_6_ ) ;
 assign n_n240 = ( (~ i_10_)  &  (~ i_7_)  &  i_8_ ) ;
 assign wire330 = ( i_4_  &  (~ i_2_) ) ;
 assign n_n771 = ( i_4_  &  (~ i_2_)  &  (~ i_0_) ) ;
 assign n_n606 = ( (~ i_5_)  &  (~ i_6_)  &  (~ i_2_) ) ;
 assign n_n813 = ( (~ i_9_)  &  i_5_  &  i_4_ ) ;
 assign wire290 = ( (~ i_6_)  &  i_0_ ) ;
 assign wire308 = ( i_9_  &  i_13_  &  (~ i_12_) ) ;
 assign wire318 = ( (~ i_9_)  &  i_8_  &  i_4_ ) ;
 assign n_n768 = ( (~ i_9_)  &  i_8_  &  i_5_ ) ;
 assign wire6748 = ( i_2_  &  i_0_ ) ;
 assign wire494 = ( wire33  &  n_n768 ) | ( n_n769  &  wire6748 ) ;
 assign wire360 = ( i_10_  &  (~ i_5_)  &  (~ i_11_) ) ;
 assign wire1637 = ( wire308  &  wire1639 ) | ( wire308  &  wire1640 ) ;
 assign wire1643 = ( n_n658  &  wire25 ) | ( wire25  &  n_n683 ) | ( wire25  &  wire1644 ) ;
 assign wire6640 = ( n_n675  &  wire6637 ) | ( n_n358  &  wire6638 ) ;
 assign wire497 = ( wire1637 ) | ( n_n665  &  wire1643 ) | ( n_n665  &  wire6640 ) ;
 assign wire1634 = ( i_13_  &  (~ i_12_)  &  n_n675  &  wire360 ) ;
 assign wire1635 = ( i_13_  &  (~ i_12_)  &  (~ i_11_)  &  wire6636 ) ;
 assign n_n1250 = ( wire1634 ) | ( wire1635 ) | ( (~ i_11_)  &  wire497 ) ;
 assign wire294 = ( (~ i_10_)  &  (~ i_13_)  &  (~ i_12_)  &  i_11_ ) ;
 assign wire296 = ( (~ i_4_)  &  i_1_  &  i_2_  &  i_0_ ) ;
 assign wire503 = ( wire22  &  wire6622 ) | ( n_n735  &  wire6623 ) ;
 assign wire1669 = ( (~ i_4_)  &  i_2_  &  wire317 ) ;
 assign wire6624 = ( n_n746  &  wire6620 ) | ( n_n346  &  wire6621 ) ;
 assign wire277 = ( (~ i_3_)  &  (~ i_4_) ) ;
 assign wire501 = ( (~ i_5_)  &  n_n847  &  wire277 ) | ( i_5_  &  n_n852  &  wire277 ) ;
 assign wire272 = ( i_3_  &  (~ i_4_)  &  i_1_  &  i_2_ ) ;
 assign wire298 = ( i_3_  &  (~ i_4_)  &  (~ i_1_)  &  i_2_ ) ;
 assign wire311 = ( i_10_  &  (~ i_6_) ) ;
 assign wire363 = ( i_10_  &  (~ i_6_)  &  (~ i_11_) ) ;
 assign wire1274 = ( i_9_  &  wire272 ) | ( i_9_  &  wire1277 ) ;
 assign wire6893 = ( (~ i_12_)  &  wire298 ) | ( wire22  &  wire334 ) ;
 assign wire6896 = ( wire1267 ) | ( wire6894 ) | ( n_n526  &  wire298 ) ;
 assign wire104 = ( i_9_  &  i_10_  &  i_12_  &  i_11_ ) ;
 assign wire270 = ( i_9_  &  i_8_  &  i_12_ ) ;
 assign wire379 = ( i_3_  &  i_1_  &  i_11_ ) ;
 assign wire507 = ( i_10_  &  (~ i_8_)  &  i_6_ ) | ( i_10_  &  (~ i_8_)  &  (~ i_11_) ) ;
 assign wire1263 = ( (~ i_8_)  &  wire1266 ) | ( (~ i_8_)  &  wire15  &  n_n415 ) ;
 assign wire6902 = ( n_n609  &  (~ wire96) ) | ( n_n597  &  wire6901 ) ;
 assign wire6905 = ( wire1255 ) | ( wire6904 ) | ( wire507  &  wire6899 ) ;
 assign wire181 = ( (~ i_6_) ) | ( (~ i_12_) ) ;
 assign wire364 = ( i_10_  &  (~ i_7_)  &  (~ i_8_)  &  (~ i_6_) ) ;
 assign wire512 = ( i_3_  &  (~ i_12_)  &  i_2_ ) | ( i_3_  &  i_1_  &  i_2_ ) ;
 assign wire516 = ( (~ i_6_)  &  (~ i_11_) ) | ( (~ i_12_)  &  (~ i_11_) ) ;
 assign wire513 = ( (~ i_12_)  &  i_2_ ) | ( i_1_  &  i_2_ ) ;
 assign n_n822 = ( (~ i_10_)  &  i_12_  &  i_11_ ) ;
 assign n_n840 = ( i_1_  &  i_2_  &  (~ i_0_) ) ;
 assign n_n710 = ( (~ i_5_)  &  (~ i_3_)  &  i_4_ ) ;
 assign wire520 = ( i_6_  &  n_n847  &  wire27 ) | ( (~ i_6_)  &  wire27  &  n_n840 ) ;
 assign wire1629 = ( (~ i_13_)  &  i_12_  &  n_n741  &  wire6647 ) ;
 assign wire1630 = ( n_n844  &  n_n719  &  n_n837 ) ;
 assign wire519 = ( wire1629 ) | ( wire1630 ) | ( n_n725  &  wire520 ) ;
 assign wire6644 = ( i_7_  &  (~ i_8_)  &  (~ i_3_) ) ;
 assign wire518 = ( n_n837  &  wire277 ) | ( wire22  &  wire6644 ) ;
 assign n_n735 = ( (~ i_5_)  &  (~ i_3_)  &  (~ i_4_) ) ;
 assign wire6642 = ( (~ i_6_)  &  (~ i_3_)  &  (~ i_4_) ) ;
 assign wire517 = ( n_n843  &  n_n735 ) | ( n_n795  &  wire6642 ) ;
 assign wire1624 = ( n_n732  &  n_n837  &  _8446 ) ;
 assign wire6651 = ( wire517  &  wire6643 ) | ( wire518  &  wire6645 ) ;
 assign n_n1256 = ( wire1624 ) | ( wire6651 ) | ( n_n732  &  wire519 ) ;
 assign wire525 = ( i_0_  &  wire265  &  n_n846 ) | ( (~ i_0_)  &  wire265  &  n_n851 ) ;
 assign wire524 = ( n_n833  &  n_n846 ) | ( n_n830  &  n_n851 ) ;
 assign wire523 = ( n_n746  &  wire525 ) | ( n_n748  &  wire524 ) ;
 assign wire6756 = ( i_5_  &  (~ i_13_)  &  i_12_ ) ;
 assign wire521 = ( (~ i_13_)  &  wire296 ) | ( n_n346  &  wire6756 ) ;
 assign wire1490 = ( n_n764  &  wire1493 ) | ( n_n764  &  wire6749 ) | ( n_n764  &  wire6750 ) ;
 assign wire6752 = ( wire1488 ) | ( wire37  &  wire494 ) ;
 assign wire6759 = ( wire1474 ) | ( wire6757 ) | ( n_n755  &  wire523 ) ;
 assign wire350 = ( i_7_  &  (~ i_5_)  &  (~ i_6_)  &  (~ i_2_) ) ;
 assign wire529 = ( (~ i_6_)  &  i_0_  &  n_n741 ) | ( i_6_  &  i_0_  &  n_n566 ) ;
 assign wire16 = ( (~ i_5_)  &  i_0_ ) ;
 assign wire533 = ( n_n746  &  n_n575 ) | ( n_n843  &  n_n729 ) ;
 assign wire536 = ( (~ i_8_)  &  (~ i_3_) ) | ( (~ i_7_)  &  (~ i_2_) ) ;
 assign n_n597 = ( i_10_  &  i_7_  &  (~ i_8_) ) ;
 assign n_n651 = ( i_10_  &  i_7_  &  i_8_ ) ;
 assign wire1610 = ( _1081 ) | ( n_n725  &  n_n832  &  wire541 ) ;
 assign wire6658 = ( wire1611 ) | ( wire1620  &  wire6654 ) | ( wire6653  &  wire6654 ) ;
 assign n_n1255 = ( wire1610 ) | ( wire6658 ) | ( _1084 ) | ( _1085 ) ;
 assign wire405 = ( (~ i_13_)  &  i_11_  &  n_n835  &  n_n710 ) ;
 assign wire546 = ( i_5_  &  n_n819  &  wire277 ) | ( (~ i_5_)  &  n_n699  &  wire277 ) ;
 assign wire1603 = ( n_n849  &  n_n746  &  n_n710 ) ;
 assign wire1605 = ( (~ i_10_)  &  (~ i_12_)  &  (~ i_11_)  &  _8496 ) ;
 assign wire545 = ( wire1603 ) | ( wire1605 ) | ( wire381  &  wire546 ) ;
 assign wire544 = ( n_n833  &  n_n712 ) | ( n_n830  &  n_n710 ) ;
 assign wire543 = ( n_n847  &  n_n712 ) | ( n_n852  &  n_n710 ) ;
 assign wire571 = ( n_n712  &  wire573 ) | ( n_n710  &  wire572 ) ;
 assign wire6683 = ( wire73 ) | ( wire1569 ) | ( wire1571 ) | ( wire1572 ) ;
 assign n_n1253 = ( wire6683 ) | ( n_n849  &  wire571 ) ;
 assign wire120 = ( n_n853  &  n_n699  &  n_n678 ) ;
 assign wire6678 = ( wire113 ) | ( wire1582 ) | ( wire1583 ) | ( wire1585 ) ;
 assign wire6922 = ( i_12_  &  (~ i_1_)  &  (~ i_11_) ) ;
 assign wire553 = ( n_n35  &  wire393 ) | ( n_n756  &  wire6922 ) ;
 assign wire6921 = ( i_7_  &  i_12_ ) ;
 assign wire552 = ( n_n638  &  (~ wire181) ) | ( n_n619  &  wire6921 ) ;
 assign wire1221 = ( (~ i_6_)  &  wire1228 ) | ( (~ i_6_)  &  wire6925 ) ;
 assign wire6926 = ( wire1218 ) | ( (~ i_4_)  &  i_1_  &  wire552 ) ;
 assign n_n1128 = ( wire1221 ) | ( wire6926 ) | ( (~ i_4_)  &  wire553 ) ;
 assign wire30 = ( (~ i_7_)  &  (~ i_5_) ) ;
 assign wire352 = ( (~ i_7_)  &  i_2_ ) ;
 assign wire7249 = ( (~ i_12_)  &  i_11_  &  (~ i_0_) ) ;
 assign wire7250 = ( (~ i_7_)  &  i_5_  &  (~ i_6_)  &  i_2_ ) ;
 assign wire557 = ( n_n844  &  wire30 ) | ( wire7249  &  wire7250 ) ;
 assign wire338 = ( i_10_  &  (~ i_5_)  &  i_12_  &  i_0_ ) ;
 assign wire562 = ( i_10_  &  (~ i_7_)  &  i_5_ ) | ( i_10_  &  (~ i_7_)  &  (~ i_11_) ) ;
 assign wire561 = ( i_10_  &  i_5_  &  (~ i_6_) ) | ( i_10_  &  (~ i_6_)  &  (~ i_11_) ) ;
 assign wire560 = ( n_n840  &  wire562 ) | ( wire333  &  wire561 ) ;
 assign wire558 = ( i_10_  &  i_1_  &  (~ i_11_) ) | ( i_10_  &  i_1_  &  i_0_ ) ;
 assign wire176 = ( n_n656  &  wire180 ) | ( n_n656  &  wire182 ) ;
 assign wire7255 = ( wire11  &  wire558 ) | ( wire338  &  wire7254 ) ;
 assign n_n1000 = ( wire176 ) | ( wire7255 ) | ( (~ i_12_)  &  wire560 ) ;
 assign wire375 = ( i_5_  &  i_6_  &  (~ i_12_) ) ;
 assign wire170 = ( (~ i_5_)  &  i_6_  &  (~ i_11_)  &  (~ i_0_) ) ;
 assign wire171 = ( i_6_  &  (~ i_12_)  &  (~ i_11_)  &  (~ i_0_) ) ;
 assign wire172 = ( i_5_  &  i_6_  &  i_0_ ) ;
 assign wire565 = ( wire375 ) | ( wire170 ) | ( wire171 ) | ( wire172 ) ;
 assign wire36 = ( i_6_  &  i_0_ ) ;
 assign wire7257 = ( i_9_  &  i_10_  &  i_12_  &  (~ i_11_) ) ;
 assign wire564 = ( n_n432  &  wire36 ) | ( wire26  &  wire7257 ) ;
 assign n_n503 = ( (~ i_9_)  &  (~ i_8_)  &  i_6_ ) ;
 assign wire73 = ( (~ i_10_)  &  (~ i_7_)  &  wire17  &  n_n683 ) ;
 assign wire121 = ( (~ i_13_)  &  i_12_  &  n_n835  &  n_n712 ) ;
 assign wire573 = ( n_n830  &  n_n756 ) | ( n_n746  &  n_n840 ) ;
 assign wire572 = ( n_n838  &  n_n752 ) | ( n_n833  &  n_n756 ) ;
 assign n_n1264 = ( wire1462 ) | ( wire1463 ) | ( wire1466 ) | ( wire6766 ) ;
 assign n_n1265 = ( wire1450 ) | ( _990 ) | ( _991 ) | ( _993 ) ;
 assign n_n851 = ( (~ i_5_)  &  i_3_  &  i_4_ ) ;
 assign wire574 = ( n_n826  &  wire9 ) | ( (~ wire38)  &  n_n851 ) ;
 assign n_n624 = ( i_5_  &  i_6_  &  (~ i_2_) ) ;
 assign wire24 = ( (~ i_9_)  &  (~ i_13_)  &  i_4_ ) ;
 assign wire931 = ( (~ i_9_)  &  i_8_  &  (~ i_13_)  &  (~ i_12_) ) ;
 assign wire932 = ( (~ i_9_)  &  (~ i_8_)  &  (~ i_13_)  &  (~ i_11_) ) ;
 assign wire579 = ( wire24 ) | ( wire931 ) | ( wire932 ) ;
 assign wire6848 = ( (~ i_13_)  &  (~ i_12_)  &  (~ i_2_) ) ;
 assign wire584 = ( i_0_  &  wire33  &  n_n541 ) | ( (~ i_0_)  &  wire33  &  wire6803 ) ;
 assign wire1418 = ( n_n538  &  n_n850  &  n_n716  &  wire6799 ) ;
 assign wire1419 = ( n_n833  &  n_n538  &  n_n550  &  n_n837 ) ;
 assign wire583 = ( wire1418 ) | ( wire1419 ) | ( n_n843  &  wire584 ) ;
 assign wire410 = ( (~ i_13_)  &  (~ i_12_)  &  n_n835  &  n_n541 ) ;
 assign wire1414 = ( n_n830  &  n_n541  &  n_n550  &  n_n837 ) ;
 assign wire115 = ( i_1_  &  i_2_  &  i_0_  &  wire6807 ) ;
 assign wire1400 = ( n_n835  &  n_n498  &  wire269  &  wire307 ) ;
 assign wire1402 = ( i_9_  &  i_10_  &  wire1406 ) | ( i_9_  &  i_10_  &  wire6812 ) ;
 assign wire6814 = ( wire1403 ) | ( n_n421  &  wire268  &  wire410 ) ;
 assign n_n1234 = ( wire115 ) | ( wire1400 ) | ( wire1402 ) | ( wire6814 ) ;
 assign wire591 = ( i_9_  &  i_7_  &  i_6_ ) | ( i_7_  &  (~ i_5_)  &  i_6_ ) ;
 assign wire594 = ( i_9_  &  i_7_ ) | ( i_7_  &  (~ i_2_) ) ;
 assign wire593 = ( i_9_  &  i_10_ ) | ( i_10_  &  (~ i_7_) ) ;
 assign wire123 = ( (~ i_7_)  &  (~ i_6_)  &  i_3_  &  i_0_ ) ;
 assign wire276 = ( i_5_  &  (~ i_12_) ) ;
 assign wire291 = ( i_3_  &  i_0_ ) ;
 assign wire354 = ( (~ i_7_)  &  (~ i_12_)  &  i_11_ ) ;
 assign wire7287 = ( i_10_  &  (~ i_5_)  &  i_6_  &  i_12_ ) ;
 assign wire7288 = ( (~ i_5_)  &  i_3_  &  i_0_ ) ;
 assign wire596 = ( n_n818  &  wire7287 ) | ( n_n415  &  wire7288 ) ;
 assign n_n277 = ( (~ i_9_)  &  (~ i_7_)  &  (~ i_11_) ) ;
 assign wire6807 = ( i_9_  &  i_10_  &  i_3_  &  (~ i_4_) ) ;
 assign wire1214 = ( i_9_  &  (~ i_7_)  &  i_6_  &  i_11_ ) ;
 assign wire1215 = ( i_10_  &  i_7_  &  (~ i_6_)  &  i_12_ ) ;
 assign wire1216 = ( i_10_  &  (~ i_7_)  &  (~ i_6_)  &  i_11_ ) ;
 assign wire1217 = ( i_9_  &  i_7_  &  i_6_  &  i_12_ ) ;
 assign wire604 = ( wire1214 ) | ( wire1215 ) | ( wire1216 ) | ( wire1217 ) ;
 assign wire606 = ( wire15  &  n_n827 ) | ( n_n819  &  wire291 ) ;
 assign wire1462 = ( (~ i_9_)  &  i_4_  &  wire313  &  wire6762 ) ;
 assign wire1463 = ( n_n822  &  wire24  &  wire6763 ) ;
 assign wire1466 = ( n_n849  &  wire6764 ) | ( n_n849  &  wire9  &  wire287 ) ;
 assign wire6766 = ( wire1464 ) | ( wire37  &  wire606 ) ;
 assign wire292 = ( i_3_  &  i_1_  &  i_2_  &  i_0_ ) ;
 assign wire340 = ( (~ i_9_)  &  (~ i_10_)  &  (~ i_13_)  &  i_4_ ) ;
 assign wire359 = ( (~ i_5_)  &  i_3_  &  i_1_  &  i_2_ ) ;
 assign wire6777 = ( (~ i_9_)  &  i_4_  &  i_2_ ) ;
 assign wire612 = ( n_n818  &  n_n810 ) | ( n_n633  &  wire6777 ) ;
 assign wire1132 = ( _575 ) | ( wire615  &  _9211 ) ;
 assign wire1134 = ( i_3_  &  i_2_  &  n_n592 ) ;
 assign wire6978 = ( wire1135 ) | ( n_n432  &  wire6976 ) ;
 assign wire6979 = ( wire1133 ) | ( (~ i_8_)  &  i_3_  &  n_n656 ) ;
 assign n_n1191 = ( wire1132 ) | ( wire1134 ) | ( wire6978 ) | ( wire6979 ) ;
 assign wire1154 = ( (~ i_7_)  &  (~ i_3_)  &  i_4_  &  _9176 ) ;
 assign wire6966 = ( wire1156 ) | ( (~ i_3_)  &  wire1162 ) | ( (~ i_3_)  &  wire6964 ) ;
 assign wire351 = ( (~ i_9_)  &  i_7_  &  i_4_ ) ;
 assign wire369 = ( (~ i_10_)  &  (~ i_13_)  &  i_4_  &  i_11_ ) ;
 assign wire617 = ( n_n816  &  wire9 ) | ( wire19  &  wire294 ) ;
 assign wire616 = ( n_n761  &  wire351 ) | ( (~ i_11_)  &  n_n761  &  n_n275 ) ;
 assign wire314 = ( i_9_  &  i_10_  &  i_7_ ) ;
 assign wire275 = ( (~ i_7_)  &  (~ i_2_) ) ;
 assign wire356 = ( i_8_  &  i_12_  &  (~ i_11_) ) ;
 assign wire619 = ( n_n35  &  n_n656 ) | ( wire275  &  wire356 ) ;
 assign n_n612 = ( i_5_  &  i_1_  &  i_2_ ) ;
 assign wire626 = ( i_10_  &  (~ i_7_)  &  (~ i_11_) ) | ( i_10_  &  (~ i_7_)  &  i_2_ ) ;
 assign wire628 = ( (~ i_8_)  &  wire37 ) | ( (~ i_8_)  &  (~ i_3_)  &  n_n716 ) ;
 assign wire633 = ( (~ i_8_)  &  (~ i_3_) ) | ( (~ i_7_)  &  (~ i_2_) ) ;
 assign wire632 = ( n_n566  &  wire19 ) | ( n_n741  &  wire633 ) ;
 assign wire7129 = ( n_n712  &  n_n751 ) | ( n_n570  &  n_n827 ) ;
 assign wire7127 = ( i_7_  &  (~ i_3_)  &  i_4_  &  (~ i_0_) ) ;
 assign wire638 = ( n_n545  &  wire377 ) | ( n_n755  &  wire7127 ) ;
 assign wire7126 = ( (~ i_5_)  &  (~ i_3_)  &  (~ i_0_) ) ;
 assign wire637 = ( n_n185  &  n_n683 ) | ( n_n752  &  wire7126 ) ;
 assign wire41 = ( (~ i_6_)  &  (~ i_3_)  &  (~ i_0_) ) | ( (~ i_3_)  &  (~ i_1_)  &  (~ i_0_) ) ;
 assign wire382 = ( (~ i_10_)  &  (~ i_7_)  &  (~ i_8_)  &  (~ i_11_) ) ;
 assign wire641 = ( (~ i_6_)  &  (~ i_0_)  &  n_n242 ) | ( i_6_  &  (~ i_0_)  &  n_n277 ) ;
 assign wire324 = ( (~ i_5_)  &  (~ i_3_)  &  (~ i_1_) ) ;
 assign wire1064 = ( (~ i_11_)  &  wire7017 ) | ( (~ i_11_)  &  wire7018 ) ;
 assign wire7019 = ( (~ i_5_)  &  wire265  &  n_n242 ) | ( i_5_  &  wire265  &  n_n277 ) ;
 assign wire649 = ( (~ i_8_)  &  i_11_ ) | ( i_9_  &  i_7_  &  i_11_ ) ;
 assign wire1848 = ( i_9_  &  i_10_  &  i_1_  &  i_11_ ) ;
 assign wire1849 = ( i_3_  &  i_1_  &  i_11_  &  i_2_ ) ;
 assign wire299 = ( i_12_  &  i_2_ ) ;
 assign wire316 = ( i_10_  &  (~ i_7_)  &  i_12_ ) ;
 assign wire395 = ( i_9_  &  i_5_  &  i_6_  &  i_12_ ) ;
 assign wire304 = ( i_10_  &  (~ i_5_)  &  (~ i_6_)  &  i_11_ ) ;
 assign wire384 = ( (~ i_5_)  &  (~ i_6_)  &  i_3_  &  i_2_ ) ;
 assign wire385 = ( (~ i_5_)  &  (~ i_6_)  &  i_2_ ) ;
 assign wire347 = ( i_10_  &  (~ i_5_) ) ;
 assign wire657 = ( i_0_  &  wire33  &  wire10 ) | ( (~ i_0_)  &  wire33  &  wire7184 ) ;
 assign wire777 = ( n_n752  &  wire338 ) | ( n_n752  &  wire779 ) ;
 assign wire7185 = ( n_n638  &  wire7182 ) | ( n_n651  &  wire7183 ) ;
 assign wire655 = ( wire777 ) | ( wire7185 ) | ( i_8_  &  wire657 ) ;
 assign wire772 = ( i_10_  &  (~ i_5_)  &  n_n346  &  wire356 ) ;
 assign wire773 = ( wire296  &  wire7181 ) ;
 assign n_n991 = ( wire772 ) | ( wire773 ) | ( (~ i_4_)  &  wire655 ) ;
 assign wire660 = ( i_9_  &  i_10_  &  i_11_ ) | ( i_9_  &  i_7_  &  i_11_ ) ;
 assign wire1814 = ( (~ i_7_)  &  wire1820 ) | ( (~ i_7_)  &  wire1821 ) ;
 assign wire6506 = ( wire6504 ) | ( (~ i_7_)  &  i_2_  &  wire304 ) ;
 assign wire6507 = ( wire1816 ) | ( wire1817 ) | ( wire385  &  wire660 ) ;
 assign wire287 = ( i_7_  &  i_3_  &  i_1_  &  i_0_ ) ;
 assign wire1805 = ( n_n598  &  wire1810 ) | ( n_n598  &  wire6510 ) ;
 assign wire1806 = ( i_12_  &  i_11_ ) | ( i_11_  &  wire327 ) | ( i_11_  &  wire123 ) ;
 assign wire1808 = ( i_12_  &  wire287 ) ;
 assign wire6512 = ( n_n36  &  wire388 ) | ( n_n35  &  wire6509 ) ;
 assign wire668 = ( (~ i_5_)  &  (~ i_6_)  &  (~ i_3_) ) | ( (~ i_5_)  &  (~ i_3_)  &  (~ i_1_) ) ;
 assign wire667 = ( n_n779  &  wire288 ) | ( n_n685  &  wire30 ) ;
 assign wire7066 = ( (~ i_5_)  &  i_4_  &  (~ i_1_) ) ;
 assign wire666 = ( n_n699  &  n_n710 ) | ( n_n792  &  wire7066 ) ;
 assign wire1074 = ( (~ i_9_)  &  i_5_  &  (~ i_6_)  &  (~ i_1_) ) ;
 assign wire7013 = ( i_5_  &  (~ i_3_)  &  (~ i_1_) ) ;
 assign wire669 = ( wire1074 ) | ( n_n658  &  n_n275 ) | ( n_n275  &  wire7013 ) ;
 assign wire671 = ( wire35  &  n_n675 ) | ( n_n672  &  wire11 ) ;
 assign wire406 = ( (~ i_9_)  &  i_8_  &  i_5_  &  _9853 ) ;
 assign wire677 = ( (~ i_5_)  &  (~ i_6_) ) | ( (~ i_6_)  &  (~ i_0_) ) ;
 assign wire676 = ( wire279  &  n_n671 ) | ( n_n792  &  wire677 ) ;
 assign wire403 = ( (~ i_3_)  &  i_4_  &  (~ i_1_)  &  _8395 ) ;
 assign wire334 = ( i_9_  &  i_12_  &  i_11_ ) ;
 assign wire380 = ( (~ i_11_)  &  (~ i_0_) ) ;
 assign wire686 = ( n_n432  &  n_n176 ) | ( wire12  &  wire270 ) ;
 assign wire685 = ( i_5_  &  wire292 ) | ( i_5_  &  (~ i_12_)  &  n_n814 ) ;
 assign wire373 = ( _372 ) | ( wire689  &  _9409 ) ;
 assign wire7191 = ( wire362 ) | ( n_n818  &  wire686 ) ;
 assign n_n993 = ( wire373 ) | ( wire7191 ) | ( wire18  &  wire685 ) ;
 assign wire1012 = ( _520 ) | ( n_n827  &  _9280 ) ;
 assign wire7046 = ( n_n741  &  _9285 ) | ( (~ i_7_)  &  (~ i_2_)  &  n_n741 ) ;
 assign wire7047 = ( n_n242  &  n_n606 ) | ( n_n624  &  n_n277 ) ;
 assign wire1003 = ( i_6_  &  (~ i_1_)  &  (~ i_0_) ) | ( i_6_  &  (~ i_0_)  &  wire1009 ) ;
 assign wire1005 = ( (~ i_3_)  &  (~ i_2_)  &  (~ i_0_)  &  _9303 ) ;
 assign wire7050 = ( i_5_  &  (~ i_0_) ) | ( n_n835  &  _9304 ) ;
 assign wire7051 = ( n_n769  &  n_n671 ) | ( n_n240  &  wire698 ) ;
 assign wire696 = ( wire1003 ) | ( wire1005 ) | ( wire7050 ) | ( wire7051 ) ;
 assign wire397 = ( i_9_  &  i_5_  &  (~ i_6_)  &  i_11_ ) ;
 assign wire701 = ( i_9_  &  i_7_  &  i_6_ ) | ( i_9_  &  i_7_  &  i_11_ ) ;
 assign wire7269 = ( i_9_  &  i_3_  &  i_12_  &  i_1_ ) ;
 assign wire700 = ( n_n432  &  n_n826 ) | ( wire380  &  wire7269 ) ;
 assign wire704 = ( i_5_  &  (~ i_6_)  &  i_3_ ) | ( i_5_  &  i_3_  &  i_1_ ) ;
 assign wire366 = ( i_5_  &  i_3_  &  i_0_ ) ;
 assign wire7275 = ( (~ i_7_)  &  i_8_  &  i_5_ ) ;
 assign wire703 = ( n_n746  &  wire366 ) | ( n_n826  &  wire7275 ) ;
 assign wire706 = ( i_10_  &  (~ i_5_) ) | ( (~ i_5_)  &  (~ i_0_) ) ;
 assign wire707 = ( (~ i_5_)  &  i_0_ ) | ( i_5_  &  (~ i_12_)  &  (~ i_0_) ) ;
 assign wire7294 = ( (~ i_7_)  &  (~ i_8_)  &  (~ i_0_) ) ;
 assign wire7295 = ( i_5_  &  i_3_  &  (~ i_12_)  &  i_1_ ) ;
 assign wire7296 = ( (~ i_7_)  &  (~ i_8_)  &  (~ i_6_)  &  i_3_ ) ;
 assign wire705 = ( wire7294  &  wire7295 ) | ( wire707  &  wire7296 ) ;
 assign wire7178 = ( i_9_  &  i_5_ ) ;
 assign wire708 = ( n_n538  &  wire333 ) | ( n_n369  &  wire7178 ) ;
 assign wire785 = ( _310 ) | ( wire712  &  _9492 ) ;
 assign wire718 = ( i_9_  &  i_0_ ) | ( (~ i_5_)  &  i_0_ ) ;
 assign wire717 = ( wire20  &  wire334 ) | ( n_n415  &  wire718 ) ;
 assign wire719 = ( i_10_  &  i_12_  &  (~ i_11_) ) | ( i_10_  &  i_12_  &  i_0_ ) | ( i_12_  &  (~ i_11_)  &  (~ i_0_) ) ;
 assign wire7194 = ( i_5_  &  i_6_  &  i_0_ ) ;
 assign wire716 = ( n_n176  &  wire719 ) | ( wire270  &  wire7194 ) ;
 assign wire256 = ( (~ i_4_)  &  i_2_  &  wire716 ) ;
 assign wire7196 = ( wire255 ) | ( wire258 ) | ( (~ i_4_)  &  wire717 ) ;
 assign wire762 = ( wire863 ) | ( wire864 ) | ( n_n716  &  wire763 ) ;
 assign wire857 = ( i_5_  &  (~ i_6_)  &  wire761 ) ;
 assign wire7140 = ( wire405 ) | ( wire856 ) | ( wire859 ) ;
 assign n_n981 = ( wire857 ) | ( wire7140 ) | ( i_5_  &  wire762 ) ;
 assign wire836 = ( n_n853  &  wire51 ) | ( n_n853  &  n_n671  &  n_n810 ) ;
 assign wire7155 = ( wire834 ) | ( wire835 ) | ( wire17  &  wire6669 ) ;
 assign wire824 = ( n_n853  &  wire7157 ) | ( n_n764  &  n_n853  &  n_n791 ) ;
 assign wire825 = ( (~ i_10_)  &  (~ i_6_)  &  wire17  &  n_n671 ) ;
 assign wire7161 = ( wire68 ) | ( wire69 ) | ( wire106 ) | ( wire120 ) ;
 assign wire726 = ( (~ i_7_) ) | ( (~ i_8_)  &  (~ i_3_) ) ;
 assign wire725 = ( n_n773  &  n_n671 ) | ( n_n835  &  wire726 ) ;
 assign wire724 = ( wire37 ) | ( (~ i_3_)  &  n_n725 ) ;
 assign wire7165 = ( (~ i_10_)  &  (~ i_8_)  &  (~ i_13_)  &  i_12_ ) ;
 assign wire723 = ( wire37  &  n_n671 ) | ( n_n771  &  wire7165 ) ;
 assign wire374 = ( i_9_  &  (~ i_4_)  &  i_11_ ) ;
 assign wire246 = ( wire304  &  wire7200 ) | ( wire397  &  wire7200 ) ;
 assign wire247 = ( (~ i_7_)  &  i_5_  &  n_n826  &  wire374 ) ;
 assign wire249 = ( _301 ) | ( (~ i_8_)  &  i_5_  &  wire7203 ) ;
 assign wire808 = ( (~ i_9_)  &  i_8_  &  (~ i_13_)  &  (~ i_12_) ) ;
 assign wire809 = ( (~ i_9_)  &  (~ i_8_)  &  (~ i_13_)  &  (~ i_11_) ) ;
 assign wire735 = ( wire24 ) | ( wire808 ) | ( wire809 ) ;
 assign wire10 = ( i_9_  &  i_10_  &  i_12_ ) | ( i_10_  &  (~ i_5_)  &  i_12_ ) ;
 assign wire737 = ( wire395 ) | ( wire397 ) | ( i_6_  &  wire10 ) ;
 assign wire263 = ( i_6_  &  (~ i_0_) ) ;
 assign wire230 = ( i_1_  &  (~ i_11_)  &  i_2_  &  (~ i_0_) ) ;
 assign wire231 = ( i_10_  &  i_1_  &  i_2_  &  i_0_ ) ;
 assign wire7219 = ( i_12_  &  (~ i_11_)  &  i_2_ ) ;
 assign wire736 = ( wire230 ) | ( wire231 ) | ( wire263  &  wire7219 ) ;
 assign wire7226 = ( (~ i_5_)  &  i_12_  &  (~ i_11_)  &  (~ i_0_) ) ;
 assign wire738 = ( n_n818  &  wire304 ) | ( n_n752  &  wire7226 ) ;
 assign wire746 = ( i_13_  &  (~ i_12_) ) | ( (~ i_13_)  &  i_4_  &  i_12_ ) ;
 assign wire751 = ( (~ i_5_)  &  i_6_  &  i_3_ ) | ( (~ i_5_)  &  i_3_  &  i_1_ ) ;
 assign wire54 = ( (~ i_5_)  &  (~ i_11_) ) | ( (~ i_12_)  &  (~ i_11_) ) ;
 assign wire80 = ( i_5_  &  (~ i_12_)  &  i_1_  &  i_2_ ) ;
 assign wire81 = ( i_5_  &  i_1_  &  i_2_  &  i_0_ ) ;
 assign wire752 = ( wire80 ) | ( wire81 ) | ( n_n840  &  wire54 ) ;
 assign wire763 = ( n_n792  &  n_n683 ) | ( n_n699  &  wire7136 ) ;
 assign wire863 = ( wire37  &  wire7134 ) ;
 assign wire864 = ( (~ i_7_)  &  (~ i_8_)  &  n_n849  &  n_n791 ) ;
 assign wire7132 = ( (~ i_10_)  &  (~ i_7_)  &  (~ i_13_)  &  i_12_ ) ;
 assign wire7133 = ( (~ i_1_)  &  (~ i_0_) ) ;
 assign wire761 = ( n_n678  &  wire7132 ) | ( n_n716  &  wire7133 ) ;
 assign wire51 = ( n_n769  &  n_n771 ) | ( n_n835  &  wire318 ) ;
 assign wire317 = ( i_8_  &  (~ i_5_)  &  (~ i_6_)  &  (~ i_3_) ) ;
 assign wire319 = ( (~ i_9_)  &  i_8_  &  (~ i_13_)  &  i_4_ ) ;
 assign wire329 = ( (~ i_10_)  &  (~ i_13_)  &  (~ i_12_)  &  (~ i_11_) ) ;
 assign wire335 = ( (~ i_9_)  &  (~ i_13_)  &  (~ i_12_)  &  (~ i_11_) ) ;
 assign wire424 = ( n_n850  &  n_n751 ) | ( n_n570  &  n_n503 ) ;
 assign wire6549 = ( i_9_  &  i_8_  &  (~ i_6_) ) ;
 assign wire6550 = ( i_9_  &  (~ i_7_)  &  i_8_  &  (~ i_6_) ) ;
 assign wire423 = ( wire329  &  wire6549 ) | ( n_n729  &  wire6550 ) ;
 assign wire429 = ( i_6_  &  (~ i_0_) ) | ( (~ i_1_)  &  (~ i_0_) ) ;
 assign wire428 = ( i_6_  &  i_0_ ) | ( i_1_  &  i_0_ ) ;
 assign wire426 = ( i_5_  &  i_1_  &  i_2_ ) | ( i_1_  &  i_2_  &  i_0_ ) ;
 assign wire1740 = ( i_5_  &  (~ i_1_)  &  (~ i_2_) ) ;
 assign wire1741 = ( i_6_  &  (~ i_2_)  &  (~ i_0_) ) ;
 assign wire440 = ( (~ i_9_)  &  i_7_  &  i_8_ ) | ( (~ i_10_)  &  (~ i_7_)  &  (~ i_8_) ) ;
 assign wire447 = ( i_1_  &  wire335 ) | ( (~ i_13_)  &  i_1_  &  n_n277 ) ;
 assign wire452 = ( i_5_  &  (~ i_6_)  &  (~ i_13_) ) | ( i_5_  &  (~ i_13_)  &  i_1_ ) ;
 assign wire451 = ( n_n816  &  wire264 ) | ( n_n822  &  wire452 ) ;
 assign wire459 = ( wire279  &  wire301 ) | ( n_n852  &  wire329 ) ;
 assign wire469 = ( n_n658  &  n_n844 ) | ( n_n847  &  n_n653 ) ;
 assign wire468 = ( i_5_  &  (~ i_6_)  &  n_n838 ) | ( (~ i_5_)  &  i_6_  &  n_n830 ) ;
 assign wire479 = ( n_n852  &  n_n846 ) | ( n_n847  &  n_n851 ) ;
 assign wire6622 = ( i_8_  &  (~ i_3_)  &  i_0_ ) ;
 assign wire6623 = ( i_8_  &  i_1_ ) ;
 assign wire515 = ( i_6_  &  (~ i_12_) ) | ( (~ i_12_)  &  (~ i_11_) ) ;
 assign wire531 = ( i_7_ ) | ( i_8_  &  (~ i_3_) ) ;
 assign wire530 = ( wire23  &  n_n729 ) | ( n_n575  &  wire531 ) ;
 assign wire541 = ( (~ i_5_)  &  n_n833  &  wire277 ) | ( i_5_  &  n_n830  &  wire277 ) ;
 assign wire551 = ( (~ i_5_)  &  i_6_  &  n_n838 ) | ( i_5_  &  (~ i_6_)  &  n_n830 ) ;
 assign wire569 = ( n_n795  &  n_n570 ) | ( n_n843  &  n_n751 ) ;
 assign wire576 = ( i_5_  &  (~ i_6_)  &  i_2_ ) | ( i_5_  &  i_1_  &  i_2_ ) ;
 assign wire6803 = ( i_5_  &  i_3_  &  (~ i_4_)  &  (~ i_12_) ) ;
 assign wire615 = ( i_10_  &  i_7_  &  (~ i_8_) ) | ( i_10_  &  (~ i_8_)  &  (~ i_11_) ) ;
 assign wire622 = ( i_2_ ) | ( (~ i_12_)  &  (~ i_11_) ) ;
 assign wire636 = ( (~ i_10_)  &  (~ i_7_)  &  (~ i_11_) ) | ( (~ i_10_)  &  (~ i_12_)  &  (~ i_11_) ) ;
 assign wire635 = ( (~ i_10_)  &  (~ i_7_)  &  i_8_ ) | ( (~ i_10_)  &  (~ i_7_)  &  (~ i_11_) ) ;
 assign wire644 = ( (~ i_9_)  &  (~ i_8_)  &  i_6_ ) | ( (~ i_10_)  &  (~ i_8_)  &  (~ i_6_) ) ;
 assign wire643 = ( (~ i_7_) ) | ( (~ i_8_)  &  (~ i_3_) ) ;
 assign wire646 = ( i_6_  &  (~ i_3_)  &  (~ i_0_) ) | ( (~ i_3_)  &  (~ i_1_)  &  (~ i_0_) ) ;
 assign wire653 = ( i_8_  &  i_12_ ) | ( i_10_  &  (~ i_7_)  &  i_12_ ) ;
 assign wire7184 = ( (~ i_5_)  &  i_12_  &  (~ i_11_) ) ;
 assign wire673 = ( i_8_  &  (~ i_3_) ) | ( i_7_  &  (~ i_2_) ) ;
 assign wire680 = ( (~ i_9_)  &  i_7_  &  i_8_ ) | ( (~ i_10_)  &  (~ i_7_)  &  i_8_ ) ;
 assign wire684 = ( i_9_  &  i_7_  &  i_8_ ) | ( i_9_  &  i_7_  &  i_6_ ) ;
 assign wire1794 = ( i_9_  &  i_7_  &  i_6_  &  i_2_ ) ;
 assign wire683 = ( n_n814 ) | ( wire1794 ) | ( i_1_  &  wire684 ) ;
 assign wire7190 = ( i_9_  &  i_12_  &  (~ i_11_) ) ;
 assign wire689 = ( (~ i_5_)  &  i_0_  &  n_n432 ) | ( (~ i_5_)  &  (~ i_0_)  &  wire7190 ) ;
 assign wire698 = ( (~ i_5_)  &  (~ i_6_)  &  (~ i_3_) ) | ( (~ i_5_)  &  (~ i_3_)  &  (~ i_1_) ) ;
 assign wire712 = ( n_n541  &  wire333 ) | ( n_n369  &  wire347 ) ;
 assign wire728 = ( (~ i_9_)  &  i_4_ ) | ( (~ i_8_)  &  i_4_ ) ;
 assign wire734 = ( n_n819  &  wire381 ) | ( n_n752  &  n_n550 ) ;
 assign wire741 = ( i_9_  &  i_7_  &  i_8_ ) | ( i_7_  &  i_8_  &  (~ i_5_) ) ;
 assign wire7136 = ( (~ i_2_)  &  (~ i_0_) ) ;
 assign wire7322 = ( (~ i_8_)  &  (~ i_5_)  &  i_4_ ) ;
 assign wire57 = ( (~ i_7_)  &  (~ i_5_)  &  wire1202 ) | ( (~ i_7_)  &  (~ i_5_)  &  wire1203 ) ;
 assign wire7325 = ( (~ i_7_)  &  (~ i_8_)  &  (~ i_5_) ) ;
 assign wire59 = ( n_n699  &  wire62 ) | ( n_n699  &  wire63 ) ;
 assign wire60 = ( (~ i_1_)  &  wire329 ) ;
 assign wire7327 = ( wire325  &  n_n575 ) | ( wire281  &  wire7326 ) ;
 assign wire1202 = ( (~ i_10_)  &  i_8_  &  (~ i_13_)  &  (~ i_12_) ) ;
 assign wire1203 = ( (~ i_10_)  &  (~ i_13_)  &  i_4_ ) ;
 assign wire62 = ( (~ i_3_)  &  (~ i_13_)  &  (~ i_12_)  &  (~ i_11_) ) ;
 assign wire63 = ( (~ i_13_)  &  (~ i_11_)  &  (~ i_2_) ) ;
 assign wire82 = ( i_7_  &  i_12_  &  i_2_ ) ;
 assign wire83 = ( i_8_  &  i_3_  &  i_12_ ) ;
 assign wire7312 = ( i_9_  &  i_10_  &  i_11_  &  i_0_ ) ;
 assign wire64 = ( wire82  &  wire7312 ) | ( wire83  &  wire7312 ) ;
 assign wire84 = ( (~ i_5_)  &  i_12_  &  (~ i_11_)  &  (~ i_0_) ) ;
 assign wire7313 = ( i_9_  &  i_7_  &  i_6_  &  i_2_ ) ;
 assign wire65 = ( wire338  &  wire7313 ) | ( wire84  &  wire7313 ) ;
 assign wire86 = ( i_12_  &  (~ i_11_)  &  n_n597  &  wire751 ) ;
 assign wire95 = ( (~ i_5_)  &  i_1_  &  i_2_  &  i_0_ ) ;
 assign wire89 = ( wire126  &  wire95 ) | ( wire126  &  n_n526  &  n_n840 ) ;
 assign wire7304 = ( i_10_  &  i_11_  &  (~ i_0_) ) ;
 assign wire103 = ( i_9_  &  i_10_  &  i_13_  &  i_0_ ) ;
 assign wire107 = ( i_10_  &  (~ i_5_)  &  i_13_  &  i_0_ ) ;
 assign wire112 = ( i_9_  &  i_5_  &  i_13_  &  (~ i_12_) ) ;
 assign wire7280 = ( i_10_  &  (~ i_8_)  &  i_3_ ) ;
 assign wire127 = ( i_5_  &  (~ i_12_)  &  n_n840  &  wire7280 ) ;
 assign wire7282 = ( (~ i_7_)  &  (~ i_8_)  &  (~ i_5_) ) ;
 assign wire128 = ( i_10_  &  i_11_  &  n_n826  &  wire7282 ) ;
 assign wire136 = ( i_10_  &  (~ i_8_)  &  i_2_ ) ;
 assign wire129 = ( n_n631  &  n_n316  &  wire314 ) | ( n_n631  &  n_n316  &  wire136 ) ;
 assign wire130 = ( i_9_  &  i_10_  &  n_n639  &  wire354 ) ;
 assign wire144 = ( i_5_  &  (~ i_6_)  &  (~ i_12_)  &  i_2_ ) ;
 assign wire145 = ( i_5_  &  (~ i_6_)  &  i_2_  &  i_0_ ) ;
 assign wire139 = ( n_n194  &  wire144 ) | ( n_n194  &  wire145 ) ;
 assign wire141 = ( i_9_  &  i_5_  &  i_13_  &  i_0_ ) ;
 assign wire142 = ( i_5_  &  i_13_  &  (~ i_12_)  &  (~ i_0_) ) ;
 assign wire143 = ( i_13_  &  (~ i_12_)  &  (~ i_11_)  &  (~ i_0_) ) ;
 assign wire7264 = ( i_9_  &  i_8_  &  i_2_ ) ;
 assign wire150 = ( (~ i_12_)  &  i_11_  &  n_n639  &  wire7264 ) ;
 assign wire156 = ( i_5_  &  i_3_  &  i_11_  &  i_0_ ) ;
 assign wire154 = ( wire270  &  wire156 ) | ( n_n826  &  wire34  &  wire270 ) ;
 assign wire163 = ( i_9_  &  i_10_  &  i_1_  &  i_0_ ) ;
 assign wire166 = ( i_5_  &  (~ i_6_)  &  (~ i_12_)  &  i_2_ ) ;
 assign wire180 = ( (~ i_5_)  &  i_6_  &  i_12_  &  i_2_ ) ;
 assign wire182 = ( (~ i_5_)  &  i_1_  &  i_2_ ) ;
 assign wire190 = ( i_3_  &  i_0_  &  wire104 ) | ( i_2_  &  i_0_  &  wire104 ) ;
 assign wire194 = ( i_9_  &  i_10_  &  i_5_  &  (~ i_12_) ) ;
 assign wire1408 = ( i_9_  &  i_10_  &  (~ i_5_)  &  (~ i_11_) ) ;
 assign wire1409 = ( i_9_  &  i_10_  &  (~ i_12_)  &  (~ i_11_) ) ;
 assign wire192 = ( i_1_  &  wire194 ) | ( i_1_  &  wire1408 ) | ( i_1_  &  wire1409 ) ;
 assign wire7235 = ( i_5_  &  (~ i_6_)  &  (~ i_12_)  &  i_11_ ) ;
 assign wire198 = ( wire7235  &  _9528 ) | ( wire7235  &  _9529 ) ;
 assign wire200 = ( (~ i_8_)  &  i_5_  &  n_n598  &  wire374 ) ;
 assign wire207 = ( wire27  &  wire208 ) | ( wire27  &  wire841 ) | ( wire27  &  wire842 ) ;
 assign wire201 = ( _292 ) | ( (~ i_4_)  &  i_1_  &  wire207 ) ;
 assign wire7239 = ( i_5_  &  (~ i_12_)  &  i_11_ ) ;
 assign wire208 = ( i_9_  &  i_5_  &  i_11_  &  i_0_ ) ;
 assign wire841 = ( i_5_  &  (~ i_12_)  &  i_11_  &  (~ i_0_) ) ;
 assign wire842 = ( i_10_  &  (~ i_5_)  &  i_11_  &  i_0_ ) ;
 assign wire7223 = ( (~ i_12_)  &  i_11_  &  i_2_ ) ;
 assign wire212 = ( (~ i_6_)  &  (~ i_0_)  &  n_n538  &  wire7223 ) ;
 assign wire213 = ( i_5_  &  (~ i_6_)  &  n_n412  &  wire342 ) ;
 assign wire222 = ( i_12_  &  (~ i_11_)  &  wire223 ) | ( i_12_  &  (~ i_11_)  &  wire224 ) ;
 assign wire7229 = ( wire741  &  wire7227 ) | ( wire270  &  wire7228 ) ;
 assign wire215 = ( (~ i_4_)  &  i_1_  &  wire222 ) | ( (~ i_4_)  &  i_1_  &  wire7229 ) ;
 assign wire223 = ( i_10_  &  i_7_  &  i_8_  &  (~ i_5_) ) ;
 assign wire224 = ( i_7_  &  i_8_  &  (~ i_5_)  &  (~ i_0_) ) ;
 assign wire7215 = ( i_10_  &  i_12_  &  (~ i_11_) ) ;
 assign wire225 = ( (~ i_5_)  &  i_6_  &  n_n412  &  wire7215 ) ;
 assign wire7208 = ( i_10_  &  i_12_  &  (~ i_11_) ) | ( i_12_  &  (~ i_11_)  &  (~ i_0_) ) ;
 assign wire235 = ( i_7_  &  i_6_  &  n_n541  &  wire7208 ) ;
 assign wire236 = ( i_10_  &  i_12_  &  n_n153  &  wire591 ) ;
 assign wire241 = ( i_9_  &  i_5_  &  (~ i_12_) ) ;
 assign wire237 = ( wire360  &  wire272 ) | ( wire272  &  wire241 ) ;
 assign wire238 = ( i_1_  &  i_2_  &  i_0_  &  wire307 ) ;
 assign wire253 = ( i_5_  &  i_3_  &  (~ i_4_)  &  (~ i_0_) ) ;
 assign wire7199 = ( (~ i_7_)  &  (~ i_6_)  &  (~ i_12_)  &  i_11_ ) ;
 assign wire245 = ( wire307  &  wire7199 ) | ( wire253  &  wire7199 ) ;
 assign wire7200 = ( (~ i_7_)  &  i_3_  &  (~ i_4_)  &  i_0_ ) ;
 assign wire7203 = ( n_n346  &  wire342 ) | ( wire297  &  n_n840 ) ;
 assign wire255 = ( i_9_  &  i_12_  &  n_n752  &  wire366 ) ;
 assign wire6976 = ( i_8_  &  (~ i_4_)  &  i_2_ ) ;
 assign wire258 = ( i_6_  &  i_0_  &  n_n432  &  wire6976 ) ;
 assign wire7188 = ( i_9_  &  i_3_  &  i_12_  &  i_2_ ) ;
 assign wire362 = ( (~ i_11_)  &  (~ i_0_)  &  n_n176  &  wire7188 ) ;
 assign wire768 = ( i_9_  &  i_8_  &  (~ i_12_)  &  (~ i_11_) ) ;
 assign wire769 = ( i_9_  &  i_8_  &  (~ i_5_)  &  (~ i_11_) ) ;
 assign wire7181 = ( i_9_  &  i_8_  &  i_5_  &  i_12_ ) ;
 assign wire779 = ( i_9_  &  i_5_  &  i_12_  &  i_0_ ) ;
 assign wire790 = ( i_9_  &  i_7_  &  i_5_  &  i_12_ ) ;
 assign wire791 = ( i_10_  &  (~ i_7_)  &  (~ i_5_)  &  i_11_ ) ;
 assign wire798 = ( i_7_  &  i_0_  &  n_n658  &  wire24 ) ;
 assign wire7175 = ( i_5_  &  (~ i_6_)  &  (~ i_1_)  &  i_0_ ) ;
 assign wire800 = ( (~ i_9_)  &  (~ i_13_)  &  (~ i_11_)  &  wire7175 ) ;
 assign wire802 = ( (~ i_1_)  &  wire335 ) | ( (~ i_1_)  &  wire286  &  wire24 ) ;
 assign wire801 = ( wire20  &  wire802 ) | ( (~ i_3_)  &  wire20  &  wire734 ) ;
 assign wire814 = ( n_n853  &  n_n819  &  n_n678 ) ;
 assign wire7157 = ( n_n773  &  n_n771 ) | ( n_n683  &  wire351 ) ;
 assign wire834 = ( i_5_  &  (~ i_6_)  &  n_n581  &  wire297 ) ;
 assign wire835 = ( i_6_  &  (~ i_0_)  &  n_n764  &  wire17 ) ;
 assign wire843 = ( (~ i_5_)  &  (~ i_0_)  &  n_n819  &  wire301 ) ;
 assign wire844 = ( wire284  &  n_n671  &  n_n176 ) ;
 assign wire850 = ( wire35  &  wire853 ) | ( wire35  &  wire854 ) | ( wire35  &  wire855 ) ;
 assign wire852 = ( i_4_  &  (~ i_1_)  &  (~ i_0_)  &  _9615 ) ;
 assign wire7146 = ( n_n176  &  n_n771 ) | ( n_n671  &  wire7144 ) ;
 assign wire845 = ( n_n755  &  wire850 ) | ( n_n755  &  wire852 ) | ( n_n755  &  wire7146 ) ;
 assign wire7138 = ( (~ i_5_)  &  (~ i_1_)  &  (~ i_2_)  &  (~ i_0_) ) ;
 assign wire853 = ( i_8_  &  (~ i_1_)  &  (~ i_2_)  &  (~ i_0_) ) ;
 assign wire854 = ( i_7_  &  i_8_  &  i_6_  &  (~ i_0_) ) ;
 assign wire855 = ( i_7_  &  (~ i_3_)  &  (~ i_1_)  &  (~ i_0_) ) ;
 assign wire856 = ( (~ i_7_)  &  i_5_  &  wire37  &  n_n683 ) ;
 assign wire859 = ( i_8_  &  (~ i_3_)  &  n_n545  &  wire7138 ) ;
 assign wire7134 = ( (~ i_8_)  &  (~ i_1_)  &  (~ i_2_)  &  (~ i_0_) ) ;
 assign wire7119 = ( i_5_  &  (~ i_3_)  &  i_0_ ) ;
 assign wire7121 = ( i_5_  &  i_6_  &  (~ i_1_)  &  i_0_ ) ;
 assign wire7015 = ( (~ i_9_)  &  (~ i_8_)  &  i_5_ ) ;
 assign wire887 = ( i_5_  &  i_6_  &  wire346 ) | ( i_5_  &  i_6_  &  wire891 ) ;
 assign wire7122 = ( n_n675  &  n_n813 ) | ( n_n277  &  wire7011 ) ;
 assign wire891 = ( (~ i_9_)  &  i_7_  &  i_8_  &  i_4_ ) ;
 assign wire895 = ( _25 ) | ( n_n816  &  _9867 ) ;
 assign wire905 = ( i_7_  &  (~ i_5_)  &  (~ i_1_)  &  (~ i_2_) ) ;
 assign wire7109 = ( i_8_  &  (~ i_13_)  &  (~ i_12_)  &  i_11_ ) ;
 assign wire907 = ( (~ i_10_)  &  (~ i_5_)  &  n_n675  &  wire7109 ) ;
 assign wire912 = ( i_4_  &  (~ i_2_)  &  wire322 ) ;
 assign wire7110 = ( n_n819  &  n_n712 ) | ( n_n764  &  wire7033 ) ;
 assign wire7111 = ( n_n685  &  n_n827 ) | ( n_n624  &  n_n277 ) ;
 assign wire909 = ( n_n761  &  wire912 ) | ( n_n761  &  wire7110 ) | ( n_n761  &  wire7111 ) ;
 assign wire917 = ( n_n545  &  n_n240  &  wire668 ) ;
 assign wire7094 = ( (~ i_9_)  &  (~ i_13_)  &  (~ i_11_) ) ;
 assign wire934 = ( (~ i_9_)  &  (~ i_7_)  &  (~ i_13_)  &  (~ i_11_) ) ;
 assign wire7100 = ( i_5_  &  i_6_  &  (~ i_2_)  &  i_0_ ) ;
 assign wire927 = ( wire319  &  wire7100 ) | ( wire335  &  wire7100 ) | ( wire934  &  wire7100 ) ;
 assign wire954 = ( i_0_  &  wire957 ) | ( i_0_  &  wire958 ) ;
 assign wire7084 = ( wire11  &  n_n670 ) | ( n_n843  &  wire16 ) ;
 assign wire7085 = ( (~ i_10_)  &  (~ i_13_)  &  i_4_ ) ;
 assign wire7086 = ( (~ i_10_)  &  (~ i_8_)  &  (~ i_13_)  &  (~ i_11_) ) ;
 assign wire948 = ( (~ i_5_)  &  (~ i_6_)  &  n_n670  &  wire7086 ) ;
 assign wire957 = ( (~ i_8_)  &  (~ i_5_)  &  (~ i_6_)  &  (~ i_2_) ) ;
 assign wire958 = ( (~ i_7_)  &  (~ i_5_)  &  (~ i_6_)  &  (~ i_3_) ) ;
 assign wire7078 = ( (~ i_10_)  &  (~ i_13_)  &  (~ i_12_)  &  i_0_ ) ;
 assign wire7080 = ( n_n842  &  n_n710 ) | ( wire30  &  wire7079 ) ;
 assign wire961 = ( n_n838  &  wire7080 ) | ( (~ i_5_)  &  n_n838  &  wire530 ) ;
 assign wire7068 = ( i_5_  &  i_6_  &  (~ i_3_)  &  (~ i_12_) ) ;
 assign wire972 = ( _411 ) | ( n_n624  &  _9364 ) ;
 assign wire995 = ( (~ i_10_)  &  (~ i_7_)  &  (~ i_12_)  &  (~ i_11_) ) ;
 assign wire987 = ( n_n653  &  wire382 ) | ( n_n653  &  wire995 ) ;
 assign wire988 = ( (~ i_5_)  &  (~ i_11_)  &  (~ i_0_) ) | ( (~ i_12_)  &  (~ i_11_)  &  (~ i_0_) ) ;
 assign wire993 = ( (~ i_9_)  &  (~ i_3_) ) | ( (~ i_9_)  &  (~ i_2_) ) ;
 assign wire1009 = ( (~ i_9_)  &  i_7_  &  i_8_  &  (~ i_3_) ) ;
 assign wire1021 = ( i_7_  &  (~ i_5_)  &  (~ i_1_)  &  (~ i_2_) ) ;
 assign wire1026 = ( i_5_  &  i_6_  &  i_4_ ) | ( i_6_  &  i_4_  &  (~ i_0_) ) ;
 assign wire1027 = ( i_5_  &  (~ i_3_)  &  (~ i_12_)  &  (~ i_1_) ) ;
 assign wire1023 = ( n_n764  &  wire1026 ) | ( n_n764  &  wire1027 ) ;
 assign wire1030 = ( (~ i_3_)  &  (~ i_1_)  &  (~ i_2_)  &  _9290 ) ;
 assign wire7042 = ( n_n675  &  n_n768 ) | ( wire267  &  n_n624 ) ;
 assign wire7043 = ( (~ wire55)  &  wire322 ) | ( wire317  &  wire7041 ) ;
 assign wire1024 = ( (~ i_12_)  &  wire1030 ) | ( (~ i_12_)  &  wire7042 ) | ( (~ i_12_)  &  wire7043 ) ;
 assign wire1040 = ( (~ i_6_)  &  (~ i_0_)  &  wire1043 ) | ( (~ i_6_)  &  (~ i_0_)  &  wire1044 ) ;
 assign wire1041 = ( (~ i_3_)  &  (~ i_1_)  &  (~ i_0_)  &  wire680 ) ;
 assign wire7035 = ( wire1042 ) | ( (~ i_2_)  &  (~ i_0_)  &  n_n819 ) ;
 assign wire1033 = ( (~ i_12_)  &  wire1040 ) | ( (~ i_12_)  &  wire1041 ) | ( (~ i_12_)  &  wire7035 ) ;
 assign wire1043 = ( (~ i_10_)  &  i_7_  &  (~ i_2_) ) ;
 assign wire1044 = ( (~ i_10_)  &  (~ i_7_)  &  i_8_  &  (~ i_3_) ) ;
 assign wire1042 = ( i_7_  &  (~ i_1_)  &  (~ i_2_)  &  (~ i_0_) ) ;
 assign wire1047 = ( (~ i_9_)  &  (~ i_10_)  &  i_4_ ) ;
 assign wire7017 = ( wire1067 ) | ( n_n675  &  wire7015 ) ;
 assign wire7018 = ( wire1074 ) | ( n_n275  &  wire7013 ) | ( n_n275  &  wire646 ) ;
 assign wire1067 = ( (~ i_10_)  &  (~ i_5_)  &  (~ i_6_)  &  (~ i_1_) ) ;
 assign wire1082 = ( (~ i_6_)  &  (~ i_1_)  &  (~ i_0_) ) ;
 assign wire1089 = ( (~ i_8_)  &  wire1092 ) | ( (~ i_8_)  &  wire1093 ) ;
 assign wire7004 = ( wire1087 ) | ( (~ i_7_)  &  (~ i_5_)  &  n_n685 ) ;
 assign wire7005 = ( wire35  &  n_n675 ) | ( n_n683  &  wire7003 ) ;
 assign wire1083 = ( (~ i_10_)  &  wire1089 ) | ( (~ i_10_)  &  wire7004 ) | ( (~ i_10_)  &  wire7005 ) ;
 assign wire1087 = ( (~ i_5_)  &  i_6_  &  (~ i_12_)  &  (~ i_1_) ) ;
 assign wire1092 = ( i_4_  &  (~ i_1_)  &  (~ i_2_)  &  (~ i_0_) ) ;
 assign wire1093 = ( (~ i_5_)  &  i_4_  &  (~ i_1_)  &  (~ i_2_) ) ;
 assign wire6994 = ( (~ i_3_)  &  (~ i_13_)  &  (~ i_12_)  &  i_2_ ) ;
 assign wire1094 = ( (~ i_9_)  &  i_7_  &  i_8_  &  wire6994 ) ;
 assign wire6996 = ( n_n787  &  n_n672 ) | ( n_n755  &  wire6995 ) ;
 assign wire1103 = ( i_2_  &  wire319 ) | ( (~ i_3_)  &  i_2_  &  wire335 ) ;
 assign wire1115 = ( i_10_  &  (~ i_7_)  &  i_8_  &  i_12_ ) ;
 assign wire1116 = ( i_9_  &  i_10_  &  (~ i_8_)  &  i_11_ ) ;
 assign wire1117 = ( i_9_  &  i_7_  &  i_8_  &  i_12_ ) ;
 assign wire1108 = ( wire14  &  wire1115 ) | ( wire14  &  wire1116 ) | ( wire14  &  wire1117 ) ;
 assign wire1119 = ( i_9_  &  i_10_  &  (~ i_7_)  &  (~ i_11_) ) ;
 assign wire1109 = ( i_3_  &  wire1119 ) | ( i_3_  &  wire8  &  wire622 ) ;
 assign wire1110 = ( i_3_  &  (~ i_12_)  &  wire314 ) ;
 assign wire1130 = ( i_9_  &  i_7_  &  i_8_  &  (~ i_12_) ) ;
 assign wire6983 = ( n_n623  &  wire275 ) | ( n_n526  &  wire6982 ) ;
 assign wire1121 = ( i_3_  &  wire1130 ) | ( i_3_  &  wire6983 ) ;
 assign wire1122 = ( i_9_  &  i_10_  &  i_13_  &  i_2_ ) ;
 assign wire1123 = ( (~ i_7_)  &  i_13_  &  (~ i_11_)  &  (~ i_2_) ) ;
 assign wire1133 = ( i_9_  &  i_7_  &  i_13_  &  i_2_ ) ;
 assign wire1135 = ( i_7_  &  i_13_  &  (~ i_12_)  &  (~ i_2_) ) ;
 assign wire1152 = ( (~ i_9_)  &  (~ i_3_)  &  (~ i_13_)  &  i_4_ ) ;
 assign wire6967 = ( i_7_  &  i_2_ ) ;
 assign wire1139 = ( wire1152  &  wire6967 ) | ( wire23  &  n_n719  &  wire6967 ) ;
 assign wire1143 = ( (~ i_7_)  &  (~ i_8_)  &  wire369 ) ;
 assign wire1160 = ( (~ i_10_)  &  (~ i_7_)  &  (~ i_8_)  &  i_4_ ) ;
 assign wire1156 = ( (~ i_13_)  &  wire1160 ) | ( (~ i_13_)  &  n_n566  &  wire19 ) ;
 assign wire1162 = ( (~ i_7_)  &  wire329 ) ;
 assign wire1166 = ( (~ i_10_)  &  (~ i_12_)  &  (~ i_11_)  &  _9185 ) ;
 assign wire1171 = ( (~ i_9_)  &  i_8_  &  i_4_  &  (~ i_2_) ) ;
 assign wire1168 = ( n_n853  &  n_n672 ) | ( n_n853  &  wire1171 ) ;
 assign wire1173 = ( i_9_  &  i_7_  &  (~ i_12_) ) | ( i_7_  &  (~ i_12_)  &  (~ i_2_) ) ;
 assign wire1175 = ( (~ i_12_)  &  (~ i_11_)  &  (~ i_2_) ) ;
 assign wire6959 = ( i_10_  &  (~ i_7_)  &  (~ i_11_) ) | ( (~ i_7_)  &  (~ i_11_)  &  (~ i_2_) ) ;
 assign wire1169 = ( wire21  &  wire1173 ) | ( wire21  &  wire1175 ) | ( wire21  &  wire6959 ) ;
 assign wire1180 = ( i_9_  &  i_7_  &  i_12_  &  i_11_ ) ;
 assign wire1181 = ( i_10_  &  (~ i_7_)  &  (~ i_8_)  &  i_11_ ) ;
 assign wire1182 = ( i_9_  &  i_7_  &  (~ i_8_)  &  i_11_ ) ;
 assign wire1183 = ( i_10_  &  (~ i_7_)  &  i_12_  &  i_11_ ) ;
 assign wire6945 = ( wire635  &  wire6942 ) | ( n_n575  &  wire6944 ) ;
 assign wire1194 = ( (~ i_13_)  &  (~ i_11_)  &  n_n273  &  n_n773 ) ;
 assign wire1348 = ( (~ i_10_)  &  (~ i_7_)  &  (~ i_6_)  &  (~ i_3_) ) ;
 assign wire1196 = ( wire336  &  wire371 ) | ( wire371  &  wire1348 ) ;
 assign wire1200 = ( (~ i_3_)  &  (~ i_13_)  &  i_1_  &  (~ i_11_) ) ;
 assign wire1204 = ( (~ i_6_)  &  (~ i_11_)  &  wire298 ) ;
 assign wire1213 = ( i_12_  &  wire393 ) ;
 assign wire6920 = ( i_6_  &  (~ i_4_)  &  i_1_  &  i_2_ ) ;
 assign wire1218 = ( i_9_  &  i_8_  &  i_12_  &  wire6920 ) ;
 assign wire1228 = ( (~ i_4_)  &  i_2_  &  wire1229 ) | ( (~ i_4_)  &  i_2_  &  wire1230 ) ;
 assign wire6925 = ( n_n651  &  wire6923 ) | ( n_n346  &  wire6924 ) ;
 assign wire1229 = ( i_8_  &  i_12_  &  (~ i_1_)  &  (~ i_11_) ) ;
 assign wire1230 = ( i_10_  &  i_8_  &  i_12_  &  (~ i_11_) ) ;
 assign wire1239 = ( i_9_  &  i_10_  &  (~ i_6_)  &  (~ i_11_) ) ;
 assign wire1234 = ( i_2_  &  wire1239 ) | ( i_2_  &  wire8  &  wire515 ) ;
 assign wire1235 = ( i_9_  &  i_10_  &  i_1_  &  i_2_ ) ;
 assign wire1245 = ( n_n534  &  _9028 ) | ( n_n534  &  _9029 ) ;
 assign wire1249 = ( (~ i_7_)  &  i_6_  &  i_3_  &  (~ i_12_) ) ;
 assign wire1250 = ( (~ i_7_)  &  i_3_  &  i_1_ ) ;
 assign wire1246 = ( n_n421  &  wire1249 ) | ( n_n421  &  wire1250 ) ;
 assign wire1252 = ( i_6_  &  i_3_  &  i_12_  &  i_1_ ) ;
 assign wire6908 = ( (~ i_6_)  &  i_3_  &  (~ i_1_) ) ;
 assign wire1247 = ( n_n638  &  wire1252 ) | ( n_n638  &  n_n316  &  wire6908 ) ;
 assign wire1248 = ( i_3_  &  i_1_  &  i_11_  &  wire364 ) ;
 assign wire6897 = ( i_6_  &  i_3_  &  (~ i_1_) ) ;
 assign wire1255 = ( (~ i_12_)  &  i_11_  &  n_n592  &  wire6897 ) ;
 assign wire1266 = ( i_10_  &  i_3_  &  i_1_  &  i_2_ ) ;
 assign wire1272 = ( i_10_  &  (~ i_6_)  &  i_12_  &  i_11_ ) ;
 assign wire1267 = ( (~ i_4_)  &  i_1_  &  wire104 ) | ( (~ i_4_)  &  i_1_  &  wire1272 ) ;
 assign wire1277 = ( i_3_  &  (~ i_4_)  &  (~ i_12_)  &  i_2_ ) ;
 assign wire1279 = ( (~ i_12_)  &  (~ i_1_)  &  i_2_  &  wire493 ) ;
 assign wire1290 = ( i_9_  &  i_10_  &  i_7_  &  i_12_ ) ;
 assign wire6887 = ( n_n748  &  n_n197 ) | ( n_n638  &  wire6886 ) ;
 assign wire6875 = ( (~ i_8_)  &  i_6_  &  (~ i_4_)  &  i_2_ ) ;
 assign wire6876 = ( i_9_  &  (~ i_12_)  &  i_11_ ) | ( (~ i_12_)  &  (~ i_1_)  &  i_11_ ) ;
 assign wire1301 = ( i_9_  &  i_10_  &  (~ i_7_)  &  (~ i_8_) ) ;
 assign wire1302 = ( i_9_  &  (~ i_7_)  &  (~ i_8_)  &  i_6_ ) ;
 assign wire6879 = ( (~ i_4_)  &  i_1_  &  i_11_ ) ;
 assign wire1297 = ( (~ i_7_)  &  (~ i_8_)  &  i_6_  &  (~ i_1_) ) ;
 assign wire1298 = ( i_9_  &  (~ i_7_)  &  (~ i_8_)  &  i_6_ ) ;
 assign wire1299 = ( i_10_  &  (~ i_8_)  &  (~ i_6_)  &  i_11_ ) ;
 assign wire1300 = ( i_9_  &  (~ i_8_)  &  i_6_  &  i_11_ ) ;
 assign wire1307 = ( i_6_  &  i_13_  &  (~ i_12_)  &  (~ i_1_) ) ;
 assign wire1308 = ( i_13_  &  (~ i_12_)  &  (~ i_1_)  &  (~ i_11_) ) ;
 assign wire1314 = ( (~ i_10_)  &  (~ i_3_)  &  n_n545  &  n_n746 ) ;
 assign wire6864 = ( (~ i_10_)  &  i_8_  &  (~ i_6_)  &  (~ i_3_) ) ;
 assign wire1321 = ( (~ i_9_)  &  i_7_  &  i_8_  &  i_6_ ) ;
 assign wire1338 = ( (~ i_9_)  &  i_7_  &  i_6_  &  (~ i_3_) ) ;
 assign wire1339 = ( (~ i_9_)  &  i_8_  &  i_6_  &  (~ i_2_) ) ;
 assign wire1317 = ( wire295  &  wire1321 ) | ( wire295  &  wire1338 ) | ( wire295  &  wire1339 ) ;
 assign wire1324 = ( (~ i_13_)  &  (~ i_12_)  &  i_11_  &  _9139 ) ;
 assign wire1331 = ( (~ i_9_)  &  i_6_  &  (~ i_13_)  &  i_4_ ) ;
 assign wire1326 = ( n_n273  &  wire1331 ) | ( n_n273  &  n_n274  &  n_n503 ) ;
 assign wire1328 = ( (~ i_3_)  &  (~ i_2_)  &  n_n716  &  n_n503 ) ;
 assign wire1329 = ( wire371  &  wire1338 ) | ( wire371  &  wire1339 ) ;
 assign wire1334 = ( (~ i_3_)  &  (~ i_13_)  &  (~ i_12_)  &  i_1_ ) ;
 assign wire1336 = ( (~ i_9_)  &  (~ i_7_)  &  (~ i_2_) ) ;
 assign wire1337 = ( (~ i_9_)  &  i_7_  &  (~ i_8_)  &  (~ i_3_) ) ;
 assign wire6852 = ( (~ i_3_)  &  i_1_ ) | ( i_1_  &  (~ i_2_) ) ;
 assign wire1340 = ( (~ i_9_)  &  (~ i_13_)  &  n_n701  &  wire6852 ) ;
 assign wire6853 = ( (~ i_8_)  &  i_6_  &  (~ i_3_) ) ;
 assign wire1341 = ( (~ i_13_)  &  i_12_  &  n_n741  &  wire6853 ) ;
 assign wire1346 = ( (~ i_10_)  &  (~ i_7_)  &  (~ i_8_)  &  (~ i_6_) ) ;
 assign wire1343 = ( wire336  &  wire370 ) | ( wire370  &  wire1348 ) | ( wire370  &  wire1346 ) ;
 assign wire1361 = ( (~ i_3_)  &  i_4_  &  (~ i_1_)  &  (~ i_2_) ) ;
 assign wire6842 = ( n_n779  &  wire309 ) | ( n_n685  &  wire267 ) ;
 assign wire6843 = ( (~ i_6_)  &  (~ i_13_)  &  i_11_ ) ;
 assign wire1350 = ( wire1361  &  wire6843 ) | ( wire6842  &  wire6843 ) ;
 assign wire1351 = ( (~ i_3_)  &  i_1_  &  n_n819  &  wire381 ) ;
 assign wire1352 = ( (~ i_13_)  &  (~ i_12_)  &  n_n769  &  n_n273 ) ;
 assign wire1353 = ( _666 ) | ( i_6_  &  (~ i_2_)  &  wire447 ) ;
 assign wire6846 = ( (~ i_3_)  &  (~ i_13_)  &  i_1_  &  (~ i_11_) ) ;
 assign wire6835 = ( i_7_  &  (~ i_6_)  &  (~ i_1_)  &  (~ i_2_) ) ;
 assign wire1372 = ( n_n764  &  wire1373 ) | ( n_n764  &  n_n545  &  wire31 ) ;
 assign wire6838 = ( i_8_  &  (~ i_13_)  &  (~ i_12_)  &  i_11_ ) ;
 assign wire1373 = ( (~ i_13_)  &  i_4_  &  (~ i_1_)  &  i_11_ ) ;
 assign wire1383 = ( (~ i_7_)  &  (~ i_1_)  &  (~ i_2_) ) ;
 assign wire6831 = ( i_6_  &  (~ i_13_)  &  i_12_  &  (~ i_11_) ) ;
 assign wire1377 = ( wire17  &  n_n675 ) | ( (~ i_1_)  &  wire17  &  wire440 ) ;
 assign wire1385 = ( _870 ) | ( _871 ) ;
 assign wire1393 = ( i_5_  &  i_6_  &  i_3_  &  i_2_ ) ;
 assign wire1394 = ( i_5_  &  i_3_  &  i_1_  &  i_2_ ) ;
 assign wire1388 = ( n_n665  &  wire287 ) | ( n_n665  &  wire1393 ) | ( n_n665  &  wire1394 ) ;
 assign wire1390 = ( i_13_  &  wire292 ) ;
 assign wire6816 = ( i_6_  &  (~ i_13_)  &  (~ i_12_)  &  i_11_ ) ;
 assign wire1397 = ( (~ i_7_)  &  (~ i_5_)  &  i_3_  &  i_1_ ) ;
 assign wire1406 = ( i_13_  &  (~ i_11_)  &  wire327 ) | ( i_13_  &  (~ i_11_)  &  wire384 ) ;
 assign wire6812 = ( wire272  &  wire276 ) | ( n_n818  &  wire6811 ) ;
 assign wire1403 = ( wire272  &  wire1408 ) | ( wire272  &  wire1409 ) ;
 assign wire6794 = ( (~ i_5_)  &  (~ i_6_)  &  (~ i_11_) ) ;
 assign wire1410 = ( n_n592  &  wire272  &  wire6794 ) ;
 assign wire6799 = ( (~ i_9_)  &  (~ i_2_) ) ;
 assign wire6785 = ( (~ i_13_)  &  i_4_  &  (~ i_1_)  &  i_0_ ) ;
 assign wire1423 = ( n_n795  &  n_n822  &  wire6785 ) ;
 assign wire1432 = ( n_n822  &  wire24  &  wire576 ) ;
 assign wire1433 = ( n_n816  &  wire42  &  wire9 ) | ( n_n816  &  wire9  &  wire6788 ) ;
 assign wire1425 = ( (~ i_8_)  &  wire1432 ) | ( (~ i_8_)  &  wire1433 ) ;
 assign wire6788 = ( (~ i_5_)  &  (~ i_6_)  &  i_2_ ) | ( (~ i_6_)  &  i_2_  &  i_0_ ) ;
 assign wire1436 = ( n_n846  &  n_n822  &  _8588 ) ;
 assign wire6776 = ( i_6_  &  i_3_  &  i_2_ ) ;
 assign wire1437 = ( (~ i_9_)  &  i_4_  &  wire313  &  wire6776 ) ;
 assign wire1440 = ( (~ i_9_)  &  i_4_  &  n_n816  &  wire359 ) ;
 assign wire1441 = ( wire292  &  wire340 ) ;
 assign wire1446 = ( (~ i_9_)  &  i_3_  &  i_4_  &  i_0_ ) ;
 assign wire1447 = ( (~ i_9_)  &  (~ i_5_)  &  i_3_  &  i_4_ ) ;
 assign wire1450 = ( n_n844  &  n_n843  &  n_n842  &  n_n851 ) ;
 assign wire6770 = ( n_n850  &  n_n852 ) | ( n_n838  &  n_n837 ) ;
 assign wire6771 = ( n_n835  &  n_n837 ) | ( n_n843  &  n_n840 ) ;
 assign wire6772 = ( n_n850  &  n_n847 ) | ( n_n830  &  n_n832 ) ;
 assign wire6762 = ( i_7_  &  i_6_  &  i_3_ ) ;
 assign wire6763 = ( i_5_  &  (~ i_6_)  &  i_3_  &  i_2_ ) ;
 assign wire1464 = ( wire327  &  n_n816  &  wire9 ) | ( n_n816  &  wire9  &  wire384 ) ;
 assign wire6764 = ( n_n819  &  n_n846 ) | ( n_n814  &  n_n813 ) ;
 assign wire1472 = ( n_n850  &  n_n725  &  n_n852  &  n_n735 ) ;
 assign wire1474 = ( (~ i_8_)  &  (~ i_3_)  &  n_n741  &  wire521 ) ;
 assign wire1480 = ( (~ i_8_)  &  i_6_  &  (~ i_3_)  &  i_0_ ) ;
 assign wire1481 = ( (~ i_8_)  &  i_5_  &  i_6_  &  (~ i_3_) ) ;
 assign wire1488 = ( n_n849  &  n_n844  &  wire318 ) ;
 assign wire1493 = ( i_5_  &  (~ i_1_)  &  wire17 ) | ( i_5_  &  i_1_  &  wire37 ) ;
 assign wire6749 = ( wire295  &  wire12 ) | ( n_n853  &  n_n791 ) ;
 assign wire6750 = ( i_6_  &  (~ i_0_)  &  wire17 ) | ( i_6_  &  i_0_  &  wire37 ) ;
 assign wire1500 = ( n_n844  &  n_n751  &  n_n752  &  n_n846 ) ;
 assign wire1501 = ( (~ i_2_)  &  wire17  &  wire322 ) ;
 assign wire1502 = ( i_1_  &  i_0_  &  n_n764  &  wire37 ) ;
 assign wire6719 = ( (~ i_5_)  &  i_4_  &  i_1_ ) ;
 assign wire1524 = ( n_n816  &  n_n795  &  wire6719 ) ;
 assign wire1525 = ( wire420  &  wire24  &  _8633 ) ;
 assign wire1526 = ( (~ i_5_)  &  wire17  &  wire336 ) ;
 assign wire1527 = ( i_2_  &  wire37  &  wire322 ) ;
 assign wire1528 = ( (~ i_8_)  &  (~ i_5_)  &  n_n779  &  wire313 ) ;
 assign wire6725 = ( i_8_  &  i_1_  &  i_2_ ) ;
 assign wire1529 = ( (~ i_9_)  &  i_4_  &  wire313  &  wire6725 ) ;
 assign wire1530 = ( n_n853  &  n_n773  &  n_n771 ) ;
 assign wire1534 = ( n_n795  &  n_n498  &  wire13  &  wire298 ) ;
 assign wire6714 = ( n_n358  &  wire6712 ) | ( wire34  &  wire6713 ) ;
 assign wire6708 = ( i_10_  &  (~ i_7_)  &  (~ i_8_)  &  i_6_ ) ;
 assign wire1552 = ( i_7_  &  i_8_  &  n_n658  &  n_n835 ) ;
 assign wire1553 = ( n_n833  &  n_n653  &  n_n651 ) ;
 assign wire6698 = ( (~ i_5_)  &  (~ i_6_)  &  (~ i_3_) ) | ( (~ i_5_)  &  (~ i_3_)  &  (~ i_1_) ) ;
 assign wire1554 = ( n_n656  &  wire41 ) | ( n_n656  &  wire6698 ) ;
 assign wire1562 = ( (~ i_9_)  &  i_7_  &  wire313  &  n_n685 ) ;
 assign wire6686 = ( (~ i_3_)  &  (~ i_1_)  &  (~ i_2_)  &  i_0_ ) ;
 assign wire1563 = ( n_n822  &  wire24  &  wire6686 ) ;
 assign wire6687 = ( n_n819  &  n_n678 ) | ( n_n819  &  n_n712 ) ;
 assign wire6688 = ( n_n699  &  n_n710 ) | ( n_n683  &  wire351 ) ;
 assign wire1564 = ( n_n853  &  wire403 ) | ( n_n853  &  wire6687 ) | ( n_n853  &  wire6688 ) ;
 assign wire1565 = ( (~ i_10_)  &  (~ i_5_)  &  wire17  &  n_n675 ) ;
 assign wire1574 = ( (~ i_7_)  &  (~ i_6_)  &  (~ i_3_)  &  i_0_ ) ;
 assign wire1575 = ( (~ i_7_)  &  (~ i_3_)  &  (~ i_1_)  &  i_0_ ) ;
 assign wire1569 = ( n_n822  &  wire24  &  wire1574 ) | ( n_n822  &  wire24  &  wire1575 ) ;
 assign wire1571 = ( (~ i_7_)  &  (~ i_5_)  &  wire313  &  n_n685 ) ;
 assign wire1572 = ( n_n835  &  n_n761  &  n_n712  &  n_n752 ) ;
 assign wire1587 = ( (~ i_5_)  &  (~ i_6_)  &  (~ i_3_)  &  (~ i_2_) ) ;
 assign wire1588 = ( (~ i_6_)  &  (~ i_3_)  &  (~ i_2_)  &  (~ i_0_) ) ;
 assign wire6670 = ( i_10_  &  i_13_  &  (~ i_12_)  &  (~ i_11_) ) ;
 assign wire1582 = ( wire1587  &  wire6670 ) | ( wire1588  &  wire6670 ) ;
 assign wire6672 = ( (~ i_6_)  &  (~ i_3_)  &  (~ i_2_)  &  i_0_ ) ;
 assign wire1583 = ( n_n822  &  wire24  &  wire6672 ) ;
 assign wire6674 = ( n_n671  &  n_n810 ) | ( n_n675  &  n_n813 ) ;
 assign wire6675 = ( n_n672  &  wire6673 ) | ( n_n672  &  _8369 ) ;
 assign wire1585 = ( (~ i_10_)  &  (~ i_6_)  &  wire17  &  n_n671 ) ;
 assign wire1596 = ( n_n835  &  n_n787  &  n_n843  &  n_n710 ) ;
 assign wire1611 = ( n_n835  &  n_n716  &  n_n732  &  n_n837 ) ;
 assign wire1620 = ( (~ i_7_)  &  (~ i_8_)  &  (~ i_6_)  &  _8482 ) ;
 assign wire6647 = ( i_7_  &  (~ i_8_)  &  i_1_ ) ;
 assign wire6636 = ( (~ i_3_)  &  (~ i_1_)  &  (~ i_2_)  &  (~ i_0_) ) ;
 assign wire1639 = ( i_6_  &  (~ i_3_)  &  (~ i_2_)  &  (~ i_0_) ) ;
 assign wire1640 = ( i_5_  &  i_6_  &  (~ i_3_)  &  (~ i_2_) ) ;
 assign wire1644 = ( i_5_  &  (~ i_3_)  &  (~ i_1_) ) ;
 assign wire6630 = ( n_n852  &  wire6628 ) | ( n_n847  &  wire6629 ) ;
 assign wire6631 = ( i_10_  &  (~ i_7_)  &  i_13_  &  (~ i_12_) ) ;
 assign wire6563 = ( (~ i_7_)  &  i_13_  &  (~ i_11_) ) ;
 assign wire6632 = ( i_13_  &  i_1_  &  i_2_  &  i_0_ ) ;
 assign wire1661 = ( n_n566  &  wire296  &  _8728 ) ;
 assign wire1663 = ( n_n746  &  wire294  &  n_n735 ) ;
 assign wire1672 = ( n_n716  &  n_n847  &  wire307  &  n_n756 ) ;
 assign wire1673 = ( n_n844  &  n_n752  &  n_n550  &  n_n732 ) ;
 assign wire1675 = ( n_n835  &  n_n545  &  n_n746  &  n_n735 ) ;
 assign wire6595 = ( i_8_  &  (~ i_3_)  &  (~ i_4_) ) ;
 assign wire1684 = ( wire344  &  wire6594  &  n_n598  &  wire6595 ) ;
 assign wire1685 = ( n_n746  &  n_n844  &  n_n575  &  n_n735 ) ;
 assign wire6603 = ( wire1689 ) | ( wire1691 ) | ( wire469  &  wire6600 ) ;
 assign wire1686 = ( _941 ) | ( i_13_  &  (~ i_11_)  &  wire6603 ) ;
 assign wire6598 = ( (~ i_8_)  &  (~ i_5_)  &  (~ i_3_) ) ;
 assign wire1689 = ( n_n358  &  n_n840  &  wire6598 ) ;
 assign wire1691 = ( (~ i_7_)  &  (~ i_8_)  &  n_n835  &  n_n653 ) ;
 assign wire1704 = ( i_13_  &  (~ i_12_)  &  (~ i_1_)  &  (~ i_0_) ) ;
 assign wire1705 = ( (~ i_5_)  &  (~ i_6_)  &  i_13_ ) ;
 assign wire6588 = ( i_10_  &  (~ i_7_)  &  (~ i_8_)  &  (~ i_11_) ) ;
 assign wire1699 = ( wire1704  &  wire6588 ) | ( wire1705  &  wire6588 ) ;
 assign wire6589 = ( (~ i_7_)  &  (~ i_5_)  &  (~ i_1_) ) ;
 assign wire6578 = ( i_9_  &  i_5_ ) ;
 assign wire6579 = ( (~ i_3_)  &  i_13_  &  (~ i_11_) ) ;
 assign wire1708 = ( n_n832  &  n_n852  &  wire6578  &  wire6579 ) ;
 assign wire6582 = ( i_13_  &  i_1_  &  i_2_  &  i_0_ ) ;
 assign wire1709 = ( n_n635  &  n_n592  &  wire6582 ) ;
 assign wire6584 = ( (~ i_0_)  &  n_n633  &  wire265 ) | ( i_0_  &  n_n631  &  wire265 ) ;
 assign wire6585 = ( n_n631  &  n_n852 ) | ( n_n639  &  n_n840 ) ;
 assign wire1720 = ( (~ i_11_)  &  wire341  &  n_n752  &  n_n840 ) ;
 assign wire1724 = ( n_n570  &  n_n847  &  n_n541  &  n_n752 ) ;
 assign wire1725 = ( n_n835  &  n_n570  &  n_n541  &  n_n756 ) ;
 assign wire1722 = ( i_9_  &  i_11_  &  wire1724 ) | ( i_9_  &  i_11_  &  wire1725 ) ;
 assign wire1726 = ( (~ i_5_)  &  i_6_  &  wire294  &  wire298 ) ;
 assign wire6573 = ( i_3_  &  (~ i_4_)  &  (~ i_12_)  &  (~ i_11_) ) ;
 assign wire1729 = ( wire6573  &  _8824 ) ;
 assign wire1732 = ( i_9_  &  i_8_  &  wire434  &  wire6563 ) ;
 assign wire6558 = ( (~ i_7_)  &  (~ i_5_)  &  i_1_ ) | ( (~ i_7_)  &  i_1_  &  i_0_ ) ;
 assign wire6559 = ( i_9_  &  i_10_  &  i_8_  &  i_2_ ) ;
 assign wire1748 = ( (~ i_6_)  &  (~ i_2_)  &  (~ i_0_) ) ;
 assign wire1750 = ( (~ i_7_)  &  (~ i_6_)  &  (~ i_0_) ) ;
 assign wire1763 = ( n_n838  &  n_n748  &  n_n725  &  wire341 ) ;
 assign wire1764 = ( n_n835  &  n_n538  &  n_n850  &  n_n498 ) ;
 assign wire1767 = ( n_n538  &  n_n725  &  n_n830  &  n_n746 ) ;
 assign wire1768 = ( n_n835  &  n_n538  &  n_n748  &  n_n716 ) ;
 assign wire1765 = ( i_9_  &  wire1767 ) | ( i_9_  &  wire1768 ) ;
 assign wire1770 = ( wire341  &  n_n575  &  n_n756 ) ;
 assign wire1776 = ( i_9_  &  i_10_  &  i_1_ ) | ( i_10_  &  (~ i_6_)  &  i_1_ ) ;
 assign wire1778 = ( i_10_  &  (~ i_7_)  &  i_2_ ) ;
 assign wire1779 = ( i_9_  &  i_6_  &  i_1_ ) ;
 assign wire1780 = ( i_9_  &  i_10_  &  i_3_ ) | ( i_9_  &  i_10_  &  i_2_ ) ;
 assign wire1781 = ( i_9_  &  i_8_  &  i_3_ ) ;
 assign wire1792 = ( i_9_  &  i_10_  &  i_12_  &  i_1_ ) ;
 assign wire1803 = ( (~ i_8_)  &  i_1_  &  i_11_  &  i_0_ ) ;
 assign wire1804 = ( i_3_  &  i_1_  &  i_11_  &  i_0_ ) ;
 assign wire1796 = ( (~ i_7_)  &  wire1803 ) | ( (~ i_7_)  &  wire1804 ) ;
 assign wire6515 = ( i_10_  &  (~ i_7_) ) | ( (~ i_8_)  &  i_11_ ) ;
 assign wire6516 = ( i_9_  &  i_7_ ) | ( i_8_  &  i_12_ ) ;
 assign wire1797 = ( n_n844  &  wire6515 ) | ( n_n844  &  wire6516 ) ;
 assign wire1798 = ( i_10_  &  (~ i_6_)  &  i_1_  &  i_0_ ) ;
 assign wire6509 = ( i_7_  &  i_1_  &  i_0_ ) ;
 assign wire1810 = ( i_10_  &  (~ i_7_)  &  i_11_ ) ;
 assign wire6510 = ( (~ i_8_)  &  i_11_ ) | ( i_9_  &  i_7_  &  i_11_ ) ;
 assign wire1820 = ( (~ i_8_)  &  (~ i_5_)  &  (~ i_6_)  &  i_11_ ) ;
 assign wire1821 = ( (~ i_5_)  &  (~ i_6_)  &  i_3_  &  i_11_ ) ;
 assign wire1816 = ( i_9_  &  i_6_  &  i_1_  &  i_0_ ) ;
 assign wire1817 = ( i_9_  &  i_10_  &  i_0_ ) ;
 assign wire1829 = ( i_7_  &  i_8_  &  i_12_ ) | ( i_7_  &  i_3_  &  i_12_ ) ;
 assign wire6493 = ( i_8_  &  i_12_ ) | ( i_9_  &  i_10_  &  i_12_ ) ;
 assign wire6494 = ( i_5_  &  i_6_  &  i_2_ ) ;
 assign wire1838 = ( i_8_  &  i_5_  &  i_6_  &  i_12_ ) ;
 assign wire1839 = ( i_5_  &  i_6_  &  i_3_  &  i_12_ ) ;
 assign wire1844 = ( i_10_  &  i_1_  &  i_11_  &  i_2_ ) ;
 assign wire1845 = ( (~ i_8_)  &  i_1_  &  i_11_ ) ;
 assign wire1850 = ( i_9_  &  i_10_  &  i_3_  &  i_13_ ) ;
 assign wire1856 = ( i_9_  &  i_8_  &  (~ i_12_) ) | ( i_8_  &  (~ i_3_)  &  (~ i_12_) ) ;
 assign wire1857 = ( i_9_  &  i_10_  &  (~ i_12_)  &  (~ i_11_) ) ;
 assign wire1853 = ( (~ i_8_)  &  (~ i_3_)  &  i_13_  &  (~ i_11_) ) ;
 assign wire1863 = ( i_9_  &  i_8_  &  i_3_ ) ;
 assign wire6478 = ( i_10_  &  (~ i_8_)  &  i_3_ ) | ( i_10_  &  (~ i_8_)  &  (~ i_11_) ) ;
 assign wire6473 = ( (~ i_8_)  &  (~ i_11_) ) | ( (~ i_12_)  &  (~ i_11_) ) ;
 assign wire6488 = ( i_9_  &  i_1_  &  i_11_ ) ;
 assign wire6499 = ( i_12_  &  i_2_  &  i_0_ ) ;
 assign wire6504 = ( i_9_  &  i_5_  &  i_0_ ) | ( i_10_  &  (~ i_5_)  &  i_0_ ) ;
 assign wire6522 = ( i_7_  &  i_5_  &  i_3_  &  i_1_ ) ;
 assign wire6523 = ( i_5_  &  (~ i_6_)  &  i_1_ ) ;
 assign wire6524 = ( i_9_  &  i_7_  &  i_12_ ) ;
 assign wire6526 = ( i_12_  &  wire6522 ) | ( i_10_  &  i_12_  &  wire6523 ) ;
 assign wire6527 = ( wire376  &  wire334 ) | ( n_n612  &  wire6524 ) ;
 assign wire6554 = ( i_7_  &  i_5_  &  (~ i_1_) ) ;
 assign wire6567 = ( wire1732 ) | ( n_n665  &  wire425 ) | ( n_n665  &  wire435 ) ;
 assign wire6593 = ( wire1699 ) | ( _933 ) | ( _934 ) ;
 assign wire6600 = ( i_9_  &  i_7_  &  (~ i_8_) ) ;
 assign wire6605 = ( wire1684 ) | ( wire1685 ) | ( wire6593 ) | ( _930 ) ;
 assign wire6618 = ( i_7_  &  i_8_  &  (~ i_6_)  &  wire284 ) ;
 assign wire6620 = ( (~ i_3_)  &  (~ i_4_)  &  i_0_ ) ;
 assign wire6621 = ( i_8_  &  (~ i_5_)  &  (~ i_3_) ) ;
 assign wire6628 = ( i_8_  &  (~ i_5_)  &  i_6_  &  (~ i_3_) ) ;
 assign wire6629 = ( i_8_  &  i_5_  &  i_6_  &  (~ i_3_) ) ;
 assign wire6637 = ( i_9_  &  i_5_ ) ;
 assign wire6638 = ( (~ i_3_)  &  (~ i_0_) ) ;
 assign wire6643 = ( i_1_  &  i_2_  &  i_0_  &  _8457 ) ;
 assign wire6645 = ( (~ i_9_)  &  (~ i_10_)  &  (~ i_11_)  &  _8451 ) ;
 assign wire6653 = ( n_n832  &  n_n852 ) | ( n_n844  &  n_n837 ) ;
 assign wire6654 = ( i_5_  &  (~ i_3_)  &  i_4_  &  _8480 ) ;
 assign wire6660 = ( (~ i_7_)  &  i_8_  &  i_6_  &  _8492 ) ;
 assign wire6661 = ( (~ i_7_)  &  (~ i_8_)  &  i_6_  &  _8489 ) ;
 assign wire6665 = ( wire543  &  wire6660 ) | ( wire544  &  wire6661 ) ;
 assign wire6667 = ( wire1596 ) | ( wire6665 ) | ( n_n844  &  wire545 ) ;
 assign wire6673 = ( (~ i_10_)  &  (~ i_5_)  &  (~ i_6_) ) ;
 assign wire6693 = ( wire120 ) | ( wire1562 ) | ( wire1563 ) | ( wire1565 ) ;
 assign wire6712 = ( i_10_  &  i_3_  &  i_0_ ) ;
 assign wire6713 = ( i_9_  &  i_10_  &  i_3_  &  i_1_ ) ;
 assign wire6730 = ( wire68 ) | ( wire1524 ) | ( wire1528 ) | ( wire1530 ) ;
 assign wire6731 = ( wire1525 ) | ( wire1526 ) | ( wire1527 ) | ( wire1529 ) ;
 assign wire6757 = ( wire1472 ) | ( _1018 ) | ( _1019 ) ;
 assign wire6780 = ( wire1440 ) | ( wire1441 ) | ( n_n849  &  wire612 ) ;
 assign wire6787 = ( (~ i_10_)  &  (~ i_7_)  &  (~ i_13_)  &  i_11_ ) ;
 assign wire6789 = ( wire1423 ) | ( wire574  &  wire6787 ) ;
 assign wire6806 = ( wire1410 ) | ( _808 ) | ( _810 ) ;
 assign wire6811 = ( i_6_  &  i_13_  &  (~ i_12_) ) ;
 assign wire6850 = ( wire1351 ) | ( wire1352 ) | ( wire6848  &  _9093 ) ;
 assign wire6854 = ( (~ i_10_)  &  (~ i_6_)  &  (~ i_13_)  &  i_11_ ) ;
 assign wire6858 = ( wire1341 ) | ( wire1343 ) | ( n_n672  &  wire6854 ) ;
 assign wire6860 = ( wire1326 ) | ( wire1328 ) | ( wire1329 ) ;
 assign wire6865 = ( n_n816  &  wire9 ) | ( wire29  &  wire294 ) ;
 assign wire6868 = ( wire1317 ) | ( (~ i_6_)  &  wire1324 ) | ( (~ i_6_)  &  wire6865 ) ;
 assign wire6869 = ( wire1314 ) | ( wire6868 ) | ( _9141 ) ;
 assign wire6870 = ( wire6858 ) | ( wire6860 ) | ( _9168 ) ;
 assign wire6884 = ( i_10_  &  i_1_  &  i_2_ ) ;
 assign wire6885 = ( (~ i_6_)  &  i_2_ ) ;
 assign wire6886 = ( i_10_  &  (~ i_6_)  &  i_12_ ) ;
 assign wire6888 = ( wire28  &  wire6884 ) | ( n_n656  &  wire6885 ) ;
 assign wire6894 = ( wire272  &  wire311 ) | ( n_n412  &  wire363 ) ;
 assign wire6899 = ( i_3_  &  (~ i_12_)  &  (~ i_1_)  &  i_2_ ) ;
 assign wire6900 = ( i_9_  &  i_8_  &  i_6_  &  i_12_ ) ;
 assign wire6901 = ( i_3_  &  i_12_  &  i_1_ ) ;
 assign wire6904 = ( wire15  &  wire104 ) | ( i_11_  &  wire15  &  wire6900 ) ;
 assign wire6906 = ( i_9_  &  i_8_  &  i_6_ ) ;
 assign wire6911 = ( wire1245 ) | ( wire1247 ) | ( wire512  &  wire6906 ) ;
 assign wire6913 = ( i_7_  &  (~ i_6_)  &  i_3_  &  i_12_ ) ;
 assign wire6914 = ( i_9_  &  i_7_  &  (~ i_1_)  &  i_2_ ) ;
 assign wire6915 = ( wire1235 ) | ( n_n609  &  wire6913 ) ;
 assign wire6916 = ( n_n358  &  wire513 ) | ( wire516  &  wire6914 ) ;
 assign wire6918 = ( wire1234 ) | ( wire6915 ) | ( wire6916 ) ;
 assign wire6919 = ( wire1246 ) | ( wire1248 ) | ( wire6911 ) | ( wire6918 ) ;
 assign wire6923 = ( (~ i_4_)  &  i_12_  &  i_1_ ) ;
 assign wire6924 = ( i_10_  &  i_8_  &  i_12_ ) ;
 assign wire6929 = ( i_9_  &  (~ i_12_)  &  i_11_ ) | ( (~ i_12_)  &  (~ i_1_)  &  i_11_ ) ;
 assign wire6930 = ( i_12_  &  (~ i_1_)  &  (~ i_11_) ) ;
 assign wire6931 = ( (~ i_7_)  &  i_6_  &  wire6929 ) | ( i_7_  &  (~ i_6_)  &  wire6930 ) ;
 assign wire6934 = ( wire1204 ) | ( wire21  &  wire1213 ) | ( wire21  &  wire6931 ) ;
 assign wire6942 = ( (~ i_3_)  &  (~ i_13_)  &  (~ i_12_)  &  i_1_ ) ;
 assign wire6944 = ( i_7_  &  i_1_  &  (~ i_2_) ) ;
 assign wire6952 = ( (~ i_8_)  &  (~ i_4_)  &  (~ i_12_)  &  i_11_ ) ;
 assign wire6958 = ( (~ i_8_)  &  (~ i_13_)  &  i_4_  &  (~ i_2_) ) ;
 assign wire6961 = ( wire25  &  n_n412 ) | ( n_n822  &  wire6958 ) ;
 assign wire6964 = ( n_n792  &  n_n274 ) | ( n_n570  &  n_n240 ) ;
 assign wire6968 = ( (~ i_10_)  &  (~ i_3_)  &  (~ i_13_)  &  i_4_ ) ;
 assign wire6969 = ( n_n849  &  wire351 ) | ( wire352  &  wire6968 ) ;
 assign wire6970 = ( n_n764  &  wire295 ) | ( wire313  &  wire9 ) ;
 assign wire6972 = ( wire1139 ) | ( (~ i_3_)  &  wire616 ) ;
 assign wire6973 = ( wire6970 ) | ( (~ i_7_)  &  wire617 ) ;
 assign wire6982 = ( i_9_  &  i_8_  &  (~ i_2_) ) ;
 assign wire6984 = ( wire1123 ) | ( i_10_  &  (~ i_11_)  &  wire308 ) ;
 assign wire6985 = ( wire1122 ) | ( i_3_  &  i_2_  &  n_n638 ) ;
 assign wire6987 = ( wire6984 ) | ( wire6985 ) | ( i_13_  &  wire626 ) ;
 assign wire6991 = ( n_n1191 ) | ( wire1110 ) | ( (~ i_4_)  &  wire619 ) ;
 assign wire6992 = ( wire1108 ) | ( wire1109 ) | ( wire1121 ) | ( wire6987 ) ;
 assign wire6995 = ( i_8_  &  i_4_  &  (~ i_2_) ) ;
 assign wire6999 = ( n_n1189 ) | ( wire1168 ) | ( wire1169 ) | ( wire6961 ) ;
 assign wire7003 = ( (~ i_7_)  &  i_4_ ) ;
 assign wire7007 = ( n_n835  &  wire293 ) | ( n_n675  &  n_n813 ) ;
 assign wire7008 = ( wire7007 ) | ( n_n792  &  n_n791 ) ;
 assign wire7010 = ( wire41  &  wire382 ) | ( (~ i_2_)  &  wire641 ) ;
 assign wire7011 = ( i_5_  &  (~ i_1_)  &  (~ i_2_) ) ;
 assign wire7021 = ( n_n819  &  n_n678 ) | ( n_n671  &  n_n810 ) ;
 assign wire7022 = ( n_n819  &  n_n712 ) | ( n_n779  &  n_n768 ) ;
 assign wire7023 = ( n_n769  &  n_n771 ) | ( n_n835  &  wire318 ) ;
 assign wire7024 = ( n_n764  &  n_n791 ) | ( wire12  &  wire346 ) ;
 assign wire7027 = ( wire7021 ) | ( wire7024 ) | ( wire322  &  wire330 ) ;
 assign wire7028 = ( wire1047 ) | ( n_n773  &  n_n771 ) ;
 assign wire7029 = ( n_n699  &  n_n710 ) | ( n_n672  &  wire6673 ) ;
 assign wire7030 = ( wire35  &  wire336 ) | ( n_n699  &  n_n678 ) ;
 assign wire7032 = ( wire7030 ) | ( i_4_  &  wire676 ) ;
 assign wire7033 = ( i_5_  &  i_4_  &  (~ i_1_) ) ;
 assign wire7037 = ( n_n683  &  wire351 ) | ( n_n764  &  wire7033 ) ;
 assign wire7040 = ( wire1033 ) | ( wire7028 ) | ( wire7029 ) | ( wire7032 ) ;
 assign wire7041 = ( (~ i_10_)  &  (~ i_2_) ) ;
 assign wire7057 = ( (~ i_5_)  &  (~ i_3_)  &  (~ i_11_)  &  (~ i_2_) ) ;
 assign wire7058 = ( (~ i_9_)  &  i_7_  &  (~ i_12_)  &  (~ i_11_) ) ;
 assign wire7059 = ( n_n773  &  wire7057 ) | ( n_n658  &  wire7058 ) ;
 assign wire7060 = ( wire988 ) | ( n_n701  &  n_n606 ) | ( n_n701  &  wire993 ) ;
 assign wire7062 = ( wire987 ) | ( wire7059 ) | ( wire7060 ) ;
 assign wire7063 = ( wire7010 ) | ( wire7062 ) | ( _430 ) | ( _431 ) ;
 assign wire7070 = ( n_n741  &  wire326 ) | ( n_n792  &  wire7066 ) ;
 assign wire7071 = ( n_n701  &  wire323 ) | ( n_n566  &  wire325 ) ;
 assign wire7074 = ( wire7070 ) | ( wire7071 ) | ( _9382 ) ;
 assign wire7079 = ( (~ i_10_)  &  (~ i_13_)  &  (~ i_11_) ) ;
 assign wire7082 = ( _9672 ) | ( (~ i_13_)  &  (~ i_1_)  &  wire529 ) ;
 assign wire7083 = ( (~ i_5_)  &  (~ i_3_)  &  i_0_ ) ;
 assign wire7092 = ( wire340 ) | ( n_n701  &  _9541 ) ;
 assign wire7104 = ( (~ i_5_)  &  i_6_  &  (~ i_1_) ) ;
 assign wire7105 = ( n_n849  &  n_n813 ) | ( wire294  &  wire7104 ) ;
 assign wire7107 = ( wire7105 ) | ( (~ i_13_)  &  i_11_  &  wire666 ) ;
 assign wire7108 = ( wire70 ) | ( wire917 ) | ( n_n816  &  wire667 ) ;
 assign wire7113 = ( wire907 ) | ( n_n716  &  wire669 ) ;
 assign wire7114 = ( (~ i_5_)  &  (~ i_13_)  &  i_4_  &  i_11_ ) ;
 assign wire7115 = ( n_n816  &  wire671 ) | ( wire336  &  wire7114 ) ;
 assign wire7117 = ( wire7107 ) | ( wire7108 ) | ( _41 ) | ( _42 ) ;
 assign wire7118 = ( wire895 ) | ( wire909 ) | ( wire7113 ) | ( wire7115 ) ;
 assign wire7130 = ( wire26  &  wire638 ) | ( wire284  &  wire637 ) ;
 assign wire7144 = ( (~ i_5_)  &  i_6_  &  i_4_ ) ;
 assign wire7149 = ( wire843 ) | ( wire844 ) | ( wire7138  &  _9611 ) ;
 assign wire7151 = ( wire845 ) | ( wire7130 ) | ( _204 ) ;
 assign wire7163 = ( i_5_  &  (~ i_0_)  &  n_n843 ) ;
 assign wire7164 = ( i_5_  &  (~ i_13_)  &  i_12_  &  (~ i_11_) ) ;
 assign wire7174 = ( i_7_  &  i_5_  &  n_n687 ) ;
 assign wire7177 = ( wire798 ) | ( wire800 ) | ( wire735  &  wire7174 ) ;
 assign wire7182 = ( i_10_  &  i_6_  &  i_12_  &  i_0_ ) ;
 assign wire7183 = ( (~ i_5_)  &  i_6_  &  i_12_  &  (~ i_11_) ) ;
 assign wire7202 = ( i_10_  &  (~ i_8_)  &  (~ i_5_)  &  i_11_ ) ;
 assign wire7211 = ( n_n840  &  wire6803 ) | ( n_n840  &  wire6573 ) ;
 assign wire7214 = ( wire235 ) | ( wire236 ) | ( wire7211 ) ;
 assign wire7218 = ( i_3_  &  (~ i_4_)  &  i_2_  &  i_0_ ) ;
 assign wire7222 = ( wire115 ) | ( wire225 ) | ( wire737  &  wire7218 ) ;
 assign wire7227 = ( i_10_  &  i_12_  &  i_0_ ) ;
 assign wire7228 = ( i_7_  &  i_5_  &  i_0_ ) ;
 assign wire7231 = ( wire212 ) | ( wire213 ) | ( (~ i_4_)  &  wire738 ) ;
 assign wire7237 = ( i_10_  &  (~ i_4_)  &  i_11_ ) ;
 assign wire7241 = ( wire198 ) | ( wire200 ) | ( _284 ) ;
 assign wire7246 = ( (~ i_7_)  &  (~ i_5_)  &  i_2_  &  i_0_ ) ;
 assign wire7248 = ( i_10_  &  (~ i_7_)  &  (~ i_5_)  &  i_11_ ) ;
 assign wire7251 = ( n_n415  &  wire7246 ) | ( n_n598  &  wire7248 ) ;
 assign wire7253 = ( wire190 ) | ( wire7251 ) | ( i_10_  &  wire557 ) ;
 assign wire7254 = ( (~ i_7_)  &  i_6_  &  i_2_ ) ;
 assign wire7260 = ( wire163 ) | ( n_n421  &  n_n598 ) | ( n_n421  &  wire166 ) ;
 assign wire7261 = ( wire283  &  wire565 ) | ( i_2_  &  wire564 ) ;
 assign wire7262 = ( wire7260 ) | ( wire7261 ) ;
 assign wire7263 = ( n_n1000 ) | ( wire192 ) | ( wire7253 ) ;
 assign wire7266 = ( i_5_  &  i_12_  &  i_2_  &  i_0_ ) ;
 assign wire7267 = ( i_8_  &  i_3_  &  i_2_  &  i_0_ ) ;
 assign wire7268 = ( i_9_  &  i_10_  &  i_8_  &  (~ i_5_) ) ;
 assign wire7271 = ( wire397  &  wire7267 ) | ( wire292  &  wire7268 ) ;
 assign wire7272 = ( wire154 ) | ( n_n185  &  wire700 ) ;
 assign wire7273 = ( wire150 ) | ( wire7271 ) | ( wire701  &  wire7266 ) ;
 assign wire7277 = ( wire143 ) | ( wire18  &  wire354  &  wire704 ) ;
 assign wire7278 = ( wire139 ) | ( wire141 ) | ( wire142 ) ;
 assign wire7279 = ( wire7277 ) | ( i_9_  &  i_11_  &  wire703 ) ;
 assign wire7286 = ( i_10_  &  i_3_  &  i_12_  &  i_0_ ) ;
 assign wire7289 = ( n_n421  &  wire123 ) | ( n_n358  &  wire7286 ) ;
 assign wire7292 = ( wire7289 ) | ( (~ i_8_)  &  wire596 ) ;
 assign wire7293 = ( wire127 ) | ( wire128 ) | ( wire129 ) | ( wire130 ) ;
 assign wire7297 = ( n_n453  &  wire308 ) | ( n_n637  &  wire706 ) ;
 assign wire7302 = ( i_7_  &  (~ i_8_)  &  i_6_  &  i_3_ ) ;
 assign wire7303 = ( i_10_  &  (~ i_8_)  &  (~ i_5_)  &  i_12_ ) ;
 assign wire7307 = ( n_n609  &  wire359 ) | ( wire287  &  wire7303 ) ;
 assign wire7308 = ( wire86 ) | ( wire89 ) | ( wire338  &  wire7302 ) ;
 assign wire7309 = ( wire7307 ) | ( _67 ) | ( _68 ) ;
 assign wire7310 = ( wire7292 ) | ( wire7293 ) | ( wire7308 ) ;
 assign wire7311 = ( wire7297 ) | ( wire7309 ) | ( _64 ) | ( _9805 ) ;
 assign wire7314 = ( (~ i_5_)  &  i_1_  &  i_2_  &  i_0_ ) ;
 assign wire7317 = ( wire64 ) | ( wire65 ) | ( wire314  &  wire7314 ) ;
 assign wire7318 = ( wire7317 ) | ( i_9_  &  i_7_  &  wire752 ) ;
 assign wire7319 = ( wire7272 ) | ( wire7273 ) | ( wire7278 ) | ( wire7279 ) ;
 assign wire7321 = ( wire7262 ) | ( wire7263 ) | ( wire7310 ) | ( wire7311 ) ;
 assign wire7324 = ( (~ i_5_)  &  (~ i_6_)  &  (~ i_1_)  &  i_0_ ) ;
 assign wire7326 = ( (~ i_10_)  &  (~ i_7_)  &  (~ i_8_)  &  (~ i_13_) ) ;
 assign wire7335 = ( n_n970 ) | ( n_n957 ) | ( wire961 ) | ( wire7082 ) ;
 assign wire7336 = ( wire7117 ) | ( wire7118 ) | ( _9881 ) ;
 assign _25 = ( (~ i_5_)  &  wire6594  &  wire673  &  _9868 ) ;
 assign _41 = ( (~ i_10_)  &  wire301  &  wire317 ) ;
 assign _42 = ( (~ i_10_)  &  n_n545  &  wire350 ) | ( (~ i_10_)  &  n_n545  &  wire905 ) ;
 assign _52 = ( n_n716  &  n_n675  &  wire7015 ) ;
 assign _53 = ( n_n716  &  n_n503  &  _9846 ) ;
 assign _64 = ( i_10_  &  i_11_  &  wire705 ) ;
 assign _67 = ( (~ i_8_)  &  wire304  &  _9809 ) ;
 assign _68 = ( (~ i_8_)  &  n_n639  &  wire7304  &  _9811 ) ;
 assign _196 = ( (~ i_11_)  &  i_0_  &  n_n575  &  n_n606 ) ;
 assign _197 = ( n_n575  &  n_n670  &  _9640 ) ;
 assign _204 = ( n_n838  &  wire7129 ) | ( n_n838  &  _221 ) | ( n_n838  &  _222 ) ;
 assign _221 = ( i_5_  &  wire319 ) | ( i_5_  &  n_n719  &  _9628 ) ;
 assign _222 = ( i_8_  &  i_5_  &  (~ i_3_)  &  n_n550 ) ;
 assign _267 = ( i_5_  &  i_0_  &  n_n843  &  wire374 ) ;
 assign _268 = ( (~ i_4_)  &  n_n843  &  wire841 ) | ( (~ i_4_)  &  n_n843  &  wire842 ) ;
 assign _274 = ( i_0_  &  _279 ) | ( i_0_  &  n_n741  &  _9543 ) ;
 assign _279 = ( (~ i_13_)  &  n_n566  &  wire19 ) | ( (~ i_13_)  &  n_n566  &  _9544 ) ;
 assign _284 = ( n_n581  &  wire290  &  wire7237 ) | ( wire290  &  wire7237  &  _9532 ) ;
 assign _292 = ( (~ i_4_)  &  i_1_  &  wire7239  &  _9523 ) ;
 assign _296 = ( wire296  &  wire7202 ) ;
 assign _301 = ( i_9_  &  i_11_  &  wire296  &  _9504 ) ;
 assign _310 = ( i_7_  &  wire395  &  _9494 ) ;
 assign _313 = ( (~ i_4_)  &  wire287  &  wire10 ) ;
 assign _314 = ( (~ i_4_)  &  n_n826  &  wire790 ) | ( (~ i_4_)  &  n_n826  &  wire791 ) ;
 assign _319 = ( (~ i_5_)  &  i_3_  &  (~ i_4_)  &  wire736 ) ;
 assign _372 = ( i_3_  &  n_n840  &  wire768 ) | ( i_3_  &  n_n840  &  wire769 ) ;
 assign _411 = ( (~ i_9_)  &  _412 ) | ( (~ i_9_)  &  _413 ) | ( (~ i_9_)  &  _414 ) ;
 assign _412 = ( i_5_  &  (~ i_12_)  &  (~ i_1_)  &  (~ i_11_) ) ;
 assign _413 = ( i_5_  &  i_6_  &  (~ i_12_)  &  (~ i_1_) ) ;
 assign _414 = ( (~ i_10_)  &  (~ i_12_)  &  (~ i_1_)  &  (~ i_11_) ) ;
 assign _430 = ( wire644  &  _9347 ) ;
 assign _431 = ( (~ i_11_)  &  wire1082 ) | ( (~ i_11_)  &  n_n835  &  wire643 ) ;
 assign _459 = ( (~ i_3_)  &  i_4_  &  (~ i_1_)  &  n_n827 ) ;
 assign _520 = ( (~ i_10_)  &  (~ i_12_)  &  wire350 ) | ( (~ i_10_)  &  (~ i_12_)  &  wire1021 ) ;
 assign _523 = ( (~ i_9_)  &  i_7_  &  (~ i_8_)  &  _9277 ) ;
 assign _524 = ( (~ i_11_)  &  n_n503  &  _9279 ) ;
 assign _536 = ( wire14  &  wire104 ) | ( wire14  &  wire1181 ) | ( wire14  &  wire1183 ) ;
 assign _537 = ( (~ i_4_)  &  i_2_  &  wire1180 ) | ( (~ i_4_)  &  i_2_  &  wire1182 ) ;
 assign _575 = ( i_13_  &  (~ i_12_)  &  (~ i_11_)  &  (~ i_2_) ) ;
 assign _629 = ( i_6_  &  n_n716  &  wire1336 ) | ( i_6_  &  n_n716  &  wire1337 ) ;
 assign _630 = ( i_6_  &  n_n764  &  wire371 ) | ( i_6_  &  n_n764  &  wire1334 ) ;
 assign _666 = ( i_6_  &  wire6846  &  _9087 ) ;
 assign _684 = ( (~ i_6_)  &  n_n273  &  wire1202 ) | ( (~ i_6_)  &  n_n273  &  wire1203 ) ;
 assign _685 = ( (~ i_6_)  &  n_n792  &  wire371 ) | ( (~ i_6_)  &  n_n792  &  wire1200 ) ;
 assign _808 = ( wire1414  &  _8904 ) | ( _812  &  _8904 ) | ( _813  &  _8904 ) ;
 assign _810 = ( wire364  &  n_n840  &  wire6573 ) ;
 assign _812 = ( n_n538  &  n_n838  &  n_n832  &  n_n550 ) ;
 assign _813 = ( n_n835  &  n_n541  &  n_n832  &  _8793 ) ;
 assign _840 = ( wire1746  &  _8869 ) | ( _844  &  _8869 ) | ( _845  &  _8869 ) ;
 assign _844 = ( n_n835  &  n_n609 ) | ( n_n609  &  n_n606 ) | ( n_n609  &  wire1750 ) ;
 assign _845 = ( n_n609  &  wire1748 ) | ( n_n609  &  _847 ) ;
 assign _847 = ( (~ i_5_)  &  (~ i_1_)  &  (~ i_2_) ) ;
 assign _855 = ( n_n833  &  n_n541  &  wire423 ) ;
 assign _856 = ( n_n833  &  wire1770 ) | ( n_n833  &  wire424  &  _8833 ) ;
 assign _863 = ( n_n638  &  n_n541  &  wire459 ) ;
 assign _864 = ( n_n638  &  wire1726 ) | ( n_n638  &  wire1729 ) | ( n_n638  &  _865 ) ;
 assign _865 = ( i_5_  &  i_6_  &  (~ i_12_)  &  wire272 ) ;
 assign _870 = ( wire1388  &  _8807 ) | ( _872  &  _8807 ) | ( _873  &  _8807 ) ;
 assign _871 = ( wire1390  &  _8814 ) | ( _880  &  _8814 ) | ( _881  &  _8814 ) ;
 assign _872 = ( n_n637  &  wire123 ) | ( n_n637  &  wire359 ) | ( n_n637  &  wire1397 ) ;
 assign _873 = ( i_13_  &  (~ i_11_)  &  _875 ) | ( i_13_  &  (~ i_11_)  &  _876 ) ;
 assign _875 = ( (~ i_7_)  &  (~ i_5_)  &  (~ i_6_)  &  i_3_ ) ;
 assign _876 = ( (~ i_7_)  &  i_3_  &  i_1_  &  i_0_ ) ;
 assign _880 = ( n_n716  &  n_n847  &  _8808 ) ;
 assign _881 = ( n_n847  &  wire6816  &  _8812 ) ;
 assign _893 = ( n_n538  &  n_n498  &  n_n847  &  n_n843 ) ;
 assign _894 = ( n_n850  &  n_n847  &  n_n541  &  _8768 ) ;
 assign _897 = ( i_13_  &  (~ i_12_)  &  wire314  &  _8758 ) ;
 assign _901 = ( n_n538  &  wire6708  &  _8746  &  _8751 ) ;
 assign _930 = ( i_9_  &  i_10_  &  wire6557  &  wire465 ) ;
 assign _933 = ( n_n665  &  n_n830  &  n_n639  &  n_n597 ) ;
 assign _934 = ( i_13_  &  (~ i_12_)  &  wire6589  &  _8690 ) ;
 assign _941 = ( _948  &  _8681 ) | ( wire468  &  _8678  &  _8681 ) ;
 assign _948 = ( n_n833  &  n_n581  &  _8680 ) ;
 assign _951 = ( n_n665  &  n_n592  &  wire6585 ) | ( n_n665  &  n_n592  &  _8662 ) ;
 assign _952 = ( n_n665  &  n_n597  &  wire6584 ) | ( n_n665  &  n_n597  &  _8664 ) ;
 assign _986 = ( n_n816  &  wire1446  &  _8597 ) | ( n_n816  &  wire1447  &  _8597 ) ;
 assign _987 = ( n_n846  &  n_n822  &  _8598  &  _8600 ) ;
 assign _990 = ( n_n849  &  n_n846  &  wire6771 ) | ( n_n849  &  n_n846  &  wire6772 ) ;
 assign _991 = ( n_n849  &  n_n851  &  wire6770 ) | ( n_n849  &  n_n851  &  _8586 ) ;
 assign _993 = ( (~ i_9_)  &  i_4_  &  wire313 ) ;
 assign _1018 = ( n_n741  &  wire1481  &  _8562 ) ;
 assign _1019 = ( n_n741  &  wire1480  &  _8562 ) ;
 assign _1047 = ( n_n752  &  n_n755  &  n_n840  &  n_n851 ) ;
 assign _1050 = ( n_n853  &  n_n792  &  wire6735 ) | ( n_n853  &  n_n792  &  _8519 ) ;
 assign _1054 = ( (~ i_6_)  &  i_0_  &  n_n795  &  wire369 ) ;
 assign _1081 = ( n_n847  &  n_n832  &  n_n755  &  n_n710 ) ;
 assign _1084 = ( n_n755  &  n_n837  &  n_n840  &  n_n710 ) ;
 assign _1085 = ( n_n838  &  n_n725  &  n_n837  &  n_n735 ) ;
 assign _1113 = ( wire1552  &  _8421 ) | ( wire1553  &  _8421 ) | ( wire1554  &  _8421 ) ;
 assign _1114 = ( _1122  &  _8427 ) | ( wire551  &  _8424  &  _8427 ) ;
 assign _1122 = ( (~ i_3_)  &  n_n746  &  n_n840  &  _8425 ) ;
 assign _8162 = ( i_8_  &  (~ i_13_)  &  i_12_ ) ;
 assign _8227 = ( i_8_  &  i_12_  &  i_11_ ) ;
 assign _8232 = ( wire292 ) | ( wire1798 ) | ( wire6509  &  _8227 ) ;
 assign _8334 = ( (~ i_1_)  &  i_2_  &  (~ i_0_) ) ;
 assign _8369 = ( (~ i_9_)  &  i_5_  &  i_6_ ) ;
 assign _8395 = ( (~ i_9_)  &  i_7_  &  i_5_ ) ;
 assign _8407 = ( wire6678 ) | ( n_n853  &  wire6674 ) | ( n_n853  &  wire6675 ) ;
 assign _8421 = ( (~ i_12_)  &  i_13_ ) ;
 assign _8424 = ( i_10_  &  i_7_  &  i_8_  &  (~ i_3_) ) ;
 assign _8425 = ( i_5_  &  i_10_ ) ;
 assign _8427 = ( (~ i_12_)  &  i_13_ ) ;
 assign _8446 = ( (~ i_9_)  &  (~ i_13_)  &  i_12_  &  (~ i_11_) ) ;
 assign _8451 = ( (~ i_13_)  &  i_12_  &  i_0_ ) ;
 assign _8457 = ( (~ i_10_)  &  (~ i_13_)  &  (~ i_11_) ) ;
 assign _8480 = ( (~ i_9_)  &  (~ i_13_)  &  i_11_ ) ;
 assign _8482 = ( (~ i_1_)  &  (~ i_2_)  &  i_0_ ) ;
 assign _8489 = ( (~ i_9_)  &  (~ i_13_)  &  i_11_ ) ;
 assign _8492 = ( (~ i_10_)  &  (~ i_13_)  &  i_12_ ) ;
 assign _8496 = ( (~ i_9_)  &  (~ i_3_)  &  (~ i_13_)  &  (~ i_4_) ) ;
 assign _8509 = ( (~ i_9_)  &  (~ i_7_)  &  (~ i_8_)  &  i_4_ ) ;
 assign _8519 = ( (~ i_5_)  &  i_4_  &  (~ i_1_) ) ;
 assign _8521 = ( wire69 ) | ( wire70 ) | ( wire106 ) | ( _1050 ) ;
 assign _8562 = ( (~ i_13_)  &  (~ i_4_)  &  i_12_  &  i_2_ ) ;
 assign _8586 = ( i_7_  &  (~ i_8_)  &  (~ i_6_)  &  n_n833 ) ;
 assign _8588 = ( (~ i_9_)  &  (~ i_7_)  &  (~ i_13_)  &  i_1_ ) ;
 assign _8597 = ( (~ i_6_)  &  (~ i_7_) ) ;
 assign _8598 = ( (~ i_13_)  &  (~ i_9_) ) ;
 assign _8600 = ( (~ i_6_)  &  (~ i_7_) ) ;
 assign _8610 = ( wire1436 ) | ( wire1437 ) | ( _986 ) | ( _987 ) ;
 assign _8633 = ( (~ i_10_)  &  (~ i_8_)  &  i_12_  &  i_11_ ) ;
 assign _8662 = ( (~ i_1_)  &  i_2_  &  (~ i_0_)  &  n_n633 ) ;
 assign _8664 = ( (~ i_5_)  &  (~ i_6_)  &  i_3_  &  n_n833 ) ;
 assign _8678 = ( i_9_  &  (~ i_7_)  &  (~ i_8_)  &  (~ i_3_) ) ;
 assign _8680 = ( i_5_  &  i_6_  &  (~ i_3_) ) ;
 assign _8681 = ( (~ i_11_)  &  i_13_ ) ;
 assign _8690 = ( i_10_  &  (~ i_8_)  &  (~ i_11_) ) ;
 assign _8728 = ( i_8_  &  (~ i_3_)  &  (~ i_13_) ) ;
 assign _8746 = ( (~ i_1_)  &  i_2_  &  i_0_ ) ;
 assign _8747 = ( i_10_  &  (~ i_11_)  &  n_n538  &  _8746 ) ;
 assign _8751 = ( (~ i_9_)  &  (~ i_13_)  &  (~ i_12_) ) ;
 assign _8758 = ( i_5_  &  i_6_  &  i_3_ ) ;
 assign _8768 = ( i_10_  &  (~ i_13_)  &  (~ i_12_)  &  i_11_ ) ;
 assign _8774 = ( n_n1243 ) | ( wire1686 ) | ( wire6605 ) ;
 assign _8793 = ( (~ i_12_)  &  (~ i_13_) ) ;
 assign _8807 = ( i_10_  &  i_9_ ) ;
 assign _8808 = ( i_5_  &  (~ i_6_)  &  i_3_  &  (~ i_4_) ) ;
 assign _8812 = ( (~ i_5_)  &  i_3_  &  (~ i_4_) ) ;
 assign _8814 = ( i_10_  &  i_9_ ) ;
 assign _8824 = ( i_6_  &  i_1_  &  i_2_  &  (~ i_0_) ) ;
 assign _8833 = ( i_10_  &  (~ i_11_)  &  n_n538 ) ;
 assign _8842 = ( wire1764 ) | ( wire1763 ) ;
 assign _8852 = ( wire1720 ) | ( n_n844  &  n_n752  &  wire307 ) ;
 assign _8853 = ( wire1722 ) | ( wire1765 ) | ( _8842 ) | ( _8852 ) ;
 assign _8854 = ( _855 ) | ( _856 ) | ( _863 ) | ( _864 ) ;
 assign _8869 = ( (~ i_12_)  &  i_13_ ) ;
 assign _8904 = ( i_11_  &  i_10_ ) ;
 assign _8905 = ( wire1744 ) | ( _840 ) | ( i_10_  &  wire583 ) ;
 assign _8908 = ( n_n1234 ) | ( wire1385 ) | ( _8853 ) | ( _8854 ) ;
 assign _8989 = ( i_6_  &  wire1274 ) | ( i_6_  &  wire6893 ) ;
 assign _9006 = ( (~ i_6_)  &  wire1263 ) | ( (~ i_6_)  &  wire6902 ) ;
 assign _9028 = ( i_9_  &  i_8_  &  (~ i_12_)  &  (~ i_11_) ) ;
 assign _9029 = ( i_9_  &  i_8_  &  (~ i_6_)  &  (~ i_11_) ) ;
 assign _9050 = ( wire6896 ) | ( wire6905 ) | ( _8989 ) | ( _9006 ) ;
 assign _9055 = ( (~ i_6_)  &  (~ i_13_)  &  i_1_  &  (~ i_2_) ) ;
 assign _9087 = ( (~ i_9_)  &  i_7_  &  (~ i_8_) ) ;
 assign _9093 = ( (~ i_9_)  &  i_7_  &  i_6_  &  i_1_ ) ;
 assign _9115 = ( (~ i_6_)  &  (~ i_3_)  &  (~ i_1_)  &  (~ i_2_) ) ;
 assign _9128 = ( i_6_  &  (~ i_13_)  &  i_12_ ) ;
 assign _9139 = ( (~ i_9_)  &  (~ i_10_)  &  i_8_  &  (~ i_3_) ) ;
 assign _9141 = ( wire301  &  wire6864 ) | ( wire346  &  _9128 ) ;
 assign _9151 = ( i_7_  &  (~ i_13_)  &  i_1_  &  (~ i_2_) ) ;
 assign _9152 = ( n_n849  &  n_n810 ) | ( n_n566  &  _9151 ) ;
 assign _9168 = ( wire1340 ) | ( _629 ) | ( _630 ) | ( _9152 ) ;
 assign _9176 = ( (~ i_10_)  &  (~ i_13_)  &  i_11_ ) ;
 assign _9183 = ( (~ i_8_)  &  (~ i_3_)  &  (~ i_13_) ) ;
 assign _9185 = ( (~ i_9_)  &  (~ i_3_)  &  (~ i_13_) ) ;
 assign _9186 = ( wire340 ) | ( n_n741  &  _9183 ) ;
 assign _9187 = ( wire1154 ) | ( i_2_  &  wire1166 ) | ( i_2_  &  _9186 ) ;
 assign _9198 = ( (~ i_7_)  &  i_8_  &  (~ i_3_) ) ;
 assign _9200 = ( i_7_  &  (~ i_13_)  &  i_12_ ) ;
 assign _9211 = ( i_3_  &  (~ i_12_)  &  (~ i_2_) ) ;
 assign _9277 = ( i_5_  &  i_6_  &  (~ i_3_)  &  (~ i_11_) ) ;
 assign _9279 = ( i_5_  &  (~ i_3_)  &  (~ i_2_) ) ;
 assign _9280 = ( (~ i_12_)  &  (~ i_1_)  &  (~ i_2_) ) ;
 assign _9285 = ( (~ i_3_)  &  (~ i_8_) ) ;
 assign _9288 = ( wire7046 ) | ( wire7047 ) | ( _523 ) | ( _524 ) ;
 assign _9290 = ( (~ i_10_)  &  i_8_  &  (~ i_5_) ) ;
 assign _9296 = ( (~ i_2_)  &  i_7_ ) ;
 assign _9297 = ( wire1023 ) | ( n_n566  &  wire19 ) | ( n_n566  &  _9296 ) ;
 assign _9303 = ( (~ i_10_)  &  i_8_  &  (~ i_6_) ) ;
 assign _9304 = ( (~ i_3_)  &  i_8_ ) ;
 assign _9309 = ( wire1012 ) | ( wire1024 ) | ( _9288 ) | ( _9297 ) ;
 assign _9324 = ( wire7019 ) | ( wire382  &  wire324 ) ;
 assign _9328 = ( wire7022 ) | ( wire7023 ) | ( wire7037 ) | ( _459 ) ;
 assign _9347 = ( (~ i_3_)  &  (~ i_11_)  &  (~ i_2_)  &  (~ i_0_) ) ;
 assign _9362 = ( wire1064 ) | ( wire7027 ) | ( _9324 ) | ( _9328 ) ;
 assign _9364 = ( (~ i_9_)  &  (~ i_12_)  &  (~ i_11_) ) ;
 assign _9376 = ( (~ i_10_)  &  (~ i_8_)  &  (~ i_5_)  &  (~ i_11_) ) ;
 assign _9380 = ( (~ i_9_)  &  i_7_  &  i_8_ ) ;
 assign _9382 = ( n_n675  &  _9376 ) | ( wire7068  &  _9380 ) ;
 assign _9386 = ( wire7076 ) | ( _9309 ) | ( (~ i_12_)  &  wire696 ) ;
 assign _9409 = ( i_7_  &  i_8_  &  i_6_  &  i_3_ ) ;
 assign _9492 = ( i_7_  &  i_12_  &  (~ i_11_) ) ;
 assign _9494 = ( i_3_  &  (~ i_4_)  &  i_0_ ) ;
 assign _9496 = ( _313 ) | ( _314 ) | ( wire354  &  wire708 ) ;
 assign _9504 = ( i_5_  &  (~ i_8_) ) ;
 assign _9512 = ( wire246 ) | ( wire247 ) | ( wire245 ) | ( _296 ) ;
 assign _9523 = ( i_9_  &  (~ i_7_)  &  (~ i_8_) ) ;
 assign _9528 = ( (~ i_8_)  &  (~ i_4_)  &  i_2_  &  (~ i_0_) ) ;
 assign _9529 = ( i_9_  &  (~ i_8_)  &  (~ i_4_)  &  i_2_ ) ;
 assign _9532 = ( (~ i_8_)  &  (~ i_5_)  &  i_2_ ) ;
 assign _9535 = ( wire249 ) | ( wire201 ) | ( _9512 ) ;
 assign _9536 = ( wire785 ) | ( wire7241 ) | ( _9496 ) ;
 assign _9537 = ( wire7232 ) | ( wire215 ) | ( wire7222 ) | ( _319 ) ;
 assign _9539 = ( i_5_  &  (~ i_13_)  &  i_12_ ) ;
 assign _9541 = ( (~ i_9_)  &  (~ i_13_)  &  (~ i_2_) ) ;
 assign _9542 = ( n_n741  &  _9183 ) | ( n_n701  &  _9185 ) ;
 assign _9543 = ( (~ i_7_)  &  (~ i_13_)  &  (~ i_2_) ) ;
 assign _9544 = ( (~ i_2_)  &  i_7_ ) ;
 assign _9545 = ( wire937 ) | ( i_0_  &  wire7092 ) | ( i_0_  &  _9542 ) ;
 assign _9570 = ( wire7168 ) | ( wire7167 ) ;
 assign _9589 = ( wire801 ) | ( wire7177 ) | ( _274 ) | ( _9545 ) ;
 assign _9611 = ( i_7_  &  (~ i_13_)  &  (~ i_12_)  &  i_11_ ) ;
 assign _9615 = ( i_7_  &  i_8_  &  (~ i_5_) ) ;
 assign _9628 = ( (~ i_3_)  &  (~ i_8_) ) ;
 assign _9640 = ( i_8_  &  (~ i_5_)  &  (~ i_6_) ) ;
 assign _9669 = ( (~ i_9_)  &  (~ i_13_)  &  (~ i_1_)  &  i_0_ ) ;
 assign _9672 = ( wire350  &  wire7078 ) | ( n_n701  &  _9669 ) ;
 assign _9676 = ( n_n981 ) | ( wire7149 ) | ( wire7151 ) ;
 assign _9805 = ( wire103 ) | ( wire107 ) | ( wire112 ) ;
 assign _9809 = ( i_3_  &  i_2_  &  i_0_ ) ;
 assign _9811 = ( i_2_  &  (~ i_12_) ) ;
 assign _9837 = ( wire925 ) | ( i_5_  &  i_0_  &  wire578 ) ;
 assign _9846 = ( i_5_  &  (~ i_3_)  &  (~ i_2_) ) ;
 assign _9853 = ( i_4_  &  (~ i_1_)  &  (~ i_2_) ) ;
 assign _9856 = ( wire881 ) | ( wire882 ) | ( _52 ) | ( _53 ) ;
 assign _9867 = ( (~ i_9_)  &  (~ i_5_)  &  i_4_ ) ;
 assign _9868 = ( (~ i_10_)  &  (~ i_9_) ) ;
 assign _9881 = ( wire7102 ) | ( wire884 ) | ( _9837 ) | ( _9856 ) ;
 assign _9885 = ( wire7337 ) | ( wire7335 ) | ( _9676 ) ;


endmodule

