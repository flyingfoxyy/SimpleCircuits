module apex4_2 (
	i_7_, i_8_, i_5_, i_6_, i_3_, i_4_, i_1_, i_2_, 
	i_0_, o_1_, o_2_, o_0_, o_12_, o_11_, o_14_, o_13_, o_16_, o_15_, 
	o_18_, o_17_, o_10_, o_9_, o_7_, o_8_, o_5_, o_6_, o_3_, o_4_);

input i_7_, i_8_, i_5_, i_6_, i_3_, i_4_, i_1_, i_2_, i_0_;

output o_1_, o_2_, o_0_, o_12_, o_11_, o_14_, o_13_, o_16_, o_15_, o_18_, o_17_, o_10_, o_9_, o_7_, o_8_, o_5_, o_6_, o_3_, o_4_;

wire n_n105, n_n127, n_n720, n_n842, wire4717, wire4735, n_n889, wire4767, n_n912, n_n580, n_n445, n_n513, n_n303, n_n372, n_n192, n_n244, n_n1324, n_n94, n_n1176, n_n78, n_n1254, n_n93, n_n1132, n_n92, n_n1259, wire4614, n_n856, n_n855, n_n846, n_n999, n_n97, n_n1004, n_n95, n_n995, n_n63, n_n77, n_n101, n_n1216, n_n975, n_n987, n_n504, n_n964, n_n814, n_n809, n_n804, n_n1060, n_n83, n_n58, n_n1055, n_n82, n_n1160, n_n1181, n_n771, n_n874, n_n1092, n_n730, n_n726, wire4608, n_n81, n_n1009, n_n1011, n_n1087, n_n1082, n_n1217, n_n84, n_n951, n_n956, n_n943, n_n676, n_n665, n_n658, n_n661, wire4879, n_n90, n_n967, n_n957, n_n602, n_n591, n_n601, n_n584, wire4935, n_n990, n_n991, n_n986, n_n102, n_n1100, n_n1095, n_n1184, n_n96, n_n1283, n_n1058, wire5164, n_n530, n_n529, n_n531, n_n71, n_n968, n_n969, n_n1045, n_n1046, n_n1043, wire5034, n_n80, n_n953, n_n954, n_n952, n_n54, n_n1006, n_n1074, n_n91, n_n1077, n_n1068, n_n1169, n_n1088, wire5324, n_n1047, n_n1042, n_n87, n_n1147, n_n994, n_n322, n_n311, n_n958, n_n962, n_n1048, n_n1164, n_n1105, n_n257, wire5389, wire5393, n_n252, n_n254, n_n246, n_n66, n_n974, n_n980, n_n67, n_n1146, n_n1145, n_n40, n_n1122, wire5337, n_n205, n_n195, n_n202, n_n208, n_n196, n_n1022, n_n1204, wire4411, n_n144, n_n131, n_n141, n_n147, wire4354, n_n106, n_n99, n_n100, n_n939, n_n85, n_n79, n_n86, n_n76, n_n75, n_n960, n_n74, n_n103, n_n973, n_n981, n_n989, n_n1134, n_n1163, n_n1172, n_n64, n_n937, wire4762, n_n918, n_n1109, n_n1032, wire4743, n_n890, n_n892, n_n853, n_n852, n_n854, n_n950, n_n955, n_n940, n_n815, n_n941, n_n1040, n_n1039, n_n1128, wire4462, n_n1085, n_n1091, n_n1078, n_n1153, n_n1170, n_n554, wire4570, n_n732, n_n727, n_n722, n_n735, n_n1018, n_n1081, n_n664, n_n662, n_n666, n_n652, n_n590, n_n588, n_n587, wire4956, n_n1001, n_n993, n_n1079, n_n1193, n_n1188, n_n1279, wire5168, n_n527, n_n533, n_n532, n_n518, n_n971, n_n1035, wire5060, n_n466, n_n465, n_n654, n_n451, n_n947, n_n944, n_n1013, n_n1010, n_n421, n_n1177, n_n390, n_n389, wire5268, n_n1144, n_n977, n_n983, n_n970, n_n365, n_n1331, n_n310, n_n942, n_n1057, n_n1156, wire5415, n_n256, wire5420, n_n984, wire5341, n_n204, n_n198, n_n1330, n_n137, n_n134, n_n133, n_n135, n_n128, wire4164, n_n70, n_n982, n_n52, n_n73, n_n1173, n_n946, n_n1125, wire4670, n_n966, n_n1070, n_n812, wire4681, n_n811, wire4685, n_n1036, n_n1075, n_n1185, n_n728, n_n949, wire4873, wire4813, n_n670, n_n1267, wire5003, n_n978, n_n53, n_n1158, wire5176, n_n526, wire5108, n_n523, n_n525, n_n959, wire5010, wire5056, wire5102, n_n1014, n_n1294, n_n1028, n_n1130, n_n320, n_n1215, wire5192, wire5216, n_n309, wire5255, n_n1030, n_n259, n_n258, n_n295, n_n248, n_n1019, n_n1020, n_n136, n_n1281, wire4181, n_n1093, n_n1103, n_n1297, n_n1286, n_n1369, wire4715, wire4690, n_n808, wire4694, n_n1021, n_n1054, n_n961, n_n716, wire4877, n_n663, n_n582, n_n595, n_n1025, n_n1026, wire5017, n_n453, n_n455, n_n446, n_n458, n_n1120, n_n1117, n_n1002, n_n321, wire5198, n_n312, n_n206, n_n1174, n_n109, n_n775, n_n773, n_n770, n_n765, n_n774, wire4524, n_n1052, n_n669, n_n598, n_n521, wire5042, wire5048, n_n456, wire5054, n_n976, n_n1121, wire5203, n_n315, n_n308, n_n319, n_n325, wire5444, wire5365, n_n882, n_n145, wire4211, n_n110, n_n1108, n_n1118, n_n849, n_n776, n_n668, n_n641, n_n599, wire5130, wire5208, n_n314, n_n250, n_n146, n_n850, n_n734, n_n733, n_n671, n_n672, wire4836, n_n1101, n_n600, wire4985, wire4977, n_n1312, n_n519, n_n520, wire5136, n_n463, wire5079, n_n464, n_n324, wire5234, wire5214, n_n140, wire4662, n_n769, n_n768, wire4556, n_n594, wire5178, n_n460, wire5092, n_n459, wire5100, n_n318, wire5242, wire5405, wire4296, n_n1059, n_n395, wire5294, n_n384, n_n392, n_n378, n_n379, wire5290, wire5437, n_n262, n_n261, n_n904, wire5301, n_n385, n_n374, n_n386, wire5333, wire5375, n_n199, n_n142, n_n393, n_n382, wire5306, n_n143, wire5315, wire4664, wire5350, n_n201, wire4934, n_n388, wire5331, wire4909, n_n596, wire4914, _19, _20, _21, _22, _23, _24, _25, _26, _27, _28, _29, _30, _31, _32, _33, _34, _35, _36, _37, _38, _39, _40, _41, _42, _43, _44, _45, _46, _47, _48, _49, _50, _51, _52, _53, _54, _55, _56, _57, _58, _59, _60, _61, _62, _63, _64, _65, _66, _67, _68, _69, _70, _71, _72, _73, _74, _75, _76, _77, _78, _79, _80, _81, _82, _83, _84, _85, _86, _87, _88, _89, _90, _91, _92, _93, _94, _95, _96, _97, _98, _99, _100, _102, _103, _104, _107, _108, _109, _110, _111, _112, _113, _114, _115, _116, _117, _119, _121, _122, _123, _124, _125, _126, _127, _128, _129, _130, _131, _132, _133, _134, _135, _136, _137, _138, _140, _142, _143, _144, _145, _147, _148, _149, _150, _151, _152, _153, _154, _155, _156, _157, _158, _159, _160, _161, _162, _163, _164, _165, _166, _167, _168, _169, _170, _171, _172, _173, _174, _176, _177, _178, _180, _181, _182, _183, _184, _185, _186, _187, _188, _189, _190, _191, _192, _193, _194, _195, _196, _197, _198, _199, _200, _201, _202, _203, _204, _205, _206, _207, _208, _209, _210, _211, _212, _213, _214, _215, _216, _217, _218, _219, _220, _221, _222, _223, _224, _226, _227, _228, _230, _231, _232, _233, _235, _236, _237, _238, _239, _240, _243, _244, _245, _246, _248, _249, _250, _252, _254, _255, _257, _259, _260, _261, _262, _263, _264, _265, _267, _268, _269, _270, _271, _272, _273, _274, _275, _276, _277, _278, _279, _282, _283, _284, _286, _287, _288, _289, _290, _291, _293, _295, _296, _297, _298, _299, _300, _301, _302, _303, _304, _305, _306, _307, _308, _309, _310, _311, _312, _313, _314, _315, _316, _317, _318, _319, _320, _321, _322, _323, _324, _325, _326, _327, _328, _329, _330, _331, _332, _333, _334, _335, _336, _337, _338, _339, _340, _341, _342, _343, _344, _345, _346, _347, _348, _349, _350, _351, _352, _353, _354, _355, _356, _357, _358, _359, _360, _361, _362, _363, _364, _365, _366, _367, _368, _369, _370, _371, _372, _373, _374, _381, _382, _387, _388, _389, _392, _398, _399, _404, _410, _411, _416, _422, _423, _424, _430, _431, _437, _445, _447, _453, _454, _461, _468, _475, _476, _481, _482, _489, _497, _501, _502, _507, _513, _520, _522, _524, _531, _537, _538, _543, _549, _556, _557, _561, _567, _568, _569, _573, _574, _581, _583, _590, _596, _604, _610, _611, _616, _617, _624, _632, _634, _635, _636, _640, _646, _652, _658, _659, _660, _664, _671, _675, _676, _681, _687, _693, _696, _702, _709, _710, _717, _722, _723, _724, _732, _734, _740, _741, _747, _748, _749, _753, _758, _759, _765, _766, _767, _768, _769, _771, _778, _780, _786, _792, _794, _795, _796, _797, _798, _799, _800, _804, _812, _818, _825, _827, _833, _834, _839, _841, _848, _850, _852, _854, _856, _864, _865, _870, _876, _878, _884, _885, _892, _899, _901, _903, _911, _913, _915, _917, _923, _925, _927, _935, _943, _951, _952, _953, _958, _959, _960, _968, _969, _970, _971, _972, _973, _978, _986, _987, _988, _990, _991, _996, _1004, _1010, _1017, _1018, _1019, _1021, _1023, _1030, _1032, _1034, _1035, _1036, _1037, _1041, _1042, _1046, _1047, _1048, _1049, _1052, _1053, _1054, _1056, _1057, _4385, _4386, _4387, _4388, _4389, _4390, _4391, _4392, _4393, _4394, _4395, _4396, _4397, _4398, _4399, _4400, _4401, _4402, _4403, _4404, _4405, _4406, _4407, _4408, _4409, _4410, _4411, _4412, _4413, _4414, _4415, _4416, _4417, _4418, _4419, _4420, _4421, _4422, _4423, _4424, _4425, _4426, _4427, _4428, _4429, _4430, _4431, _4432, _4433, _4434, _4435, _4436, _4437, _4438, _4439, _4440, _4441, _4442, _4443, _4444, _4445, _4446, _4447, _4448, _4449, _4450, _4451, _4452, _4453, _4454, _4455, _4456, _4457, _4458, _4459, _4460, _4461, _4462, _4463, _4464, _4465, _4466, _4467, _4468, _4469, _4470, _4471, _4472, _4473, _4474, _4475, _4476, _4477, _4478, _4479, _4480, _4481, _4482, _4483, _4484, _4485, _4486, _4487, _4488, _4489, _4490, _4491, _4492, _4493, _4494, _4495, _4496, _4497, _4498, _4499, _4500, _4501, _4502, _4503, _4504, _4505, _4506, _4507, _4508, _4509, _4510, _4511, _4512, _4513, _4514, _4515, _4516, _4517, _4518, _4519, _4520, _4521, _4522, _4523, _4524, _4525, _4526, _4527, _4528, _4529, _4530, _4531, _4532, _4533, _4534, _4535, _4536, _4537, _4538, _4539, _4540, _4541, _4542, _4543, _4544, _4545, _4546, _4547, _4548, _4549, _4550, _4551, _4552, _4553, _4554, _4555, _4556, _4557, _4558, _4559, _4560, _4561, _4562, _4563, _4564, _4565, _4566, _4567, _4568, _4569, _4570, _4571, _4572, _4573, _4574, _4575, _4576, _4577, _4578, _4579, _4580, _4581, _4582, _4583, _4584, _4585, _4586, _4587, _4588, _4589, _4590, _4591, _4592, _4593, _4594, _4595, _4596, _4597, _4598, _4599, _4600, _4601, _4602, _4603, _4604, _4605, _4606, _4607, _4608, _4609, _4610, _4611, _4612, _4613, _4614, _4615, _4616, _4617, _4618, _4619, _4620, _4621, _4622, _4623, _4624, _4625, _4626, _4627, _4628, _4629, _4630, _4631, _4632, _4633, _4634, _4635, _4636, _4637, _4638, _4639, _4640, _4641, _4642, _4643, _4644, _4645, _4646, _4647, _4648, _4649, _4650, _4651, _4652, _4653, _4654, _4655, _4656, _4657, _4658, _4659, _4660, _4661, _4662, _4663, _4664, _4665, _4666, _4667, _4668, _4669, _4670, _4671, _4672, _4673, _4674, _4675, _4676, _4677, _4678, _4679, _4680, _4681, _4682, _4683, _4684, _4685, _4686, _4687, _4688, _4689, _4690, _4691, _4692, _4693, _4694, _4695, _4696, _4697, _4698, _4699, _4700, _4701, _4702, _4703, _4704, _4705, _4706, _4707, _4708, _4709, _4710, _4711, _4712, _4713, _4714, _4715, _4716, _4717, _4718, _4719, _4720, _4721, _4722, _4723, _4724, _4725, _4726, _4727, _4728, _4729, _4730, _4731, _4732, _4733, _4734, _4735, _4736, _4737, _4738, _4739, _4740, _4741, _4742, _4743, _4744, _4745, _4746, _4747, _4748, _4749, _4750, _4751, _4752, _4753, _4754, _4755, _4756, _4757, _4758, _4759, _4760, _4761, _4762, _4763, _4764, _4765, _4766, _4767, _4768, _4769, _4770, _4771, _4772, _4773, _4774, _4775, _4776, _4777, _4778, _4779, _4780, _4781, _4782, _4783, _4784, _4785, _4786, _4787, _4788, _4789, _4790, _4791, _4792, _4793, _4794, _4795, _4796, _4797, _4798, _4799, _4800, _4801, _4802, _4803, _4804, _4805, _4806, _4807, _4808, _4809, _4810, _4811, _4812, _4813, _4814, _4815, _4816, _4817, _4818, _4819, _4820, _4821, _4822, _4823, _4824, _4825, _4826, _4827, _4828, _4829, _4830, _4831, _4832, _4833, _4834, _4835, _4836, _4837, _4838, _4839, _4840, _4841, _4842, _4843, _4844, _4845, _4846, _4847, _4848, _4849, _4850, _4851, _4852, _4853, _4854, _4855, _4856, _4857, _4858, _4859, _4860, _4861, _4862, _4863, _4864, _4865, _4866, _4867, _4868, _4869, _4870, _4871, _4872, _4873, _4874, _4875, _4876, _4877, _4878, _4879, _4880, _4881, _4882, _4883, _4884, _4885, _4886, _4887, _4888, _4889, _4890, _4891, _4892, _4893, _4894, _4895, _4896, _4897, _4898, _4899, _4900, _4901, _4902, _4903, _4904, _4905, _4906, _4907, _4908, _4909, _4910, _4911, _4912, _4913, _4914, _4915, _4916, _4917, _4918, _4919, _4920, _4921, _4922, _4923, _4924, _4925, _4926, _4927, _4928, _4929, _4930, _4931, _4932, _4933, _4934, _4935, _4936, _4937, _4938, _4939, _4940, _4941, _4942, _4943, _4944, _4945, _4946, _4947, _4948, _4949, _4950, _4951, _4952, _4953, _4954, _4955, _4956, _4957, _4958, _4959, _4960, _4961, _4962, _4963, _4964, _4965, _4966, _4967, _4968, _4969, _4970, _4971, _4972, _4973, _4974, _4975, _4976, _4977, _4978, _4979, _4980, _4981, _4982, _4983, _4984, _4985, _4986, _4987, _4988, _4989, _4990, _4991, _4992, _4993, _4994, _4995, _4996, _4997, _4998, _4999, _5000, _5001, _5002, _5003, _5004, _5005, _5006, _5007, _5008, _5009, _5010, _5011, _5012, _5013, _5014, _5015, _5016, _5017, _5018, _5019, _5020, _5021, _5022, _5023, _5024, _5025, _5026, _5027, _5028, _5029, _5030, _5031, _5032, _5033, _5034, _5035, _5036, _5037, _5038, _5039, _5040, _5041, _5042, _5043, _5044, _5045, _5046, _5047, _5048, _5049, _5050, _5051, _5052, _5053, _5054, _5055, _5056, _5057, _5058, _5059, _5060, _5061, _5062, _5063, _5064, _5065, _5066, _5067, _5068, _5069, _5070, _5071, _5072, _5073, _5074, _5075, _5076, _5077, _5078, _5079, _5080, _5081, _5082, _5083, _5084, _5085, _5086, _5087, _5088, _5089, _5090, _5091, _5092, _5093, _5094, _5095, _5096, _5097, _5098, _5099, _5100, _5101, _5102, _5103, _5104, _5105, _5106, _5107, _5108, _5109, _5110, _5111, _5112, _5113, _5114, _5115, _5116, _5117, _5118, _5119, _5120, _5121, _5122, _5123, _5124, _5125, _5126, _5127, _5128, _5129, _5130, _5131, _5132, _5133, _5134, _5135, _5136, _5137, _5138, _5139, _5140, _5141, _5142, _5143, _5144, _5145, _5146, _5147, _5148, _5149, _5150, _5151, _5152, _5153, _5154, _5155, _5156, _5157, _5158, _5159, _5160, _5161, _5162, _5163, _5164, _5165, _5166, _5167, _5168, _5169, _5170, _5171, _5172, _5173, _5174, _5175, _5176, _5177, _5178, _5179, _5180, _5181, _5182, _5183, _5184, _5185, _5186, _5187, _5188, _5189, _5190, _5191, _5192, _5193, _5194, _5195, _5196, _5197, _5198, _5199, _5200, _5201, _5202, _5203, _5204, _5205, _5206, _5207, _5208, _5209, _5210, _5211, _5212, _5213, _5214, _5215, _5216, _5217, _5218, _5219, _5220, _5221, _5222, _5223, _5224, _5225, _5226, _5227, _5228, _5229, _5230, _5231, _5232, _5233, _5234, _5235, _5236, _5237, _5238, _5239, _5240, _5241, _5242, _5243, _5244, _5245, _5246, _5247, _5248, _5249, _5250, _5251, _5252, _5253, _5254, _5255, _5256, _5257, _5258, _5259, _5260, _5261, _5262, _5263, _5264, _5265, _5266, _5267, _5268, _5269, _5270, _5271, _5272, _5273, _5274, _5275, _5276, _5277, _5278, _5279, _5280, _5281, _5282, _5283, _5284, _5285, _5286, _5287, _5288, _5289, _5290, _5291, _5292, _5293, _5294, _5295, _5296, _5297, _5298, _5299, _5300, _5301, _5302, _5303, _5304, _5305, _5306, _5307, _5308, _5309, _5310, _5311, _5312, _5313, _5314, _5315, _5316, _5317, _5318, _5319, _5320, _5321, _5322, _5323, _5324, _5325, _5326, _5327, _5328, _5329, _5330, _5331, _5332, _5333, _5334, _5335, _5336, _5337, _5338, _5339, _5340, _5341, _5342, _5343, _5344, _5345, _5346, _5347, _5348, _5349, _5350, _5351, _5352, _5353, _5354, _5355, _5356, _5357, _5358, _5359, _5360, _5361, _5362, _5363, _5364, _5365, _5366, _5367, _5368, _5369, _5370, _5371, _5372, _5373, _5374, _5375, _5376, _5377, _5378, _5379, _5380, _5381, _5382, _5383, _5384, _5385, _5386, _5387, _5388, _5389, _5390, _5391, _5392, _5393, _5394, _5395, _5396, _5397, _5398, _5399, _5400, _5401, _5402, _5403, _5404, _5405, _5406, _5407, _5408, _5409, _5410, _5411, _5412, _5413, _5414, _5415, _5416, _5417, _5418, _5419, _5420, _5421, _5422, _5423, _5424, _5425, _5426, _5427, _5428, _5429, _5430, _5431, _5432, _5433, _5434, _5435, _5436, _5437, _5438, _5439, _5440, _5441, _5442, _5443, _5444, _5445, _5446, _5447, _5448, _5449, _5450, _5451, _5452, _5453, _5454, _5455, _5456, _5457, _5458, _5459, _5460, _5461, _5462, _5463, _5464, _5465, _5466, _5467, _5468, _5469, _5470, _5471, _5472, _5473, _5474, _5475, _5476, _5477, _5478, _5479, _5480, _5481, _5482, _5483, _5484, _5485, _5486, _5487, _5488, _5489, _5490, _5491, _5492, _5493, _5494, _5495, _5496, _5497, _5498, _5499, _5500, _5501, _5502, _5503, _5504, _5505, _5506, _5507, _5508, _5509, _5510, _5511, _5512, _5513, _5514, _5515, _5516, _5517, _5518, _5519, _5520, _5521, _5522, _5523, _5524, _5525, _5526, _5527, _5528, _5529, _5530, _5531, _5532, _5533, _5534, _5535, _5536, _5537, _5538, _5539, _5540, _5541, _5542, _5543, _5544, _5545, _5546, _5547, _5548, _5549, _5550, _5551, _5552, _5553, _5554, _5555, _5556, _5557, _5558, _5559, _5560, _5561, _5562, _5563, _5564, _5565, _5566, _5567, _5568, _5569, _5570, _5571, _5572, _5573, _5574, _5575, _5576, _5577, _5578, _5579, _5580, _5581, _5582, _5583, _5584, _5585, _5586, _5587, _5588, _5589, _5590, _5591, _5592, _5593, _5594, _5595, _5596, _5597, _5598, _5599, _5600, _5601, _5602, _5603, _5604, _5605, _5606, _5607, _5608, _5609, _5610, _5611, _5612, _5613, _5614, _5615, _5616, _5617, _5618, _5619, _5620, _5621, _5622, _5623, _5624, _5625, _5626, _5627, _5628, _5629, _5630, _5631, _5632, _5633, _5634, _5635, _5636, _5637, _5638, _5639, _5640, _5641, _5642, _5643, _5644, _5645, _5646, _5647, _5648, _5649, _5650, _5651, _5652, _5653, _5654, _5655, _5656, _5657, _5658, _5659, _5660, _5661, _5662, _5663, _5664, _5665, _5666, _5667, _5668, _5669, _5670, _5671, _5672, _5673, _5674, _5675, _5676, _5677, _5678, _5679, _5680, _5681, _5682, _5683, _5684, _5685, _5686, _5687, _5688, _5689, _5690, _5691, _5692, _5693, _5694, _5695, _5696, _5697, _5698, _5699, _5700, _5701, _5702, _5703, _5704, _5705, _5706, _5707;

assign o_1_ = ( n_n105 ) | ( _4425 ) ;
 assign o_2_ = ( n_n127 ) | ( _4553 ) ;
 assign o_0_ =((~ i_7_) & i_7_);
 assign o_12_ = ( wire4524 ) | ( _4617 ) ;
 assign o_11_ = ( n_n720 ) | ( _4689 ) ;
 assign o_14_ = ( n_n842 ) | ( _4759 ) ;
 assign o_13_ = ( wire4717 ) | ( _4819 ) ;
 assign o_16_ = ( wire4735 ) | ( _4832 ) ;
 assign o_15_ = ( _4854 ) | ( _4855 ) ;
 assign o_18_ = ( wire4767 ) | ( _4871 ) ;
 assign o_17_ = ( n_n912 ) | ( _4879 ) ;
 assign o_10_ = ( _4982 ) | ( _4983 ) ;
 assign o_9_ = ( n_n580 ) | ( _5108 ) ;
 assign o_7_ = ( n_n445 ) | ( _5223 ) ;
 assign o_8_ = ( n_n513 ) | ( _5328 ) ;
 assign o_5_ = ( wire5255 ) | ( _5438 ) ;
 assign o_6_ = ( n_n372 ) | ( _5544 ) ;
 assign o_3_ = ( n_n192 ) | ( _5619 ) ;
 assign o_4_ = ( n_n244 ) | ( _5707 ) ;
 assign n_n105 = ( _4409 ) | ( _4410 ) ;
 assign n_n127 = ( wire4354 ) | ( _4502 ) ;
 assign n_n720 = ( wire4608 ) | ( _4678 ) ;
 assign n_n842 = ( wire4664 ) | ( _4749 ) ;
 assign wire4717 = ( n_n804 ) | ( _4801 ) ;
 assign wire4735 = ( n_n904 ) | ( _4826 ) ;
 assign n_n889 = ( _4835 ) | ( _4836 ) ;
 assign wire4767 = ( n_n918 ) | ( _4865 ) ;
 assign n_n912 = ( _4876 ) | ( _4877 ) ;
 assign n_n580 = ( _5042 ) | ( _5043 ) ;
 assign n_n445 = ( wire5102 ) | ( _5166 ) ;
 assign n_n513 = ( wire5178 ) | ( _5279 ) ;
 assign n_n303 = ( wire5216 ) | ( _5379 ) ;
 assign n_n372 = ( wire5333 ) | ( _5496 ) ;
 assign n_n192 = ( _5601 ) | ( _5602 ) ;
 assign n_n244 = ( wire5444 ) | ( _5675 ) ;
 assign n_n1324 = ( n_n93  &  _38 ) ;
 assign n_n94 = ( (~ i_2_)  &  _305 ) ;
 assign n_n1176 = ( n_n91  &  _318 ) ;
 assign n_n78 = ( (~ i_6_)  &  n_n86 ) ;
 assign n_n1254 = ( n_n78  &  _308 ) ;
 assign n_n93 = ( i_6_  &  n_n86 ) ;
 assign n_n1132 = ( n_n93  &  _321 ) ;
 assign n_n92 = ( (~ i_4_)  &  _302 ) ;
 assign n_n1259 = ( n_n63  &  _308 ) ;
 assign wire4614 = ( _4709 ) | ( _4710 ) ;
 assign n_n856 = ( wire4614 ) | ( _4712 ) ;
 assign n_n855 = ( _4716 ) | ( _4717 ) ;
 assign n_n846 = ( _4723 ) | ( _4724 ) ;
 assign n_n999 = ( n_n93  &  _323 ) ;
 assign n_n97 = ( i_2_  &  _304 ) ;
 assign n_n1004 = ( n_n91  &  _44 ) ;
 assign n_n95 = ( i_6_  &  n_n64 ) ;
 assign n_n995 = ( n_n95  &  _311 ) ;
 assign n_n63 = ( (~ i_6_)  &  n_n75 ) ;
 assign n_n77 = ( i_5_  &  _35 ) ;
 assign n_n101 = ( i_6_  &  n_n70 ) ;
 assign n_n1216 = ( n_n101  &  _311 ) ;
 assign n_n975 = ( n_n84  &  _334 ) ;
 assign n_n987 = ( n_n93  &  _23 ) ;
 assign n_n504 = ( n_n984 ) | ( _4802 ) ;
 assign n_n964 = ( n_n95  &  _331 ) ;
 assign n_n814 = ( _4804 ) | ( _4805 ) ;
 assign n_n809 = ( _4765 ) | ( _4766 ) ;
 assign n_n804 = ( _4779 ) | ( _4780 ) ;
 assign n_n1060 = ( n_n63  &  _312 ) ;
 assign n_n83 = ( i_2_  &  _330 ) ;
 assign n_n58 = ( (~ i_6_)  &  n_n64 ) ;
 assign n_n1055 = ( n_n58  &  _299 ) ;
 assign n_n82 = ( (~ i_6_)  &  n_n70 ) ;
 assign n_n1160 = ( n_n81  &  _334 ) ;
 assign n_n1181 = ( n_n78  &  _299 ) ;
 assign n_n771 = ( _4570 ) | ( _4571 ) ;
 assign n_n874 = ( _136 ) | ( _913 ) ;
 assign n_n1092 = ( n_n91  &  _28 ) ;
 assign n_n730 = ( _4621 ) | ( _4622 ) ;
 assign n_n726 = ( _4683 ) | ( _4684 ) ;
 assign wire4608 = ( n_n722 ) | ( _4657 ) ;
 assign n_n81 = ( i_4_  &  _302 ) ;
 assign n_n1009 = ( n_n95  &  _25 ) ;
 assign n_n1011 = ( n_n103  &  _4432 ) ;
 assign n_n1087 = ( n_n63  &  _317 ) ;
 assign n_n1082 = ( n_n63  &  _44 ) ;
 assign n_n1217 = ( n_n101  &  _312 ) ;
 assign n_n84 = ( i_3_  &  _329 ) ;
 assign n_n951 = ( n_n92  &  _309 ) ;
 assign n_n956 = ( n_n78  &  _43 ) ;
 assign n_n943 = ( n_n93  &  _308 ) ;
 assign n_n676 = ( _4905 ) | ( _4906 ) ;
 assign n_n665 = ( _4885 ) | ( _4886 ) ;
 assign n_n658 = ( _4901 ) | ( _4902 ) ;
 assign n_n661 = ( _4920 ) | ( _4921 ) ;
 assign wire4879 = ( _4960 ) | ( _4961 ) ;
 assign n_n90 = ( i_2_  &  _306 ) ;
 assign n_n967 = ( n_n93  &  _24 ) ;
 assign n_n957 = ( n_n91  &  _41 ) ;
 assign n_n602 = ( _5012 ) | ( _5013 ) ;
 assign n_n591 = ( _5059 ) | ( _5060 ) ;
 assign n_n601 = ( _4987 ) | ( _4988 ) ;
 assign n_n584 = ( _5007 ) | ( _5008 ) ;
 assign wire4935 = ( n_n602 ) | ( _5021 ) ;
 assign n_n990 = ( n_n74  &  _350 ) ;
 assign n_n991 = ( n_n82  &  _25 ) ;
 assign n_n986 = ( n_n63  &  _316 ) ;
 assign n_n102 = ( (~ i_5_)  &  _314 ) ;
 assign n_n1100 = ( n_n82  &  _24 ) ;
 assign n_n1095 = ( n_n91  &  _27 ) ;
 assign n_n1184 = ( n_n95  &  _307 ) ;
 assign n_n96 = ( (~ i_4_)  &  _297 ) ;
 assign n_n1283 = ( n_n91  &  _321 ) ;
 assign n_n1058 = ( n_n58  &  _318 ) ;
 assign wire5164 = ( _5226 ) | ( _5227 ) ;
 assign n_n530 = ( _5244 ) | ( _5245 ) ;
 assign n_n529 = ( _5249 ) | ( _5250 ) ;
 assign n_n531 = ( _5255 ) | ( _5256 ) ;
 assign n_n71 = ( i_6_  &  _329 ) ;
 assign n_n968 = ( n_n80  &  _4492 ) ;
 assign n_n969 = ( n_n77  &  _319 ) ;
 assign n_n1045 = ( _307  &  _325 ) ;
 assign n_n1046 = ( n_n101  &  _38 ) ;
 assign n_n1043 = ( n_n91  &  _322 ) ;
 assign wire5034 = ( _5188 ) | ( _5189 ) ;
 assign n_n80 = ( i_0_  &  _4405 ) ;
 assign n_n953 = ( n_n79  &  _5014 ) ;
 assign n_n954 = ( n_n78  &  _317 ) ;
 assign n_n952 = ( n_n81  &  _352 ) ;
 assign n_n54 = ( (~ i_6_)  &  _313 ) ;
 assign n_n1006 = ( n_n95  &  _318 ) ;
 assign n_n1074 = ( n_n101  &  _318 ) ;
 assign n_n91 = ( i_6_  &  n_n75 ) ;
 assign n_n1077 = ( n_n91  &  _311 ) ;
 assign n_n1068 = ( n_n95  &  _34 ) ;
 assign n_n1169 = ( n_n91  &  _38 ) ;
 assign n_n1088 = ( n_n91  &  _349 ) ;
 assign wire5324 = ( _5442 ) | ( _5443 ) ;
 assign n_n1047 = ( n_n63  &  _301 ) ;
 assign n_n1042 = ( n_n92  &  _30 ) ;
 assign n_n87 = ( (~ i_6_)  &  _328 ) ;
 assign n_n1147 = ( _339  &  _340 ) ;
 assign n_n994 = ( n_n91  &  _310 ) ;
 assign n_n322 = ( _5402 ) | ( _5403 ) ;
 assign n_n311 = ( _5333 ) | ( _5334 ) ;
 assign n_n958 = ( n_n77  &  _351 ) ;
 assign n_n962 = ( n_n74  &  _348 ) ;
 assign n_n1048 = ( n_n95  &  _299 ) ;
 assign n_n1164 = ( n_n93  &  _43 ) ;
 assign n_n1105 = ( n_n58  &  _317 ) ;
 assign n_n257 = ( _5624 ) | ( _5625 ) ;
 assign wire5389 = ( _5678 ) | ( _5679 ) ;
 assign wire5393 = ( _5682 ) | ( _5683 ) ;
 assign n_n252 = ( wire5393 ) | ( _5685 ) ;
 assign n_n254 = ( _5690 ) | ( _5691 ) ;
 assign n_n246 = ( _5694 ) | ( _5695 ) ;
 assign n_n66 = ( i_6_  &  _313 ) ;
 assign n_n974 = ( n_n66  &  _4907 ) ;
 assign n_n980 = ( n_n84  &  _309 ) ;
 assign n_n67 = ( (~ i_3_)  &  _330 ) ;
 assign n_n1146 = ( n_n96  &  _335 ) ;
 assign n_n1145 = ( _31  &  _314 ) ;
 assign n_n40 = ( i_4_  &  _4385 ) ;
 assign n_n1122 = ( n_n101  &  _331 ) ;
 assign wire5337 = ( _5547 ) | ( _5548 ) ;
 assign n_n205 = ( _5553 ) | ( _5554 ) ;
 assign n_n195 = ( _5563 ) | ( _5564 ) ;
 assign n_n202 = ( _5568 ) | ( _5569 ) ;
 assign n_n208 = ( _5573 ) | ( _5574 ) ;
 assign n_n196 = ( _5585 ) | ( _5586 ) ;
 assign n_n1022 = ( n_n58  &  _322 ) ;
 assign n_n1204 = ( n_n95  &  _354 ) ;
 assign wire4411 = ( _4508 ) | ( _4509 ) ;
 assign n_n144 = ( _4441 ) | ( _4442 ) ;
 assign n_n131 = ( n_n143 ) | ( _4459 ) ;
 assign n_n141 = ( _4467 ) | ( _4468 ) ;
 assign n_n147 = ( _4430 ) | ( _4431 ) ;
 assign wire4354 = ( n_n131 ) | ( _4484 ) ;
 assign n_n106 = ( _4415 ) | ( _4416 ) ;
 assign n_n99 = ( (~ i_4_)  &  _303 ) ;
 assign n_n100 = ( (~ i_2_)  &  _330 ) ;
 assign n_n939 = ( _327  &  _357 ) ;
 assign n_n85 = ( (~ i_2_)  &  _304 ) ;
 assign n_n79 = ( (~ i_6_)  &  _329 ) ;
 assign n_n86 = ( (~ i_7_)  &  (~ i_8_) ) ;
 assign n_n76 = ( (~ i_6_)  &  _302 ) ;
 assign n_n75 = ( (~ i_7_)  &  i_8_ ) ;
 assign n_n960 = ( n_n75  &  _358 ) ;
 assign n_n74 = ( (~ i_5_)  &  _35 ) ;
 assign n_n103 = ( i_2_  &  _305 ) ;
 assign n_n973 = ( n_n82  &  _312 ) ;
 assign n_n981 = ( n_n95  &  _45 ) ;
 assign n_n989 = ( n_n91  &  _317 ) ;
 assign n_n1134 = ( n_n58  &  _311 ) ;
 assign n_n1163 = ( n_n84  &  _32 ) ;
 assign n_n1172 = ( n_n95  &  _301 ) ;
 assign n_n64 = ( i_7_  &  i_8_ ) ;
 assign n_n937 = ( (~ i_2_)  &  _306 ) ;
 assign wire4762 = ( _4858 ) | ( _4859 ) ;
 assign n_n918 = ( wire4762 ) | ( _4861 ) ;
 assign n_n1109 = ( n_n101  &  _46 ) ;
 assign n_n1032 = ( n_n93  &  _46 ) ;
 assign wire4743 = ( _4839 ) | ( _4840 ) ;
 assign n_n890 = ( _4844 ) | ( _4845 ) ;
 assign n_n892 = ( _4849 ) | ( _4850 ) ;
 assign n_n853 = ( _4728 ) | ( _4729 ) ;
 assign n_n852 = ( _4734 ) | ( _4735 ) ;
 assign n_n854 = ( _4740 ) | ( _4741 ) ;
 assign n_n950 = ( n_n95  &  _310 ) ;
 assign n_n955 = ( n_n99  &  _4554 ) ;
 assign n_n940 = ( n_n95  &  _43 ) ;
 assign n_n815 = ( _4809 ) | ( _4810 ) ;
 assign n_n941 = ( n_n96  &  _30 ) ;
 assign n_n1040 = ( n_n96  &  _351 ) ;
 assign n_n1039 = ( n_n78  &  _36 ) ;
 assign n_n1128 = ( n_n78  &  _307 ) ;
 assign wire4462 = ( _4574 ) | ( _4575 ) ;
 assign n_n1085 = ( n_n63  &  _36 ) ;
 assign n_n1091 = ( _336  &  _343 ) ;
 assign n_n1078 = ( n_n78  &  _300 ) ;
 assign n_n1153 = ( n_n58  &  _38 ) ;
 assign n_n1170 = ( n_n93  &  _41 ) ;
 assign n_n554 = ( _167 ) | ( _4630 ) ;
 assign wire4570 = ( _4633 ) | ( _4634 ) ;
 assign n_n732 = ( _4627 ) | ( _4628 ) ;
 assign n_n727 = ( _4639 ) | ( _4640 ) ;
 assign n_n722 = ( _4647 ) | ( _4648 ) ;
 assign n_n735 = ( _4662 ) | ( _4663 ) ;
 assign n_n1018 = ( n_n95  &  _24 ) ;
 assign n_n1081 = ( _39  &  _344 ) ;
 assign n_n664 = ( _4969 ) | ( _4970 ) ;
 assign n_n662 = ( _4973 ) | ( _4974 ) ;
 assign n_n666 = ( _4891 ) | ( _4892 ) ;
 assign n_n652 = ( _178 ) | ( _5015 ) ;
 assign n_n590 = ( _5065 ) | ( _5066 ) ;
 assign n_n588 = ( _5047 ) | ( _5048 ) ;
 assign n_n587 = ( _5052 ) | ( _5053 ) ;
 assign wire4956 = ( _5055 ) | ( _5056 ) ;
 assign n_n1001 = ( n_n63  &  _300 ) ;
 assign n_n993 = ( _25  &  _338 ) ;
 assign n_n1079 = ( n_n93  &  _320 ) ;
 assign n_n1193 = ( n_n58  &  _307 ) ;
 assign n_n1188 = ( n_n58  &  _301 ) ;
 assign n_n1279 = ( n_n78  &  _46 ) ;
 assign wire5168 = ( _5230 ) | ( _5231 ) ;
 assign n_n527 = ( wire5168 ) | ( _5233 ) ;
 assign n_n533 = ( _5260 ) | ( _5261 ) ;
 assign n_n532 = ( _5266 ) | ( _5267 ) ;
 assign n_n518 = ( _5271 ) | ( _5272 ) ;
 assign n_n971 = ( n_n100  &  _4664 ) ;
 assign n_n1035 = ( n_n74  &  _335 ) ;
 assign wire5060 = ( _5111 ) | ( _5112 ) ;
 assign n_n466 = ( wire5060 ) | ( _5114 ) ;
 assign n_n465 = ( _5118 ) | ( _5119 ) ;
 assign n_n654 = ( n_n939 ) | ( _222 ) ;
 assign n_n451 = ( _5122 ) | ( _5123 ) ;
 assign n_n947 = ( _305  &  _339 ) ;
 assign n_n944 = ( n_n91  &  _23 ) ;
 assign n_n1013 = ( n_n93  &  _337 ) ;
 assign n_n1010 = ( n_n78  &  _33 ) ;
 assign n_n421 = ( _693 ) | ( _5144 ) ;
 assign n_n1177 = ( n_n78  &  _316 ) ;
 assign n_n390 = ( _5510 ) | ( _5511 ) ;
 assign n_n389 = ( _5516 ) | ( _5517 ) ;
 assign wire5268 = ( _5520 ) | ( _5521 ) ;
 assign n_n1144 = ( (~ i_1_)  &  _324 ) ;
 assign n_n977 = ( n_n67  &  _360 ) ;
 assign n_n983 = ( n_n95  &  _357 ) ;
 assign n_n970 = ( n_n85  &  _4908 ) ;
 assign n_n365 = ( _58 ) | ( _5380 ) ;
 assign n_n1331 = ( n_n91  &  _46 ) ;
 assign n_n310 = ( _5337 ) | ( _5338 ) ;
 assign n_n942 = ( n_n91  &  _316 ) ;
 assign n_n1057 = ( n_n82  &  _301 ) ;
 assign n_n1156 = ( n_n91  &  _331 ) ;
 assign wire5415 = ( _5629 ) | ( _5630 ) ;
 assign n_n256 = ( wire5415 ) | ( _5632 ) ;
 assign wire5420 = ( _5637 ) | ( _5638 ) ;
 assign n_n984 = ( n_n63  &  _310 ) ;
 assign wire5341 = ( _5557 ) | ( _5558 ) ;
 assign n_n204 = ( wire5341 ) | ( _5560 ) ;
 assign n_n198 = ( _5606 ) | ( _5607 ) ;
 assign n_n1330 = ( n_n95  &  _38 ) ;
 assign n_n137 = ( _4515 ) | ( _4516 ) ;
 assign n_n134 = ( _4521 ) | ( _4522 ) ;
 assign n_n133 = ( _4527 ) | ( _4528 ) ;
 assign n_n135 = ( _4537 ) | ( _4538 ) ;
 assign n_n128 = ( n_n135 ) | ( _4539 ) ;
 assign wire4164 = ( _4419 ) | ( _4420 ) ;
 assign n_n70 = ( i_7_  &  (~ i_8_) ) ;
 assign n_n982 = ( n_n81  &  _319 ) ;
 assign n_n52 = ( i_7_  &  i_6_ ) ;
 assign n_n73 = ( (~ i_7_)  &  (~ i_6_) ) ;
 assign n_n1173 = ( n_n91  &  _323 ) ;
 assign n_n946 = ( _315  &  _4607 ) ;
 assign n_n1125 = ( n_n78  &  _301 ) ;
 assign wire4670 = ( _4752 ) | ( _4753 ) ;
 assign n_n966 = ( n_n101  &  _23 ) ;
 assign n_n1070 = ( n_n99  &  _30 ) ;
 assign n_n812 = ( _4785 ) | ( _4786 ) ;
 assign wire4681 = ( _4789 ) | ( _4790 ) ;
 assign n_n811 = ( wire4681 ) | ( _4792 ) ;
 assign wire4685 = ( _4795 ) | ( _4796 ) ;
 assign n_n1036 = ( n_n91  &  _312 ) ;
 assign n_n1075 = ( n_n96  &  _4462 ) ;
 assign n_n1185 = ( n_n78  &  _28 ) ;
 assign n_n728 = ( _4645 ) | ( _4646 ) ;
 assign n_n949 = ( n_n101  &  _45 ) ;
 assign wire4873 = ( _4913 ) | ( _4914 ) ;
 assign wire4813 = ( _4897 ) | ( _4898 ) ;
 assign n_n670 = ( _4926 ) | ( _4927 ) ;
 assign n_n1267 = ( n_n101  &  _28 ) ;
 assign wire5003 = ( n_n582 ) | ( _5080 ) ;
 assign n_n978 = ( n_n92  &  _333 ) ;
 assign n_n53 = ( i_1_  &  _296 ) ;
 assign n_n1158 = ( n_n78  &  _323 ) ;
 assign wire5176 = ( _5237 ) | ( _5238 ) ;
 assign n_n526 = ( wire5176 ) | ( _5241 ) ;
 assign wire5108 = ( _5299 ) | ( _5300 ) ;
 assign n_n523 = ( _5306 ) | ( _5307 ) ;
 assign n_n525 = ( _5310 ) | ( _5311 ) ;
 assign n_n959 = ( n_n91  &  _33 ) ;
 assign wire5010 = ( _5172 ) | ( _5173 ) ;
 assign wire5056 = ( _5197 ) | ( _5198 ) ;
 assign wire5102 = ( n_n451 ) | ( _5143 ) ;
 assign n_n1014 = ( n_n78  &  _320 ) ;
 assign n_n1294 = ( n_n78  &  _353 ) ;
 assign n_n1028 = ( n_n63  &  _332 ) ;
 assign n_n1130 = ( n_n58  &  _45 ) ;
 assign n_n320 = ( _5407 ) | ( _5408 ) ;
 assign n_n1215 = ( n_n58  &  _354 ) ;
 assign wire5192 = ( _5341 ) | ( _5342 ) ;
 assign wire5216 = ( _5354 ) | ( _5355 ) ;
 assign n_n309 = ( _5396 ) | ( _5397 ) ;
 assign wire5255 = ( n_n308 ) | ( _5437 ) ;
 assign n_n1030 = ( n_n81  &  _309 ) ;
 assign n_n259 = ( _5642 ) | ( _5643 ) ;
 assign n_n258 = ( _5648 ) | ( _5649 ) ;
 assign n_n295 = ( n_n1002 ) | ( _632 ) ;
 assign n_n248 = ( _5653 ) | ( _5654 ) ;
 assign n_n1019 = ( _351  &  _5124 ) ;
 assign n_n1020 = ( n_n101  &  _4623 ) ;
 assign n_n136 = ( _4545 ) | ( _4546 ) ;
 assign n_n1281 = ( n_n91  &  _337 ) ;
 assign wire4181 = ( _4389 ) | ( _4390 ) ;
 assign n_n1093 = ( n_n75  &  _346 ) ;
 assign n_n1103 = ( n_n102  &  _350 ) ;
 assign n_n1297 = ( n_n95  &  _321 ) ;
 assign n_n1286 = ( n_n58  &  _316 ) ;
 assign n_n1369 = ( n_n63  &  _4613 ) ;
 assign wire4715 = ( _4813 ) | ( _4814 ) ;
 assign wire4690 = ( _4769 ) | ( _4770 ) ;
 assign n_n808 = ( wire4690 ) | ( _4772 ) ;
 assign wire4694 = ( _4775 ) | ( _4776 ) ;
 assign n_n1021 = ( n_n96  &  _352 ) ;
 assign n_n1054 = ( _29  &  _40 ) ;
 assign n_n961 = ( n_n95  &  _47 ) ;
 assign n_n716 = ( n_n959 ) | ( _4718 ) ;
 assign wire4877 = ( _4915 ) | ( _4916 ) ;
 assign n_n663 = ( _4978 ) | ( _4979 ) ;
 assign n_n582 = ( _5073 ) | ( _5074 ) ;
 assign n_n595 = ( _5089 ) | ( _5090 ) ;
 assign n_n1025 = ( n_n74  &  _309 ) ;
 assign n_n1026 = ( _4433  &  _4434 ) ;
 assign wire5017 = ( _5176 ) | ( _5177 ) ;
 assign n_n453 = ( wire5017 ) | ( _5180 ) ;
 assign n_n455 = ( _5184 ) | ( _5185 ) ;
 assign n_n446 = ( wire5034 ) | ( _5194 ) ;
 assign n_n458 = ( wire5054 ) | ( _5206 ) ;
 assign n_n1120 = ( n_n92  &  _350 ) ;
 assign n_n1117 = ( _31  &  _4474 ) ;
 assign n_n1002 = ( i_0_  &  _324 ) ;
 assign n_n321 = ( _5413 ) | ( _5414 ) ;
 assign wire5198 = ( _5346 ) | ( _5347 ) ;
 assign n_n312 = ( wire5198 ) | ( _5349 ) ;
 assign n_n206 = ( _5579 ) | ( _5580 ) ;
 assign n_n1174 = ( n_n93  &  _300 ) ;
 assign n_n109 = ( _4395 ) | ( _4396 ) ;
 assign n_n775 = ( _4558 ) | ( _4559 ) ;
 assign n_n773 = ( _4581 ) | ( _4582 ) ;
 assign n_n770 = ( _4587 ) | ( _4588 ) ;
 assign n_n765 = ( n_n768 ) | ( _4601 ) ;
 assign n_n774 = ( _4564 ) | ( _4565 ) ;
 assign wire4524 = ( n_n765 ) | ( _4606 ) ;
 assign n_n1052 = ( n_n63  &  _318 ) ;
 assign n_n669 = ( _4932 ) | ( _4933 ) ;
 assign n_n598 = ( _4993 ) | ( _4994 ) ;
 assign n_n521 = ( _5284 ) | ( _5285 ) ;
 assign wire5042 = ( _5210 ) | ( _5211 ) ;
 assign wire5048 = ( _5214 ) | ( _5215 ) ;
 assign n_n456 = ( wire5048 ) | ( _5217 ) ;
 assign wire5054 = ( _5203 ) | ( _5204 ) ;
 assign n_n976 = ( _338  &  _359 ) ;
 assign n_n1121 = ( n_n90  &  _4934 ) ;
 assign wire5203 = ( _5358 ) | ( _5359 ) ;
 assign n_n315 = ( wire5203 ) | ( _5361 ) ;
 assign n_n308 = ( n_n321 ) | ( _5415 ) ;
 assign n_n319 = ( wire5242 ) | ( _5421 ) ;
 assign n_n325 = ( _5385 ) | ( _5386 ) ;
 assign wire5444 = ( n_n248 ) | ( _5659 ) ;
 assign wire5365 = ( _5582 ) | ( _5583 ) ;
 assign n_n882 = ( _181 ) | ( _4485 ) ;
 assign n_n145 = ( _4490 ) | ( _4491 ) ;
 assign wire4211 = ( _4400 ) | ( _4401 ) ;
 assign n_n110 = ( wire4211 ) | ( _4404 ) ;
 assign n_n1108 = ( n_n93  &  _301 ) ;
 assign n_n1118 = ( n_n91  &  _4935 ) ;
 assign n_n849 = ( _4694 ) | ( _4695 ) ;
 assign n_n776 = ( _4611 ) | ( _4612 ) ;
 assign n_n668 = ( _4938 ) | ( _4939 ) ;
 assign n_n641 = ( _76 ) | ( _4940 ) ;
 assign n_n599 = ( _5027 ) | ( _5028 ) ;
 assign wire5130 = ( _5289 ) | ( _5290 ) ;
 assign wire5208 = ( _5365 ) | ( _5366 ) ;
 assign n_n314 = ( wire5208 ) | ( _5368 ) ;
 assign n_n250 = ( _5697 ) | ( _5698 ) ;
 assign n_n146 = ( _4499 ) | ( _4500 ) ;
 assign n_n850 = ( _4700 ) | ( _4701 ) ;
 assign n_n734 = ( _4669 ) | ( _4670 ) ;
 assign n_n733 = ( _4675 ) | ( _4676 ) ;
 assign n_n671 = ( _4944 ) | ( _4945 ) ;
 assign n_n672 = ( _4950 ) | ( _4951 ) ;
 assign wire4836 = ( _4955 ) | ( _4956 ) ;
 assign n_n1101 = ( n_n70  &  _346 ) ;
 assign n_n600 = ( _5033 ) | ( _5034 ) ;
 assign wire4985 = ( _5092 ) | ( _5093 ) ;
 assign wire4977 = ( _5069 ) | ( _5070 ) ;
 assign n_n1312 = ( n_n101  &  _321 ) ;
 assign n_n519 = ( _5314 ) | ( _5315 ) ;
 assign n_n520 = ( _5295 ) | ( _5296 ) ;
 assign wire5136 = ( _5320 ) | ( _5321 ) ;
 assign n_n463 = ( _5128 ) | ( _5129 ) ;
 assign wire5079 = ( _5133 ) | ( _5134 ) ;
 assign n_n464 = ( _5137 ) | ( _5138 ) ;
 assign n_n324 = ( _5390 ) | ( _5391 ) ;
 assign wire5234 = ( _5424 ) | ( _5425 ) ;
 assign wire5214 = ( _5373 ) | ( _5374 ) ;
 assign n_n140 = ( _4472 ) | ( _4473 ) ;
 assign wire4662 = ( _4705 ) | ( _4706 ) ;
 assign n_n769 = ( _4593 ) | ( _4594 ) ;
 assign n_n768 = ( _4599 ) | ( _4600 ) ;
 assign wire4556 = ( _4651 ) | ( _4652 ) ;
 assign n_n594 = ( _5101 ) | ( _5102 ) ;
 assign wire5178 = ( n_n518 ) | ( _5274 ) ;
 assign n_n460 = ( _5149 ) | ( _5150 ) ;
 assign wire5092 = ( _5153 ) | ( _5154 ) ;
 assign n_n459 = ( wire5092 ) | ( _5156 ) ;
 assign wire5100 = ( _5160 ) | ( _5161 ) ;
 assign n_n318 = ( _5430 ) | ( _5431 ) ;
 assign wire5242 = ( _5418 ) | ( _5419 ) ;
 assign wire5405 = ( _5701 ) | ( _5702 ) ;
 assign wire4296 = ( _4478 ) | ( _4479 ) ;
 assign n_n1059 = ( _344  &  _4443 ) ;
 assign n_n395 = ( _5499 ) | ( _5500 ) ;
 assign wire5294 = ( _5452 ) | ( _5453 ) ;
 assign n_n384 = ( wire5294 ) | ( _5455 ) ;
 assign n_n392 = ( _5527 ) | ( _5528 ) ;
 assign n_n378 = ( _5537 ) | ( _5538 ) ;
 assign n_n379 = ( _5505 ) | ( _5506 ) ;
 assign wire5290 = ( n_n378 ) | ( _5543 ) ;
 assign wire5437 = ( _5662 ) | ( _5663 ) ;
 assign n_n262 = ( wire5437 ) | ( _5665 ) ;
 assign n_n261 = ( _5669 ) | ( _5670 ) ;
 assign n_n904 = ( _4824 ) | ( _4825 ) ;
 assign wire5301 = ( _5458 ) | ( _5459 ) ;
 assign n_n385 = ( wire5301 ) | ( _5461 ) ;
 assign n_n374 = ( n_n382 ) | ( _5477 ) ;
 assign n_n386 = ( wire5331 ) | ( _5449 ) ;
 assign wire5333 = ( _5485 ) | ( _5486 ) ;
 assign wire5375 = ( _5611 ) | ( _5612 ) ;
 assign n_n199 = ( wire5375 ) | ( _5614 ) ;
 assign n_n142 = ( _4450 ) | ( _4451 ) ;
 assign n_n393 = ( _5532 ) | ( _5533 ) ;
 assign n_n382 = ( _5466 ) | ( _5467 ) ;
 assign wire5306 = ( _5480 ) | ( _5481 ) ;
 assign n_n143 = ( _4457 ) | ( _4458 ) ;
 assign wire5315 = ( _5470 ) | ( _5471 ) ;
 assign wire4664 = ( n_n846 ) | ( _4743 ) ;
 assign wire5350 = ( _5589 ) | ( _5590 ) ;
 assign n_n201 = ( _5595 ) | ( _5596 ) ;
 assign wire4934 = ( _282 ) | ( _5038 ) ;
 assign n_n388 = ( _5490 ) | ( _5491 ) ;
 assign wire5331 = ( _5446 ) | ( _5447 ) ;
 assign wire4909 = ( _4997 ) | ( _4998 ) ;
 assign n_n596 = ( wire4909 ) | ( _5000 ) ;
 assign wire4914 = ( _5003 ) | ( _5004 ) ;
 assign _19 = ( n_n77  &  n_n103 ) ;
 assign _20 = ( n_n93  &  n_n85 ) ;
 assign _21 = ( n_n83  &  n_n99 ) ;
 assign _22 = ( n_n97  &  n_n81 ) ;
 assign _23 = ( n_n97  &  n_n102 ) ;
 assign _24 = ( n_n77  &  n_n100 ) ;
 assign _25 = ( n_n81  &  n_n103 ) ;
 assign _26 = ( i_3_  &  i_2_ ) ;
 assign _27 = ( n_n92  &  n_n103 ) ;
 assign _28 = ( n_n84  &  n_n100 ) ;
 assign _29 = ( n_n84  &  n_n103 ) ;
 assign _30 = ( n_n94  &  n_n93 ) ;
 assign _31 = ( n_n94  &  n_n82 ) ;
 assign _32 = ( n_n83  &  n_n91 ) ;
 assign _33 = ( n_n97  &  n_n84 ) ;
 assign _34 = ( n_n99  &  n_n85 ) ;
 assign _35 = ( (~ i_3_)  &  i_4_ ) ;
 assign _36 = ( n_n94  &  n_n102 ) ;
 assign _37 = ( n_n77  &  n_n90 ) ;
 assign _38 = ( n_n90  &  n_n102 ) ;
 assign _39 = ( n_n54  &  n_n64 ) ;
 assign _40 = ( i_7_  &  (~ i_6_) ) ;
 assign _41 = ( n_n92  &  n_n100 ) ;
 assign _42 = ( n_n92  &  n_n85 ) ;
 assign _43 = ( n_n97  &  n_n96 ) ;
 assign _44 = ( n_n97  &  n_n74 ) ;
 assign _45 = ( n_n84  &  n_n85 ) ;
 assign _46 = ( n_n90  &  n_n74 ) ;
 assign _47 = ( n_n102  &  n_n100 ) ;
 assign _48 = ( n_n101  &  _347 ) ;
 assign _49 = ( _1034 ) | ( _1035 ) ;
 assign _50 = ( n_n95  &  _347 ) ;
 assign _51 = ( n_n52  &  _316 ) ;
 assign _52 = ( n_n966 ) | ( _287 ) ;
 assign _53 = ( n_n79  &  _4713 ) ;
 assign _54 = ( _289 ) | ( _901 ) ;
 assign _55 = ( n_n102  &  _334 ) ;
 assign _56 = ( _293 ) | ( _848 ) ;
 assign _57 = ( n_n962 ) | ( _778 ) ;
 assign _58 = ( n_n67  &  _4984 ) ;
 assign _59 = ( n_n91  &  _307 ) ;
 assign _60 = ( _326  &  _349 ) ;
 assign _61 = ( n_n87  &  _355 ) ;
 assign _62 = ( n_n54  &  _5130 ) ;
 assign _63 = ( n_n63  &  _349 ) ;
 assign _64 = ( n_n101  &  _301 ) ;
 assign _65 = ( n_n1185 ) | ( _1054 ) ;
 assign _66 = ( n_n95  &  _317 ) ;
 assign _67 = ( n_n78  &  _310 ) ;
 assign _68 = ( n_n71  &  _355 ) ;
 assign _69 = ( n_n40  &  _4460 ) ;
 assign _70 = ( _968 ) | ( _969 ) ;
 assign _71 = ( n_n100  &  _336 ) ;
 assign _72 = ( n_n78  &  _321 ) ;
 assign _73 = ( n_n77  &  _333 ) ;
 assign _74 = ( n_n84  &  _333 ) ;
 assign _75 = ( n_n78  &  _337 ) ;
 assign _76 = ( n_n100  &  _4402 ) ;
 assign _77 = ( n_n96  &  _4946 ) ;
 assign _78 = ( n_n77  &  _335 ) ;
 assign _79 = ( n_n91  &  _320 ) ;
 assign _80 = ( n_n102  &  _309 ) ;
 assign _81 = ( n_n101  &  _323 ) ;
 assign _82 = ( n_n58  &  _331 ) ;
 assign _83 = ( n_n82  &  _311 ) ;
 assign _84 = ( n_n63  &  _359 ) ;
 assign _85 = ( _299  &  _327 ) ;
 assign _86 = ( _422 ) | ( _423 ) ;
 assign _87 = ( n_n93 ) | ( n_n101 ) ;
 assign _88 = ( _986 ) | ( _987 ) ;
 assign _89 = ( n_n947 ) | ( _769 ) ;
 assign _90 = ( _290 ) | ( _988 ) ;
 assign _91 = ( _634 ) | ( _635 ) ;
 assign _92 = ( _796 ) | ( _797 ) ;
 assign _93 = ( n_n91  &  _308 ) ;
 assign _94 = ( _1052 ) | ( _1053 ) ;
 assign _95 = ( n_n82  &  _308 ) ;
 assign _96 = ( n_n941 ) | ( n_n942 ) ;
 assign _97 = ( n_n954 ) | ( n_n952 ) ;
 assign _98 = ( n_n999 ) | ( _522 ) ;
 assign _99 = ( n_n975 ) | ( n_n973 ) ;
 assign _100 = ( _343  &  _4760 ) ;
 assign _102 = ( n_n1082 ) | ( _1019 ) ;
 assign _103 = ( _21  &  _338 ) ;
 assign _104 = ( _958 ) | ( _959 ) ;
 assign _107 = ( n_n53  &  _356 ) ;
 assign _108 = ( n_n95  &  _320 ) ;
 assign _109 = ( n_n91  &  _354 ) ;
 assign _110 = ( n_n78  &  _322 ) ;
 assign _111 = ( n_n75  &  _323 ) ;
 assign _112 = ( _767 ) | ( _768 ) ;
 assign _113 = ( n_n81  &  _335 ) ;
 assign _114 = ( n_n84  &  _4475 ) ;
 assign _115 = ( n_n70  &  _322 ) ;
 assign _116 = ( _284 ) | ( _876 ) ;
 assign _117 = ( n_n92  &  _319 ) ;
 assign _119 = ( n_n95  &  _300 ) ;
 assign _121 = ( n_n63  &  _337 ) ;
 assign _122 = ( n_n101  &  _308 ) ;
 assign _123 = ( n_n73  &  _347 ) ;
 assign _124 = ( n_n66  &  _5199 ) ;
 assign _125 = ( n_n93  &  _353 ) ;
 assign _126 = ( n_n53  &  _4922 ) ;
 assign _127 = ( n_n70  &  _307 ) ;
 assign _128 = ( n_n81  &  _4397 ) ;
 assign _129 = ( n_n82  &  _4436 ) ;
 assign _130 = ( _288 ) | ( _852 ) ;
 assign _131 = ( n_n92  &  _31 ) ;
 assign _132 = ( n_n983 ) | ( n_n982 ) ;
 assign _133 = ( n_n1279 ) | ( n_n1281 ) ;
 assign _134 = ( n_n82  &  _22 ) ;
 assign _135 = ( n_n84  &  _30 ) ;
 assign _136 = ( n_n1109 ) | ( _915 ) ;
 assign _137 = ( n_n102  &  _4529 ) ;
 assign _138 = ( n_n103  &  _4881 ) ;
 assign _140 = ( n_n58  &  _25 ) ;
 assign _142 = ( n_n78  &  _29 ) ;
 assign _143 = ( n_n95  &  _21 ) ;
 assign _144 = ( n_n1018 ) | ( n_n1021 ) ;
 assign _145 = ( n_n1035 ) | ( n_n1036 ) ;
 assign _147 = ( n_n82  &  _23 ) ;
 assign _148 = ( n_n95  &  _33 ) ;
 assign _149 = ( n_n101  &  _44 ) ;
 assign _150 = ( _794 ) | ( _795 ) ;
 assign _151 = ( n_n95  &  _41 ) ;
 assign _152 = ( n_n1048 ) | ( _1032 ) ;
 assign _153 = ( n_n103  &  _5512 ) ;
 assign _154 = ( n_n91  &  _29 ) ;
 assign _155 = ( n_n63  &  _43 ) ;
 assign _156 = ( n_n103  &  _5286 ) ;
 assign _157 = ( n_n78  &  _24 ) ;
 assign _158 = ( n_n92  &  _20 ) ;
 assign _159 = ( n_n77  &  _32 ) ;
 assign _160 = ( n_n93  &  _44 ) ;
 assign _161 = ( n_n102  &  _20 ) ;
 assign _162 = ( _356  &  _4503 ) ;
 assign _163 = ( n_n82  &  _19 ) ;
 assign _164 = ( n_n63  &  _19 ) ;
 assign _165 = ( _765 ) | ( _766 ) ;
 assign _166 = ( n_n99  &  _4744 ) ;
 assign _167 = ( n_n85  &  _4629 ) ;
 assign _168 = ( n_n52  &  _36 ) ;
 assign _169 = ( n_n93  &  _19 ) ;
 assign _170 = ( _348  &  _4530 ) ;
 assign _171 = ( n_n74  &  _32 ) ;
 assign _172 = ( n_n100  &  _4531 ) ;
 assign _173 = ( n_n95  &  _46 ) ;
 assign _174 = ( n_n90  &  _4962 ) ;
 assign _176 = ( _291 ) | ( _899 ) ;
 assign _177 = ( n_n95  &  _28 ) ;
 assign _178 = ( n_n95  &  _23 ) ;
 assign _180 = ( n_n100  &  _5075 ) ;
 assign _181 = ( n_n78  &  _23 ) ;
 assign _182 = ( n_n91  &  _24 ) ;
 assign _183 = ( n_n93  &  _37 ) ;
 assign _184 = ( n_n52  &  _22 ) ;
 assign _185 = ( n_n63  &  _23 ) ;
 assign _186 = ( n_n91  &  _36 ) ;
 assign _187 = ( _39  &  _4532 ) ;
 assign _188 = ( n_n101  &  _27 ) ;
 assign _189 = ( n_n1267 ) | ( _911 ) ;
 assign _190 = ( n_n63  &  _45 ) ;
 assign _191 = ( _39  &  _5167 ) ;
 assign _192 = ( n_n74  &  _5168 ) ;
 assign _193 = ( n_n63  &  _5322 ) ;
 assign _194 = ( n_n91  &  _43 ) ;
 assign _195 = ( _360  &  _4452 ) ;
 assign _196 = ( n_n91  &  _5157 ) ;
 assign _197 = ( _336  &  _5178 ) ;
 assign _198 = ( n_n82  &  _21 ) ;
 assign _199 = ( n_n91  &  _45 ) ;
 assign _200 = ( n_n1040 ) | ( _1030 ) ;
 assign _201 = ( _39  &  _4702 ) ;
 assign _202 = ( n_n97  &  _5200 ) ;
 assign _203 = ( n_n1369 ) | ( _923 ) ;
 assign _204 = ( n_n1312 ) | ( _850 ) ;
 assign _205 = ( n_n1312 ) | ( _581 ) ;
 assign _206 = ( n_n937 ) | ( n_n946 ) ;
 assign _207 = ( n_n941 ) | ( _925 ) ;
 assign _208 = ( n_n58  &  _36 ) ;
 assign _209 = ( n_n968 ) | ( n_n969 ) ;
 assign _210 = ( n_n960 ) | ( n_n961 ) ;
 assign _211 = ( n_n987 ) | ( n_n989 ) ;
 assign _212 = ( n_n1028 ) | ( n_n1030 ) ;
 assign _213 = ( n_n1020 ) | ( n_n1025 ) ;
 assign _214 = ( n_n951 ) | ( n_n949 ) ;
 assign _215 = ( n_n964 ) | ( n_n967 ) ;
 assign _216 = ( n_n52  &  _34 ) ;
 assign _217 = ( n_n1042 ) | ( n_n1040 ) ;
 assign _218 = ( n_n1160 ) | ( n_n1163 ) ;
 assign _219 = ( n_n1009 ) | ( n_n1013 ) ;
 assign _220 = ( n_n76  &  _4486 ) ;
 assign _221 = ( n_n956 ) | ( n_n958 ) ;
 assign _222 = ( n_n940 ) | ( _854 ) ;
 assign _223 = ( n_n101  &  _29 ) ;
 assign _224 = ( n_n99  &  _5061 ) ;
 assign _226 = ( n_n1039 ) | ( _520 ) ;
 assign _227 = ( n_n1046 ) | ( n_n1047 ) ;
 assign _228 = ( n_n82  &  _38 ) ;
 assign _230 = ( n_n63  &  _47 ) ;
 assign _231 = ( n_n74  &  _30 ) ;
 assign _232 = ( n_n91  &  _21 ) ;
 assign _233 = ( n_n101  &  _33 ) ;
 assign _235 = ( n_n103  &  _5301 ) ;
 assign _236 = ( n_n1185 ) | ( _445 ) ;
 assign _237 = ( n_n100  &  _5608 ) ;
 assign _238 = ( n_n1170 ) | ( n_n1173 ) ;
 assign _239 = ( n_n95  &  _4547 ) ;
 assign _240 = ( n_n67  &  _4461 ) ;
 assign _243 = ( n_n1125 ) | ( _825 ) ;
 assign _244 = ( n_n1075 ) | ( _1021 ) ;
 assign _245 = ( n_n1085 ) | ( _732 ) ;
 assign _246 = ( n_n76  &  _4963 ) ;
 assign _248 = ( n_n63  &  _38 ) ;
 assign _249 = ( n_n78  &  _42 ) ;
 assign _250 = ( n_n77  &  _30 ) ;
 assign _252 = ( n_n95  &  _42 ) ;
 assign _254 = ( _39  &  _5343 ) ;
 assign _255 = ( n_n981 ) | ( _792 ) ;
 assign _257 = ( n_n73  &  _27 ) ;
 assign _259 = ( n_n82  &  _27 ) ;
 assign _260 = ( n_n101  &  _41 ) ;
 assign _261 = ( n_n78  &  _44 ) ;
 assign _262 = ( n_n58  &  _19 ) ;
 assign _263 = ( n_n91  &  _19 ) ;
 assign _264 = ( n_n978 ) | ( n_n976 ) ;
 assign _265 = ( n_n101  &  _5234 ) ;
 assign _267 = ( n_n85  &  _5169 ) ;
 assign _268 = ( n_n58  &  _5022 ) ;
 assign _269 = ( n_n53  &  _5350 ) ;
 assign _270 = ( n_n66  &  _4541 ) ;
 assign _271 = ( n_n54  &  _4406 ) ;
 assign _272 = ( n_n58  &  _37 ) ;
 assign _273 = ( n_n103  &  _4887 ) ;
 assign _274 = ( n_n78  &  _22 ) ;
 assign _275 = ( n_n101  &  _25 ) ;
 assign _276 = ( n_n91  &  _42 ) ;
 assign _277 = ( n_n74  &  _20 ) ;
 assign _278 = ( n_n85  &  _5362 ) ;
 assign _279 = ( n_n53  &  _5023 ) ;
 assign _282 = ( n_n943 ) | ( _96 ) ;
 assign _283 = ( n_n85  &  _39 ) ;
 assign _284 = ( n_n91  &  _34 ) ;
 assign _286 = ( _67 ) | ( _839 ) ;
 assign _287 = ( _19  &  _5009 ) ;
 assign _288 = ( n_n95  &  _37 ) ;
 assign _289 = ( n_n74  &  _31 ) ;
 assign _290 = ( n_n91  &  _22 ) ;
 assign _291 = ( n_n99  &  _31 ) ;
 assign _293 = ( n_n93  &  _27 ) ;
 assign _295 = ( n_n87  &  _5145 ) ;
 assign _296 = ( (~ i_3_)  &  i_2_ ) ;
 assign _297 = ( i_5_  &  (~ i_3_) ) ;
 assign _298 = ( i_3_  &  i_0_ ) ;
 assign _299 = ( n_n94  &  n_n96 ) ;
 assign _300 = ( n_n97  &  n_n99 ) ;
 assign _301 = ( n_n81  &  n_n90 ) ;
 assign _302 = ( i_5_  &  i_3_ ) ;
 assign _303 = ( (~ i_5_)  &  (~ i_3_) ) ;
 assign _304 = ( i_1_  &  i_0_ ) ;
 assign _305 = ( i_1_  &  (~ i_0_) ) ;
 assign _306 = ( (~ i_1_)  &  (~ i_0_) ) ;
 assign _307 = ( n_n94  &  n_n84 ) ;
 assign _308 = ( n_n92  &  n_n90 ) ;
 assign _309 = ( n_n83  &  n_n82 ) ;
 assign _310 = ( n_n102  &  n_n103 ) ;
 assign _311 = ( n_n100  &  n_n74 ) ;
 assign _312 = ( n_n74  &  n_n103 ) ;
 assign _313 = ( i_5_  &  (~ i_4_) ) ;
 assign _314 = ( i_3_  &  i_4_ ) ;
 assign _315 = ( (~ i_3_)  &  (~ i_4_) ) ;
 assign _316 = ( n_n94  &  n_n92 ) ;
 assign _317 = ( n_n94  &  n_n81 ) ;
 assign _318 = ( n_n94  &  n_n74 ) ;
 assign _319 = ( n_n93  &  n_n83 ) ;
 assign _320 = ( n_n81  &  n_n100 ) ;
 assign _321 = ( n_n90  &  n_n96 ) ;
 assign _322 = ( n_n102  &  n_n85 ) ;
 assign _323 = ( n_n96  &  n_n103 ) ;
 assign _324 = ( n_n79  &  _4510 ) ;
 assign _325 = ( i_8_  &  (~ i_6_) ) ;
 assign _326 = ( (~ i_8_)  &  i_6_ ) ;
 assign _327 = ( (~ i_8_)  &  (~ i_6_) ) ;
 assign _328 = ( i_5_  &  i_4_ ) ;
 assign _329 = ( (~ i_5_)  &  (~ i_4_) ) ;
 assign _330 = ( (~ i_1_)  &  i_0_ ) ;
 assign _331 = ( n_n94  &  n_n99 ) ;
 assign _332 = ( n_n97  &  n_n77 ) ;
 assign _333 = ( n_n63  &  n_n83 ) ;
 assign _334 = ( n_n101  &  n_n83 ) ;
 assign _335 = ( n_n101  &  n_n85 ) ;
 assign _336 = ( n_n87  &  n_n64 ) ;
 assign _337 = ( n_n99  &  n_n103 ) ;
 assign _338 = ( (~ i_7_)  &  i_6_ ) ;
 assign _339 = ( n_n87  &  _5035 ) ;
 assign _340 = ( i_1_  &  (~ i_2_) ) ;
 assign _341 = ( n_n40  &  _4386 ) ;
 assign _342 = ( (~ i_1_)  &  _296 ) ;
 assign _343 = ( (~ i_2_)  &  _298 ) ;
 assign _344 = ( i_0_  &  _26 ) ;
 assign _345 = ( n_n71  &  _4964 ) ;
 assign _346 = ( n_n54  &  _4576 ) ;
 assign _347 = ( n_n94  &  n_n77 ) ;
 assign _348 = ( n_n78  &  n_n83 ) ;
 assign _349 = ( n_n92  &  n_n97 ) ;
 assign _350 = ( n_n95  &  n_n83 ) ;
 assign _351 = ( n_n95  &  n_n85 ) ;
 assign _352 = ( n_n82  &  n_n85 ) ;
 assign _353 = ( n_n84  &  n_n90 ) ;
 assign _354 = ( n_n96  &  n_n100 ) ;
 assign _355 = ( n_n67  &  n_n75 ) ;
 assign _356 = ( n_n40  &  n_n64 ) ;
 assign _357 = ( n_n99  &  n_n100 ) ;
 assign _358 = ( n_n85  &  n_n76 ) ;
 assign _359 = ( n_n85  &  n_n74 ) ;
 assign _360 = ( n_n79  &  n_n64 ) ;
 assign _361 = ( _43 ) | ( _299 ) ;
 assign _362 = ( _28 ) | ( _33 ) ;
 assign _363 = ( _24 ) | ( _300 ) ;
 assign _364 = ( _41 ) | ( _4412 ) ;
 assign _365 = ( _43 ) | ( _299 ) ;
 assign _366 = ( n_n81 ) | ( n_n99 ) ;
 assign _367 = ( n_n83 ) | ( n_n85 ) ;
 assign _368 = ( _28 ) | ( _33 ) ;
 assign _369 = ( _24 ) | ( _300 ) ;
 assign _370 = ( n_n81 ) | ( n_n99 ) ;
 assign _371 = ( _31 ) | ( _32 ) ;
 assign _372 = ( _722 ) | ( _723 ) ;
 assign _373 = ( _1017 ) | ( _1018 ) ;
 assign _374 = ( n_n101  &  _19 ) ;
 assign _381 = ( n_n92  &  _32 ) ;
 assign _382 = ( n_n58  &  _22 ) ;
 assign _387 = ( n_n81  &  _371 ) ;
 assign _388 = ( n_n101  &  _47 ) ;
 assign _389 = ( n_n78  &  _25 ) ;
 assign _392 = ( n_n101  &  _24 ) ;
 assign _398 = ( n_n70  &  _320 ) ;
 assign _399 = ( n_n81  &  _20 ) ;
 assign _404 = ( n_n82  &  _5634 ) ;
 assign _410 = ( n_n77  &  _5626 ) ;
 assign _411 = ( n_n86  &  _332 ) ;
 assign _416 = ( n_n101  &  _21 ) ;
 assign _422 = ( n_n103  &  _5615 ) ;
 assign _423 = ( n_n102  &  _319 ) ;
 assign _424 = ( n_n93  &  _312 ) ;
 assign _430 = ( n_n53  &  _360 ) ;
 assign _431 = ( n_n58  &  _22 ) ;
 assign _437 = ( n_n75  &  _25 ) ;
 assign _445 = ( n_n93  &  _25 ) ;
 assign _447 = ( n_n52  &  _29 ) ;
 assign _453 = ( n_n58  &  _5522 ) ;
 assign _454 = ( n_n85  &  _91 ) ;
 assign _461 = ( (~ i_5_)  &  _319 ) ;
 assign _468 = ( (~ i_3_)  &  _334 ) ;
 assign _475 = ( n_n64  &  _358 ) ;
 assign _476 = ( n_n52  &  _29 ) ;
 assign _481 = ( _47  &  _87 ) ;
 assign _482 = ( n_n63  &  _41 ) ;
 assign _489 = ( n_n93  &  _29 ) ;
 assign _497 = ( _39  &  _330 ) ;
 assign _501 = ( _35  &  _352 ) ;
 assign _502 = ( _297  &  _348 ) ;
 assign _507 = ( n_n74  &  _5439 ) ;
 assign _513 = ( _344  &  _5432 ) ;
 assign _520 = ( _36  &  _326 ) ;
 assign _522 = ( n_n83  &  _5398 ) ;
 assign _524 = ( n_n73  &  _322 ) ;
 assign _531 = ( n_n93  &  _5370 ) ;
 assign _537 = ( _20  &  _297 ) ;
 assign _538 = ( n_n58  &  _33 ) ;
 assign _543 = ( n_n93  &  _25 ) ;
 assign _549 = ( n_n101  &  _24 ) ;
 assign _556 = ( n_n58  &  _5344 ) ;
 assign _557 = ( _20  &  _370 ) ;
 assign _561 = ( n_n93  &  _29 ) ;
 assign _567 = ( n_n93  &  _311 ) ;
 assign _568 = ( n_n77  &  _309 ) ;
 assign _569 = ( n_n81  &  _31 ) ;
 assign _573 = ( n_n91  &  _47 ) ;
 assign _574 = ( n_n78  &  _38 ) ;
 assign _581 = ( n_n101  &  _19 ) ;
 assign _583 = ( n_n94  &  _5316 ) ;
 assign _590 = ( n_n101  &  _299 ) ;
 assign _596 = ( n_n101  &  _300 ) ;
 assign _604 = ( _35  &  _352 ) ;
 assign _610 = ( n_n70  &  _345 ) ;
 assign _611 = ( _41  &  _327 ) ;
 assign _616 = ( n_n86  &  _21 ) ;
 assign _617 = ( n_n99  &  _20 ) ;
 assign _624 = ( n_n70  &  _33 ) ;
 assign _632 = ( n_n85  &  _91 ) ;
 assign _634 = ( n_n74  &  n_n64 ) ;
 assign _635 = ( n_n86  &  n_n76 ) ;
 assign _636 = ( n_n91  &  _5239 ) ;
 assign _640 = ( n_n86  &  _332 ) ;
 assign _646 = ( n_n79  &  _5207 ) ;
 assign _652 = ( n_n58  &  _368 ) ;
 assign _658 = ( n_n77  &  _309 ) ;
 assign _659 = ( _40  &  _46 ) ;
 assign _660 = ( n_n81  &  _32 ) ;
 assign _664 = ( _25  &  _87 ) ;
 assign _671 = ( n_n58  &  _24 ) ;
 assign _675 = ( n_n81  &  _333 ) ;
 assign _676 = ( n_n70  &  _320 ) ;
 assign _681 = ( n_n64  &  _345 ) ;
 assign _687 = ( _36  &  _326 ) ;
 assign _693 = ( n_n103  &  _356 ) ;
 assign _696 = ( (~ i_3_)  &  _334 ) ;
 assign _702 = ( n_n86  &  _358 ) ;
 assign _709 = ( n_n40  &  _5095 ) ;
 assign _710 = ( _343  &  _5096 ) ;
 assign _717 = ( (~ i_5_)  &  _372 ) ;
 assign _722 = ( n_n101  &  _342 ) ;
 assign _723 = ( n_n90  &  n_n91 ) ;
 assign _724 = ( n_n85  &  _5084 ) ;
 assign _732 = ( n_n103  &  _5082 ) ;
 assign _734 = ( _297  &  _348 ) ;
 assign _740 = ( _41  &  _327 ) ;
 assign _741 = ( _29  &  _87 ) ;
 assign _747 = ( n_n58  &  _362 ) ;
 assign _748 = ( n_n101  &  _363 ) ;
 assign _749 = ( n_n64  &  _345 ) ;
 assign _753 = ( _20  &  _366 ) ;
 assign _758 = ( n_n92  &  _32 ) ;
 assign _759 = ( n_n93  &  _28 ) ;
 assign _765 = ( n_n102  &  _32 ) ;
 assign _766 = ( n_n58  &  _27 ) ;
 assign _767 = ( n_n93  &  _312 ) ;
 assign _768 = ( n_n91  &  _47 ) ;
 assign _769 = ( n_n97  &  _5037 ) ;
 assign _771 = ( n_n64  &  _359 ) ;
 assign _778 = ( n_n73  &  _322 ) ;
 assign _780 = ( i_8_  &  _341 ) ;
 assign _786 = ( n_n103  &  _356 ) ;
 assign _792 = ( n_n70  &  _33 ) ;
 assign _794 = ( n_n78  &  _38 ) ;
 assign _795 = ( n_n82  &  _28 ) ;
 assign _796 = ( n_n81  &  _333 ) ;
 assign _797 = ( _46  &  _325 ) ;
 assign _798 = ( n_n101  &  _365 ) ;
 assign _799 = ( n_n91  &  _300 ) ;
 assign _800 = ( n_n93  &  _28 ) ;
 assign _804 = ( n_n70  &  _345 ) ;
 assign _812 = ( n_n85  &  _4952 ) ;
 assign _818 = ( i_8_  &  _341 ) ;
 assign _825 = ( n_n73  &  _37 ) ;
 assign _827 = ( _4909  &  _4910 ) ;
 assign _833 = ( n_n95  &  _4894 ) ;
 assign _834 = ( _313  &  _355 ) ;
 assign _839 = ( n_n58  &  _28 ) ;
 assign _841 = ( n_n86  &  _45 ) ;
 assign _848 = ( _342  &  _4880 ) ;
 assign _850 = ( _40  &  _46 ) ;
 assign _852 = ( n_n81  &  _30 ) ;
 assign _854 = ( n_n101  &  _310 ) ;
 assign _856 = ( _40  &  _310 ) ;
 assign _864 = ( n_n82  &  _42 ) ;
 assign _865 = ( n_n63  &  _22 ) ;
 assign _870 = ( n_n93  &  _47 ) ;
 assign _876 = ( n_n79  &  _4761 ) ;
 assign _878 = ( n_n64  &  _358 ) ;
 assign _884 = ( n_n86  &  _341 ) ;
 assign _885 = ( n_n77  &  _20 ) ;
 assign _892 = ( n_n82  &  _42 ) ;
 assign _899 = ( n_n77  &  _20 ) ;
 assign _901 = ( _342  &  _4679 ) ;
 assign _903 = ( n_n82  &  _34 ) ;
 assign _911 = ( n_n85  &  _336 ) ;
 assign _913 = ( n_n52  &  _332 ) ;
 assign _915 = ( n_n73  &  _357 ) ;
 assign _917 = ( n_n63  &  _22 ) ;
 assign _923 = ( n_n63  &  _34 ) ;
 assign _925 = ( n_n101  &  _310 ) ;
 assign _927 = ( n_n93  &  _47 ) ;
 assign _935 = ( n_n86  &  _21 ) ;
 assign _943 = ( n_n73  &  _21 ) ;
 assign _951 = ( n_n101  &  _369 ) ;
 assign _952 = ( _20  &  _297 ) ;
 assign _953 = ( n_n86  &  _45 ) ;
 assign _958 = ( n_n85  &  _4540 ) ;
 assign _959 = ( n_n70  &  _42 ) ;
 assign _960 = ( n_n75  &  _25 ) ;
 assign _968 = ( n_n82  &  _34 ) ;
 assign _969 = ( n_n58  &  _24 ) ;
 assign _970 = ( _47  &  _325 ) ;
 assign _971 = ( n_n63  &  _28 ) ;
 assign _972 = ( n_n78  &  _25 ) ;
 assign _973 = ( n_n101  &  _21 ) ;
 assign _978 = ( n_n82  &  _28 ) ;
 assign _986 = ( _40  &  _353 ) ;
 assign _987 = ( n_n75  &  _299 ) ;
 assign _988 = ( i_1_  &  _324 ) ;
 assign _990 = ( n_n80  &  _4504 ) ;
 assign _991 = ( n_n100  &  _4505 ) ;
 assign _996 = ( n_n77  &  _4494 ) ;
 assign _1004 = ( n_n73  &  _37 ) ;
 assign _1010 = ( _304  &  _373 ) ;
 assign _1017 = ( n_n95  &  _302 ) ;
 assign _1018 = ( n_n81  &  n_n86 ) ;
 assign _1019 = ( n_n73  &  _21 ) ;
 assign _1021 = ( _40  &  _310 ) ;
 assign _1023 = ( (~ i_5_)  &  _319 ) ;
 assign _1030 = ( n_n85  &  _4453 ) ;
 assign _1032 = ( n_n58  &  _4446 ) ;
 assign _1034 = ( n_n78  &  _4444 ) ;
 assign _1035 = ( n_n40  &  _4445 ) ;
 assign _1036 = ( n_n91  &  _4422 ) ;
 assign _1037 = ( n_n101  &  _361 ) ;
 assign _1041 = ( _367  &  _4417 ) ;
 assign _1042 = ( n_n58  &  _27 ) ;
 assign _1046 = ( n_n100  &  _4411 ) ;
 assign _1047 = ( n_n63  &  _364 ) ;
 assign _1048 = ( n_n93  &  _311 ) ;
 assign _1049 = ( n_n91  &  _300 ) ;
 assign _1052 = ( n_n95  &  _312 ) ;
 assign _1053 = ( n_n81  &  _30 ) ;
 assign _1054 = ( n_n73  &  _332 ) ;
 assign _1056 = ( n_n86  &  _341 ) ;
 assign _1057 = ( n_n102  &  _32 ) ;
 assign _4385 = ( (~ i_6_)  &  (~ i_5_) ) ;
 assign _4386 = ( _298  &  (~ i_1_) ) ;
 assign _4387 = ( _81 ) | ( n_n1281 ) ;
 assign _4388 = ( _119 ) | ( _117 ) ;
 assign _4389 = ( _1057 ) | ( _1056 ) ;
 assign _4390 = ( _4388 ) | ( _4387 ) ;
 assign _4391 = ( n_n1267 ) | ( n_n1217 ) ;
 assign _4392 = ( _182 ) | ( n_n1174 ) ;
 assign _4393 = ( _275 ) | ( _194 ) ;
 assign _4394 = ( _65 ) | ( _293 ) ;
 assign _4395 = ( _4392 ) | ( _4391 ) ;
 assign _4396 = ( _4394 ) | ( _4393 ) ;
 assign _4397 = ( n_n83  &  n_n73 ) ;
 assign _4398 = ( n_n1134 ) | ( n_n1164 ) ;
 assign _4399 = ( n_n1156 ) | ( n_n1091 ) ;
 assign _4400 = ( _128 ) | ( n_n1120 ) ;
 assign _4401 = ( _4399 ) | ( _4398 ) ;
 assign _4402 = ( n_n54  &  n_n70 ) ;
 assign _4403 = ( n_n1021 ) | ( n_n956 ) ;
 assign _4404 = ( _4403 ) | ( _76 ) ;
 assign _4405 = ( (~ i_2_)  &  (~ i_3_) ) ;
 assign _4406 = ( n_n80  &  n_n75 ) ;
 assign _4407 = ( _151 ) | ( _55 ) ;
 assign _4408 = ( _4407 ) | ( _271 ) ;
 assign _4409 = ( wire4181 ) | ( _4408 ) ;
 assign _4410 = ( n_n110 ) | ( n_n109 ) ;
 assign _4411 = ( n_n82  &  _314 ) ;
 assign _4412 = ( _34 ) | ( _28 ) ;
 assign _4413 = ( _1046 ) | ( _208 ) ;
 assign _4414 = ( _1049 ) | ( _1048 ) ;
 assign _4415 = ( _4413 ) | ( _94 ) ;
 assign _4416 = ( _1047 ) | ( _4414 ) ;
 assign _4417 = ( n_n81  &  n_n52 ) ;
 assign _4418 = ( _260 ) | ( _177 ) ;
 assign _4419 = ( _1041 ) | ( _261 ) ;
 assign _4420 = ( _4418 ) | ( _1042 ) ;
 assign _4421 = ( i_2_  &  (~ i_1_) ) ;
 assign _4422 = ( n_n81  &  _4421 ) ;
 assign _4423 = ( _1037 ) | ( _1036 ) ;
 assign _4424 = ( wire4164 ) | ( _4423 ) ;
 assign _4425 = ( _4424 ) | ( n_n106 ) ;
 assign _4426 = ( n_n943 ) | ( n_n951 ) ;
 assign _4427 = ( n_n952 ) | ( n_n957 ) ;
 assign _4428 = ( n_n940 ) | ( n_n950 ) ;
 assign _4429 = ( _210 ) | ( n_n959 ) ;
 assign _4430 = ( _4427 ) | ( _4426 ) ;
 assign _4431 = ( _4429 ) | ( _4428 ) ;
 assign _4432 = ( n_n95  &  _297 ) ;
 assign _4433 = ( n_n70  &  (~ i_3_) ) ;
 assign _4434 = ( n_n71  &  _305 ) ;
 assign _4435 = ( i_1_  &  (~ i_4_) ) ;
 assign _4436 = ( _4435  &  _298 ) ;
 assign _4437 = ( n_n1011 ) | ( _129 ) ;
 assign _4438 = ( n_n1025 ) | ( n_n1022 ) ;
 assign _4439 = ( _68 ) | ( n_n1026 ) ;
 assign _4440 = ( _219 ) | ( _184 ) ;
 assign _4441 = ( _4438 ) | ( _4437 ) ;
 assign _4442 = ( _4440 ) | ( _4439 ) ;
 assign _4443 = ( n_n71  &  n_n86 ) ;
 assign _4444 = ( _340  &  _303 ) ;
 assign _4445 = ( n_n80  &  (~ i_8_) ) ;
 assign _4446 = ( n_n83  &  (~ i_3_) ) ;
 assign _4447 = ( n_n1054 ) | ( n_n1068 ) ;
 assign _4448 = ( n_n1059 ) | ( n_n1052 ) ;
 assign _4449 = ( _49 ) | ( _143 ) ;
 assign _4450 = ( _4447 ) | ( _152 ) ;
 assign _4451 = ( _4449 ) | ( _4448 ) ;
 assign _4452 = ( i_0_  &  i_2_ ) ;
 assign _4453 = ( _40  &  _35 ) ;
 assign _4454 = ( n_n1043 ) | ( n_n1046 ) ;
 assign _4455 = ( _195 ) | ( n_n1042 ) ;
 assign _4456 = ( _145 ) | ( _1023 ) ;
 assign _4457 = ( _4454 ) | ( _200 ) ;
 assign _4458 = ( _4456 ) | ( _4455 ) ;
 assign _4459 = ( n_n142 ) | ( n_n144 ) ;
 assign _4460 = ( n_n83  &  n_n75 ) ;
 assign _4461 = ( n_n93  &  (~ i_4_) ) ;
 assign _4462 = ( n_n83  &  _40 ) ;
 assign _4463 = ( n_n1078 ) | ( n_n1077 ) ;
 assign _4464 = ( n_n1079 ) | ( n_n1081 ) ;
 assign _4465 = ( _69 ) | ( n_n1070 ) ;
 assign _4466 = ( _244 ) | ( _240 ) ;
 assign _4467 = ( _4464 ) | ( _4463 ) ;
 assign _4468 = ( _4466 ) | ( _4465 ) ;
 assign _4469 = ( _111 ) | ( n_n1092 ) ;
 assign _4470 = ( _147 ) | ( _115 ) ;
 assign _4471 = ( _102 ) | ( _257 ) ;
 assign _4472 = ( _4469 ) | ( _1010 ) ;
 assign _4473 = ( _4471 ) | ( _4470 ) ;
 assign _4474 = ( i_3_  &  (~ i_5_) ) ;
 assign _4475 = ( n_n83  &  n_n64 ) ;
 assign _4476 = ( n_n1117 ) | ( n_n1130 ) ;
 assign _4477 = ( _114 ) | ( n_n1108 ) ;
 assign _4478 = ( _1004 ) | ( _190 ) ;
 assign _4479 = ( _4477 ) | ( _4476 ) ;
 assign _4480 = ( n_n1105 ) | ( n_n1100 ) ;
 assign _4481 = ( _4480 ) | ( n_n1103 ) ;
 assign _4482 = ( wire4296 ) | ( _4481 ) ;
 assign _4483 = ( n_n140 ) | ( n_n141 ) ;
 assign _4484 = ( _4483 ) | ( _4482 ) ;
 assign _4485 = ( _64 ) | ( n_n995 ) ;
 assign _4486 = ( n_n97  &  (~ i_7_) ) ;
 assign _4487 = ( n_n991 ) | ( n_n1004 ) ;
 assign _4488 = ( n_n1006 ) | ( n_n986 ) ;
 assign _4489 = ( _220 ) | ( n_n989 ) ;
 assign _4490 = ( _4488 ) | ( _4487 ) ;
 assign _4491 = ( n_n882 ) | ( _4489 ) ;
 assign _4492 = ( n_n71  &  n_n70 ) ;
 assign _4493 = ( i_2_  &  i_7_ ) ;
 assign _4494 = ( _4493  &  i_0_ ) ;
 assign _4495 = ( n_n975 ) | ( _996 ) ;
 assign _4496 = ( n_n968 ) | ( n_n967 ) ;
 assign _4497 = ( n_n984 ) | ( n_n973 ) ;
 assign _4498 = ( _264 ) | ( n_n982 ) ;
 assign _4499 = ( _4496 ) | ( _4495 ) ;
 assign _4500 = ( _4498 ) | ( _4497 ) ;
 assign _4501 = ( n_n145 ) | ( n_n147 ) ;
 assign _4502 = ( _4501 ) | ( n_n146 ) ;
 assign _4503 = ( _26  &  i_1_ ) ;
 assign _4504 = ( _313  &  n_n86 ) ;
 assign _4505 = ( n_n78  &  i_5_ ) ;
 assign _4506 = ( n_n1172 ) | ( _990 ) ;
 assign _4507 = ( _162 ) | ( n_n1153 ) ;
 assign _4508 = ( _991 ) | ( _163 ) ;
 assign _4509 = ( _4507 ) | ( _4506 ) ;
 assign _4510 = ( _26  &  n_n75 ) ;
 assign _4511 = ( n_n1204 ) | ( n_n1181 ) ;
 assign _4512 = ( _67 ) | ( _66 ) ;
 assign _4513 = ( _185 ) | ( _142 ) ;
 assign _4514 = ( _90 ) | ( _186 ) ;
 assign _4515 = ( _4512 ) | ( _4511 ) ;
 assign _4516 = ( _4514 ) | ( _4513 ) ;
 assign _4517 = ( n_n1279 ) | ( n_n1324 ) ;
 assign _4518 = ( _79 ) | ( n_n1297 ) ;
 assign _4519 = ( _289 ) | ( _171 ) ;
 assign _4520 = ( _88 ) | ( _978 ) ;
 assign _4521 = ( _4518 ) | ( _4517 ) ;
 assign _4522 = ( _4520 ) | ( _4519 ) ;
 assign _4523 = ( _93 ) | ( n_n1330 ) ;
 assign _4524 = ( _259 ) | ( _131 ) ;
 assign _4525 = ( _971 ) | ( _970 ) ;
 assign _4526 = ( _973 ) | ( _972 ) ;
 assign _4527 = ( _4524 ) | ( _4523 ) ;
 assign _4528 = ( _4526 ) | ( _4525 ) ;
 assign _4529 = ( n_n93  &  _305 ) ;
 assign _4530 = ( i_3_  &  (~ i_5_) ) ;
 assign _4531 = ( n_n63  &  _314 ) ;
 assign _4532 = ( _304  &  (~ i_3_) ) ;
 assign _4533 = ( _169 ) | ( _137 ) ;
 assign _4534 = ( _172 ) | ( _170 ) ;
 assign _4535 = ( _276 ) | ( _187 ) ;
 assign _4536 = ( _70 ) | ( _960 ) ;
 assign _4537 = ( _4534 ) | ( _4533 ) ;
 assign _4538 = ( _4536 ) | ( _4535 ) ;
 assign _4539 = ( n_n134 ) | ( n_n133 ) ;
 assign _4540 = ( n_n87  &  n_n75 ) ;
 assign _4541 = ( n_n83  &  n_n75 ) ;
 assign _4542 = ( _140 ) | ( n_n1215 ) ;
 assign _4543 = ( _952 ) | ( _270 ) ;
 assign _4544 = ( _104 ) | ( _953 ) ;
 assign _4545 = ( _4542 ) | ( _951 ) ;
 assign _4546 = ( _4544 ) | ( _4543 ) ;
 assign _4547 = ( n_n97  &  _35 ) ;
 assign _4548 = ( _164 ) | ( _149 ) ;
 assign _4549 = ( _4548 ) | ( _239 ) ;
 assign _4550 = ( wire4411 ) | ( _4549 ) ;
 assign _4551 = ( n_n136 ) | ( n_n137 ) ;
 assign _4552 = ( _4551 ) | ( _4550 ) ;
 assign _4553 = ( _4552 ) | ( n_n128 ) ;
 assign _4554 = ( n_n90  &  i_6_ ) ;
 assign _4555 = ( n_n969 ) | ( n_n956 ) ;
 assign _4556 = ( n_n978 ) | ( n_n955 ) ;
 assign _4557 = ( _99 ) | ( n_n961 ) ;
 assign _4558 = ( _4555 ) | ( _215 ) ;
 assign _4559 = ( _4557 ) | ( _4556 ) ;
 assign _4560 = ( n_n991 ) | ( n_n1004 ) ;
 assign _4561 = ( n_n1014 ) | ( n_n981 ) ;
 assign _4562 = ( _181 ) | ( _64 ) ;
 assign _4563 = ( _144 ) | ( _184 ) ;
 assign _4564 = ( _4561 ) | ( _4560 ) ;
 assign _4565 = ( _4563 ) | ( _4562 ) ;
 assign _4566 = ( n_n1164 ) | ( n_n1181 ) ;
 assign _4567 = ( n_n1172 ) | ( n_n1146 ) ;
 assign _4568 = ( _134 ) | ( n_n1158 ) ;
 assign _4569 = ( _218 ) | ( _135 ) ;
 assign _4570 = ( _4567 ) | ( _4566 ) ;
 assign _4571 = ( _4569 ) | ( _4568 ) ;
 assign _4572 = ( n_n1095 ) | ( n_n1132 ) ;
 assign _4573 = ( n_n1128 ) | ( n_n1134 ) ;
 assign _4574 = ( _161 ) | ( n_n1130 ) ;
 assign _4575 = ( _4573 ) | ( _4572 ) ;
 assign _4576 = ( _296  &  (~ i_0_) ) ;
 assign _4577 = ( n_n1055 ) | ( n_n1060 ) ;
 assign _4578 = ( n_n1032 ) | ( n_n1022 ) ;
 assign _4579 = ( n_n1036 ) | ( n_n1039 ) ;
 assign _4580 = ( _217 ) | ( _943 ) ;
 assign _4581 = ( _4578 ) | ( _4577 ) ;
 assign _4582 = ( _4580 ) | ( _4579 ) ;
 assign _4583 = ( n_n1204 ) | ( n_n1217 ) ;
 assign _4584 = ( n_n1188 ) | ( n_n1193 ) ;
 assign _4585 = ( _185 ) | ( _160 ) ;
 assign _4586 = ( _65 ) | ( _290 ) ;
 assign _4587 = ( _4584 ) | ( _4583 ) ;
 assign _4588 = ( _4586 ) | ( _4585 ) ;
 assign _4589 = ( n_n1259 ) | ( n_n1254 ) ;
 assign _4590 = ( _140 ) | ( _73 ) ;
 assign _4591 = ( _188 ) | ( _187 ) ;
 assign _4592 = ( _70 ) | ( _935 ) ;
 assign _4593 = ( _4590 ) | ( _4589 ) ;
 assign _4594 = ( _4592 ) | ( _4591 ) ;
 assign _4595 = ( _110 ) | ( _83 ) ;
 assign _4596 = ( _232 ) | ( _159 ) ;
 assign _4597 = ( _259 ) | ( _252 ) ;
 assign _4598 = ( _133 ) | ( _927 ) ;
 assign _4599 = ( _4596 ) | ( _4595 ) ;
 assign _4600 = ( _4598 ) | ( _4597 ) ;
 assign _4601 = ( n_n769 ) | ( n_n770 ) ;
 assign _4602 = ( n_n1085 ) | ( n_n1088 ) ;
 assign _4603 = ( _4602 ) | ( n_n1093 ) ;
 assign _4604 = ( wire4462 ) | ( _4603 ) ;
 assign _4605 = ( n_n773 ) | ( n_n771 ) ;
 assign _4606 = ( _4605 ) | ( _4604 ) ;
 assign _4607 = ( _306  &  (~ i_6_) ) ;
 assign _4608 = ( n_n946 ) | ( n_n937 ) ;
 assign _4609 = ( n_n950 ) | ( n_n943 ) ;
 assign _4610 = ( _4608 ) | ( n_n942 ) ;
 assign _4611 = ( _214 ) | ( _207 ) ;
 assign _4612 = ( _4610 ) | ( _4609 ) ;
 assign _4613 = ( _306  &  _303 ) ;
 assign _4614 = ( _203 ) | ( _917 ) ;
 assign _4615 = ( n_n776 ) | ( _4614 ) ;
 assign _4616 = ( n_n774 ) | ( n_n775 ) ;
 assign _4617 = ( _4616 ) | ( _4615 ) ;
 assign _4618 = ( n_n1134 ) | ( n_n1092 ) ;
 assign _4619 = ( n_n1103 ) | ( n_n1093 ) ;
 assign _4620 = ( _103 ) | ( n_n1120 ) ;
 assign _4621 = ( _4619 ) | ( _4618 ) ;
 assign _4622 = ( n_n874 ) | ( _4620 ) ;
 assign _4623 = ( n_n94  &  _314 ) ;
 assign _4624 = ( n_n1032 ) | ( n_n1022 ) ;
 assign _4625 = ( n_n1039 ) | ( n_n1040 ) ;
 assign _4626 = ( _145 ) | ( n_n1052 ) ;
 assign _4627 = ( _4624 ) | ( _213 ) ;
 assign _4628 = ( _4626 ) | ( _4625 ) ;
 assign _4629 = ( n_n81  &  _325 ) ;
 assign _4630 = ( _161 ) | ( _135 ) ;
 assign _4631 = ( n_n1164 ) | ( n_n1184 ) ;
 assign _4632 = ( n_n1172 ) | ( n_n1146 ) ;
 assign _4633 = ( n_n1170 ) | ( n_n1153 ) ;
 assign _4634 = ( _4632 ) | ( _4631 ) ;
 assign _4635 = ( _169 ) | ( _159 ) ;
 assign _4636 = ( _183 ) | ( _170 ) ;
 assign _4637 = ( _284 ) | ( _233 ) ;
 assign _4638 = ( _189 ) | ( _903 ) ;
 assign _4639 = ( _4636 ) | ( _4635 ) ;
 assign _4640 = ( _4638 ) | ( _4637 ) ;
 assign _4641 = ( n_n1217 ) | ( n_n1216 ) ;
 assign _4642 = ( _140 ) | ( _123 ) ;
 assign _4643 = ( _188 ) | ( _185 ) ;
 assign _4644 = ( _65 ) | ( _290 ) ;
 assign _4645 = ( _4642 ) | ( _4641 ) ;
 assign _4646 = ( _4644 ) | ( _4643 ) ;
 assign _4647 = ( wire4570 ) | ( n_n554 ) ;
 assign _4648 = ( n_n728 ) | ( n_n727 ) ;
 assign _4649 = ( n_n1091 ) | ( n_n1085 ) ;
 assign _4650 = ( n_n1075 ) | ( n_n1078 ) ;
 assign _4651 = ( _168 ) | ( _69 ) ;
 assign _4652 = ( _4650 ) | ( _4649 ) ;
 assign _4653 = ( n_n1058 ) | ( n_n1055 ) ;
 assign _4654 = ( _4653 ) | ( n_n1054 ) ;
 assign _4655 = ( wire4556 ) | ( _4654 ) ;
 assign _4656 = ( n_n732 ) | ( n_n730 ) ;
 assign _4657 = ( _4656 ) | ( _4655 ) ;
 assign _4658 = ( n_n946 ) | ( n_n937 ) ;
 assign _4659 = ( n_n943 ) | ( n_n951 ) ;
 assign _4660 = ( n_n940 ) | ( n_n939 ) ;
 assign _4661 = ( _4658 ) | ( n_n941 ) ;
 assign _4662 = ( _4659 ) | ( _97 ) ;
 assign _4663 = ( _4661 ) | ( _4660 ) ;
 assign _4664 = ( n_n78  &  _315 ) ;
 assign _4665 = ( n_n981 ) | ( n_n957 ) ;
 assign _4666 = ( n_n971 ) | ( n_n955 ) ;
 assign _4667 = ( n_n984 ) | ( n_n983 ) ;
 assign _4668 = ( _264 ) | ( n_n959 ) ;
 assign _4669 = ( _4666 ) | ( _4665 ) ;
 assign _4670 = ( _4668 ) | ( _4667 ) ;
 assign _4671 = ( n_n991 ) | ( n_n999 ) ;
 assign _4672 = ( n_n1001 ) | ( n_n1018 ) ;
 assign _4673 = ( n_n1014 ) | ( n_n1010 ) ;
 assign _4674 = ( _211 ) | ( _184 ) ;
 assign _4675 = ( _4672 ) | ( _4671 ) ;
 assign _4676 = ( _4674 ) | ( _4673 ) ;
 assign _4677 = ( n_n734 ) | ( n_n735 ) ;
 assign _4678 = ( _4677 ) | ( n_n733 ) ;
 assign _4679 = ( n_n66  &  n_n86 ) ;
 assign _4680 = ( n_n1331 ) | ( n_n1324 ) ;
 assign _4681 = ( _177 ) | ( _55 ) ;
 assign _4682 = ( _54 ) | ( _263 ) ;
 assign _4683 = ( _4680 ) | ( _176 ) ;
 assign _4684 = ( _4682 ) | ( _4681 ) ;
 assign _4685 = ( _122 ) | ( _93 ) ;
 assign _4686 = ( _272 ) | ( _262 ) ;
 assign _4687 = ( _4685 ) | ( _892 ) ;
 assign _4688 = ( _4687 ) | ( _4686 ) ;
 assign _4689 = ( n_n726 ) | ( _4688 ) ;
 assign _4690 = ( _81 ) | ( _55 ) ;
 assign _4691 = ( _83 ) | ( _82 ) ;
 assign _4692 = ( _884 ) | ( _157 ) ;
 assign _4693 = ( _54 ) | ( _885 ) ;
 assign _4694 = ( _4691 ) | ( _4690 ) ;
 assign _4695 = ( _4693 ) | ( _4692 ) ;
 assign _4696 = ( _79 ) | ( n_n1259 ) ;
 assign _4697 = ( _171 ) | ( _158 ) ;
 assign _4698 = ( _223 ) | ( _183 ) ;
 assign _4699 = ( _189 ) | ( _233 ) ;
 assign _4700 = ( _4697 ) | ( _4696 ) ;
 assign _4701 = ( _4699 ) | ( _4698 ) ;
 assign _4702 = ( _296  &  i_0_ ) ;
 assign _4703 = ( n_n1215 ) | ( n_n1193 ) ;
 assign _4704 = ( _201 ) | ( _123 ) ;
 assign _4705 = ( _878 ) | ( _216 ) ;
 assign _4706 = ( _4704 ) | ( _4703 ) ;
 assign _4707 = ( n_n980 ) | ( n_n969 ) ;
 assign _4708 = ( n_n966 ) | ( n_n971 ) ;
 assign _4709 = ( n_n976 ) | ( n_n961 ) ;
 assign _4710 = ( _4708 ) | ( _4707 ) ;
 assign _4711 = ( n_n989 ) | ( n_n986 ) ;
 assign _4712 = ( _4711 ) | ( n_n983 ) ;
 assign _4713 = ( _306  &  (~ i_3_) ) ;
 assign _4714 = ( n_n1001 ) | ( _53 ) ;
 assign _4715 = ( n_n1030 ) | ( n_n1010 ) ;
 assign _4716 = ( _4714 ) | ( _213 ) ;
 assign _4717 = ( n_n882 ) | ( _4715 ) ;
 assign _4718 = ( n_n958 ) | ( n_n957 ) ;
 assign _4719 = ( n_n939 ) | ( n_n937 ) ;
 assign _4720 = ( n_n949 ) | ( n_n944 ) ;
 assign _4721 = ( _4719 ) | ( _97 ) ;
 assign _4722 = ( n_n716 ) | ( _4720 ) ;
 assign _4723 = ( _4722 ) | ( _4721 ) ;
 assign _4724 = ( n_n855 ) | ( n_n856 ) ;
 assign _4725 = ( n_n1082 ) | ( n_n1092 ) ;
 assign _4726 = ( n_n1078 ) | ( n_n1095 ) ;
 assign _4727 = ( n_n1103 ) | ( n_n1079 ) ;
 assign _4728 = ( _4726 ) | ( _4725 ) ;
 assign _4729 = ( n_n874 ) | ( _4727 ) ;
 assign _4730 = ( n_n1177 ) | ( n_n1153 ) ;
 assign _4731 = ( n_n1120 ) | ( n_n1158 ) ;
 assign _4732 = ( _63 ) | ( n_n1174 ) ;
 assign _4733 = ( _238 ) | ( _167 ) ;
 assign _4734 = ( _4731 ) | ( _4730 ) ;
 assign _4735 = ( _4733 ) | ( _4732 ) ;
 assign _4736 = ( n_n1035 ) | ( n_n1058 ) ;
 assign _4737 = ( n_n1054 ) | ( n_n1070 ) ;
 assign _4738 = ( _69 ) | ( n_n1052 ) ;
 assign _4739 = ( _244 ) | ( _168 ) ;
 assign _4740 = ( _4737 ) | ( _4736 ) ;
 assign _4741 = ( _4739 ) | ( _4738 ) ;
 assign _4742 = ( n_n852 ) | ( n_n853 ) ;
 assign _4743 = ( _4742 ) | ( n_n854 ) ;
 assign _4744 = ( _306  &  n_n86 ) ;
 assign _4745 = ( _74 ) | ( _166 ) ;
 assign _4746 = ( _4745 ) | ( _169 ) ;
 assign _4747 = ( wire4662 ) | ( _4746 ) ;
 assign _4748 = ( n_n850 ) | ( n_n849 ) ;
 assign _4749 = ( _4748 ) | ( _4747 ) ;
 assign _4750 = ( _121 ) | ( n_n1330 ) ;
 assign _4751 = ( _250 ) | ( _122 ) ;
 assign _4752 = ( _262 ) | ( _261 ) ;
 assign _4753 = ( _4751 ) | ( _4750 ) ;
 assign _4754 = ( _125 ) | ( n_n1324 ) ;
 assign _4755 = ( _263 ) | ( _177 ) ;
 assign _4756 = ( _203 ) | ( _272 ) ;
 assign _4757 = ( _4755 ) | ( _4754 ) ;
 assign _4758 = ( _4757 ) | ( _4756 ) ;
 assign _4759 = ( _4758 ) | ( wire4670 ) ;
 assign _4760 = ( n_n40  &  n_n86 ) ;
 assign _4761 = ( n_n83  &  n_n86 ) ;
 assign _4762 = ( _72 ) | ( n_n1254 ) ;
 assign _4763 = ( _171 ) | ( _100 ) ;
 assign _4764 = ( _116 ) | ( _223 ) ;
 assign _4765 = ( _4762 ) | ( _133 ) ;
 assign _4766 = ( _4764 ) | ( _4763 ) ;
 assign _4767 = ( _81 ) | ( _79 ) ;
 assign _4768 = ( _157 ) | ( _82 ) ;
 assign _4769 = ( _291 ) | ( _158 ) ;
 assign _4770 = ( _4768 ) | ( _4767 ) ;
 assign _4771 = ( n_n1330 ) | ( n_n1331 ) ;
 assign _4772 = ( _4771 ) | ( _252 ) ;
 assign _4773 = ( _121 ) | ( _93 ) ;
 assign _4774 = ( _259 ) | ( _250 ) ;
 assign _4775 = ( _870 ) | ( _261 ) ;
 assign _4776 = ( _4774 ) | ( _4773 ) ;
 assign _4777 = ( _864 ) | ( _125 ) ;
 assign _4778 = ( _4777 ) | ( _865 ) ;
 assign _4779 = ( wire4694 ) | ( _4778 ) ;
 assign _4780 = ( n_n808 ) | ( n_n809 ) ;
 assign _4781 = ( n_n1128 ) | ( n_n1088 ) ;
 assign _4782 = ( n_n1070 ) | ( n_n1079 ) ;
 assign _4783 = ( _71 ) | ( n_n1130 ) ;
 assign _4784 = ( _102 ) | ( _856 ) ;
 assign _4785 = ( _4782 ) | ( _4781 ) ;
 assign _4786 = ( _4784 ) | ( _4783 ) ;
 assign _4787 = ( n_n1163 ) | ( n_n1181 ) ;
 assign _4788 = ( n_n1173 ) | ( n_n1177 ) ;
 assign _4789 = ( _63 ) | ( n_n1174 ) ;
 assign _4790 = ( _4788 ) | ( _4787 ) ;
 assign _4791 = ( n_n1160 ) | ( n_n1132 ) ;
 assign _4792 = ( _4791 ) | ( _134 ) ;
 assign _4793 = ( n_n1204 ) | ( n_n1216 ) ;
 assign _4794 = ( _73 ) | ( n_n1215 ) ;
 assign _4795 = ( _160 ) | ( _74 ) ;
 assign _4796 = ( _4794 ) | ( _4793 ) ;
 assign _4797 = ( n_n1188 ) | ( n_n1184 ) ;
 assign _4798 = ( _4797 ) | ( _216 ) ;
 assign _4799 = ( wire4685 ) | ( _4798 ) ;
 assign _4800 = ( n_n811 ) | ( n_n812 ) ;
 assign _4801 = ( _4800 ) | ( _4799 ) ;
 assign _4802 = ( n_n986 ) | ( n_n987 ) ;
 assign _4803 = ( n_n966 ) | ( n_n980 ) ;
 assign _4804 = ( _215 ) | ( _99 ) ;
 assign _4805 = ( n_n504 ) | ( _4803 ) ;
 assign _4806 = ( n_n950 ) | ( n_n937 ) ;
 assign _4807 = ( n_n944 ) | ( n_n955 ) ;
 assign _4808 = ( _221 ) | ( n_n942 ) ;
 assign _4809 = ( _4806 ) | ( _222 ) ;
 assign _4810 = ( _4808 ) | ( _4807 ) ;
 assign _4811 = ( n_n999 ) | ( _53 ) ;
 assign _4812 = ( n_n995 ) | ( n_n1004 ) ;
 assign _4813 = ( n_n1021 ) | ( n_n1030 ) ;
 assign _4814 = ( _4812 ) | ( _4811 ) ;
 assign _4815 = ( n_n1042 ) | ( n_n1060 ) ;
 assign _4816 = ( _4815 ) | ( _283 ) ;
 assign _4817 = ( wire4715 ) | ( _4816 ) ;
 assign _4818 = ( n_n815 ) | ( n_n814 ) ;
 assign _4819 = ( _4818 ) | ( _4817 ) ;
 assign _4820 = ( n_n1254 ) | ( n_n1176 ) ;
 assign _4821 = ( n_n1074 ) | ( n_n1132 ) ;
 assign _4822 = ( n_n1032 ) | ( n_n1109 ) ;
 assign _4823 = ( _206 ) | ( n_n955 ) ;
 assign _4824 = ( _4821 ) | ( _4820 ) ;
 assign _4825 = ( _4823 ) | ( _4822 ) ;
 assign _4826 = ( _130 ) | ( n_n1369 ) ;
 assign _4827 = ( n_n1331 ) | ( n_n1283 ) ;
 assign _4828 = ( n_n1297 ) | ( n_n1294 ) ;
 assign _4829 = ( _133 ) | ( _48 ) ;
 assign _4830 = ( _4827 ) | ( _204 ) ;
 assign _4831 = ( _4829 ) | ( _4828 ) ;
 assign _4832 = ( _4831 ) | ( _4830 ) ;
 assign _4833 = ( n_n1331 ) | ( n_n1369 ) ;
 assign _4834 = ( _50 ) | ( n_n1330 ) ;
 assign _4835 = ( _131 ) | ( _95 ) ;
 assign _4836 = ( _4834 ) | ( _4833 ) ;
 assign _4837 = ( n_n1259 ) | ( n_n1254 ) ;
 assign _4838 = ( n_n1057 ) | ( n_n1109 ) ;
 assign _4839 = ( _51 ) | ( n_n1125 ) ;
 assign _4840 = ( _4838 ) | ( _4837 ) ;
 assign _4841 = ( n_n1283 ) | ( n_n1324 ) ;
 assign _4842 = ( n_n1286 ) | ( n_n1297 ) ;
 assign _4843 = ( _133 ) | ( _48 ) ;
 assign _4844 = ( _4841 ) | ( _204 ) ;
 assign _4845 = ( _4843 ) | ( _4842 ) ;
 assign _4846 = ( n_n1032 ) | ( n_n1042 ) ;
 assign _4847 = ( n_n1039 ) | ( n_n955 ) ;
 assign _4848 = ( _206 ) | ( n_n942 ) ;
 assign _4849 = ( _4846 ) | ( _227 ) ;
 assign _4850 = ( _4848 ) | ( _4847 ) ;
 assign _4851 = ( n_n1169 ) | ( n_n1132 ) ;
 assign _4852 = ( _4851 ) | ( n_n1128 ) ;
 assign _4853 = ( n_n889 ) | ( _4852 ) ;
 assign _4854 = ( n_n892 ) | ( wire4743 ) ;
 assign _4855 = ( _4853 ) | ( n_n890 ) ;
 assign _4856 = ( n_n1169 ) | ( n_n1074 ) ;
 assign _4857 = ( n_n1128 ) | ( n_n1109 ) ;
 assign _4858 = ( _51 ) | ( n_n1125 ) ;
 assign _4859 = ( _4857 ) | ( _4856 ) ;
 assign _4860 = ( n_n1294 ) | ( _166 ) ;
 assign _4861 = ( _4860 ) | ( n_n1286 ) ;
 assign _4862 = ( n_n1330 ) | ( n_n1324 ) ;
 assign _4863 = ( _131 ) | ( _95 ) ;
 assign _4864 = ( _4862 ) | ( _208 ) ;
 assign _4865 = ( _4864 ) | ( _4863 ) ;
 assign _4866 = ( _53 ) | ( n_n937 ) ;
 assign _4867 = ( n_n1039 ) | ( n_n1042 ) ;
 assign _4868 = ( _4866 ) | ( n_n1057 ) ;
 assign _4869 = ( _227 ) | ( _96 ) ;
 assign _4870 = ( _4868 ) | ( _4867 ) ;
 assign _4871 = ( _4870 ) | ( _4869 ) ;
 assign _4872 = ( n_n1132 ) | ( n_n1176 ) ;
 assign _4873 = ( n_n1283 ) | ( n_n1259 ) ;
 assign _4874 = ( n_n955 ) | ( n_n1109 ) ;
 assign _4875 = ( _206 ) | ( n_n941 ) ;
 assign _4876 = ( _4873 ) | ( _4872 ) ;
 assign _4877 = ( _4875 ) | ( _4874 ) ;
 assign _4878 = ( _208 ) | ( _50 ) ;
 assign _4879 = ( _4878 ) | ( _130 ) ;
 assign _4880 = ( n_n87  &  n_n70 ) ;
 assign _4881 = ( n_n58  &  _315 ) ;
 assign _4882 = ( _51 ) | ( n_n1217 ) ;
 assign _4883 = ( _138 ) | ( _137 ) ;
 assign _4884 = ( _56 ) | ( _841 ) ;
 assign _4885 = ( _4882 ) | ( _104 ) ;
 assign _4886 = ( _4884 ) | ( _4883 ) ;
 assign _4887 = ( n_n76  &  n_n86 ) ;
 assign _4888 = ( _59 ) | ( n_n1176 ) ;
 assign _4889 = ( _185 ) | ( _162 ) ;
 assign _4890 = ( _90 ) | ( _273 ) ;
 assign _4891 = ( _4888 ) | ( _286 ) ;
 assign _4892 = ( _4890 ) | ( _4889 ) ;
 assign _4893 = ( i_2_  &  (~ i_1_) ) ;
 assign _4894 = ( _4893  &  _328 ) ;
 assign _4895 = ( _78 ) | ( _833 ) ;
 assign _4896 = ( _163 ) | ( _154 ) ;
 assign _4897 = ( _834 ) | ( _239 ) ;
 assign _4898 = ( _4896 ) | ( _4895 ) ;
 assign _4899 = ( _80 ) | ( n_n1144 ) ;
 assign _4900 = ( _4899 ) | ( _148 ) ;
 assign _4901 = ( wire4813 ) | ( _4900 ) ;
 assign _4902 = ( n_n666 ) | ( n_n665 ) ;
 assign _4903 = ( n_n943 ) | ( n_n956 ) ;
 assign _4904 = ( _97 ) | ( n_n944 ) ;
 assign _4905 = ( _214 ) | ( _207 ) ;
 assign _4906 = ( _4904 ) | ( _4903 ) ;
 assign _4907 = ( n_n83  &  n_n70 ) ;
 assign _4908 = ( n_n91  &  _328 ) ;
 assign _4909 = ( i_2_  &  i_1_ ) ;
 assign _4910 = ( _313  &  n_n64 ) ;
 assign _4911 = ( n_n990 ) | ( _827 ) ;
 assign _4912 = ( n_n993 ) | ( n_n989 ) ;
 assign _4913 = ( n_n982 ) | ( n_n977 ) ;
 assign _4914 = ( _4912 ) | ( _4911 ) ;
 assign _4915 = ( n_n962 ) | ( n_n968 ) ;
 assign _4916 = ( _215 ) | ( _210 ) ;
 assign _4917 = ( n_n973 ) | ( n_n974 ) ;
 assign _4918 = ( _4917 ) | ( n_n970 ) ;
 assign _4919 = ( _4918 ) | ( n_n716 ) ;
 assign _4920 = ( wire4877 ) | ( wire4873 ) ;
 assign _4921 = ( n_n676 ) | ( _4919 ) ;
 assign _4922 = ( n_n79  &  n_n70 ) ;
 assign _4923 = ( _60 ) | ( n_n1074 ) ;
 assign _4924 = ( _126 ) | ( _69 ) ;
 assign _4925 = ( _49 ) | ( _240 ) ;
 assign _4926 = ( _4923 ) | ( _244 ) ;
 assign _4927 = ( _4925 ) | ( _4924 ) ;
 assign _4928 = ( n_n1088 ) | ( n_n1087 ) ;
 assign _4929 = ( n_n1081 ) | ( n_n1078 ) ;
 assign _4930 = ( _71 ) | ( n_n1093 ) ;
 assign _4931 = ( _102 ) | ( _155 ) ;
 assign _4932 = ( _4929 ) | ( _4928 ) ;
 assign _4933 = ( _4931 ) | ( _4930 ) ;
 assign _4934 = ( n_n101  &  _328 ) ;
 assign _4935 = ( n_n90  &  _35 ) ;
 assign _4936 = ( n_n1118 ) | ( n_n1121 ) ;
 assign _4937 = ( _127 ) | ( _85 ) ;
 assign _4938 = ( _4936 ) | ( _243 ) ;
 assign _4939 = ( n_n874 ) | ( _4937 ) ;
 assign _4940 = ( n_n1006 ) | ( n_n1004 ) ;
 assign _4941 = ( n_n1058 ) | ( n_n1060 ) ;
 assign _4942 = ( _143 ) | ( n_n1047 ) ;
 assign _4943 = ( _152 ) | ( _818 ) ;
 assign _4944 = ( _4941 ) | ( _200 ) ;
 assign _4945 = ( _4943 ) | ( _4942 ) ;
 assign _4946 = ( n_n83  &  n_n52 ) ;
 assign _4947 = ( n_n1032 ) | ( _129 ) ;
 assign _4948 = ( n_n1026 ) | ( n_n1018 ) ;
 assign _4949 = ( _145 ) | ( _77 ) ;
 assign _4950 = ( _4947 ) | ( _212 ) ;
 assign _4951 = ( _4949 ) | ( _4948 ) ;
 assign _4952 = ( _327  &  (~ i_3_) ) ;
 assign _4953 = ( n_n999 ) | ( _812 ) ;
 assign _4954 = ( n_n1011 ) | ( n_n1009 ) ;
 assign _4955 = ( _220 ) | ( n_n1001 ) ;
 assign _4956 = ( _4954 ) | ( _4953 ) ;
 assign _4957 = ( wire4836 ) | ( n_n641 ) ;
 assign _4958 = ( n_n669 ) | ( n_n670 ) ;
 assign _4959 = ( n_n671 ) | ( n_n668 ) ;
 assign _4960 = ( _4957 ) | ( n_n672 ) ;
 assign _4961 = ( _4959 ) | ( _4958 ) ;
 assign _4962 = ( n_n95  &  _302 ) ;
 assign _4963 = ( n_n100  &  n_n64 ) ;
 assign _4964 = ( _26  &  (~ i_0_) ) ;
 assign _4965 = ( _171 ) | ( _72 ) ;
 assign _4966 = ( _173 ) | ( _172 ) ;
 assign _4967 = ( _246 ) | ( _174 ) ;
 assign _4968 = ( _88 ) | ( _804 ) ;
 assign _4969 = ( _4966 ) | ( _4965 ) ;
 assign _4970 = ( _4968 ) | ( _4967 ) ;
 assign _4971 = ( _177 ) | ( _125 ) ;
 assign _4972 = ( _800 ) | ( _799 ) ;
 assign _4973 = ( _798 ) | ( _176 ) ;
 assign _4974 = ( _4972 ) | ( _4971 ) ;
 assign _4975 = ( _55 ) | ( n_n1294 ) ;
 assign _4976 = ( _231 ) | ( _100 ) ;
 assign _4977 = ( _92 ) | ( _289 ) ;
 assign _4978 = ( _4975 ) | ( _150 ) ;
 assign _4979 = ( _4977 ) | ( _4976 ) ;
 assign _4980 = ( n_n664 ) | ( n_n662 ) ;
 assign _4981 = ( _4980 ) | ( n_n663 ) ;
 assign _4982 = ( n_n661 ) | ( n_n658 ) ;
 assign _4983 = ( wire4879 ) | ( _4981 ) ;
 assign _4984 = ( n_n66  &  n_n70 ) ;
 assign _4985 = ( n_n976 ) | ( n_n980 ) ;
 assign _4986 = ( _99 ) | ( _58 ) ;
 assign _4987 = ( _255 ) | ( _209 ) ;
 assign _4988 = ( _4986 ) | ( _4985 ) ;
 assign _4989 = ( n_n1043 ) | ( n_n1045 ) ;
 assign _4990 = ( n_n1032 ) | ( n_n1048 ) ;
 assign _4991 = ( n_n1030 ) | ( n_n1036 ) ;
 assign _4992 = ( _227 ) | ( _68 ) ;
 assign _4993 = ( _4990 ) | ( _4989 ) ;
 assign _4994 = ( _4992 ) | ( _4991 ) ;
 assign _4995 = ( n_n1070 ) | ( n_n1074 ) ;
 assign _4996 = ( _126 ) | ( _75 ) ;
 assign _4997 = ( _786 ) | ( _168 ) ;
 assign _4998 = ( _4996 ) | ( _4995 ) ;
 assign _4999 = ( n_n1077 ) | ( n_n1082 ) ;
 assign _5000 = ( _4999 ) | ( n_n1078 ) ;
 assign _5001 = ( n_n1055 ) | ( n_n1060 ) ;
 assign _5002 = ( n_n1057 ) | ( n_n1058 ) ;
 assign _5003 = ( _107 ) | ( n_n1059 ) ;
 assign _5004 = ( _5002 ) | ( _5001 ) ;
 assign _5005 = ( n_n1052 ) | ( n_n1054 ) ;
 assign _5006 = ( _5005 ) | ( _780 ) ;
 assign _5007 = ( wire4914 ) | ( _5006 ) ;
 assign _5008 = ( n_n596 ) | ( n_n598 ) ;
 assign _5009 = ( i_6_  &  i_8_ ) ;
 assign _5010 = ( n_n967 ) | ( n_n964 ) ;
 assign _5011 = ( _52 ) | ( n_n957 ) ;
 assign _5012 = ( _210 ) | ( _57 ) ;
 assign _5013 = ( _5011 ) | ( _5010 ) ;
 assign _5014 = ( n_n80  &  n_n86 ) ;
 assign _5015 = ( n_n949 ) | ( n_n950 ) ;
 assign _5016 = ( n_n956 ) | ( n_n951 ) ;
 assign _5017 = ( n_n954 ) | ( n_n953 ) ;
 assign _5018 = ( n_n955 ) | ( n_n952 ) ;
 assign _5019 = ( _5017 ) | ( _5016 ) ;
 assign _5020 = ( n_n652 ) | ( _5018 ) ;
 assign _5021 = ( _5020 ) | ( _5019 ) ;
 assign _5022 = ( n_n83  &  i_3_ ) ;
 assign _5023 = ( n_n54  &  i_7_ ) ;
 assign _5024 = ( n_n1025 ) | ( n_n1001 ) ;
 assign _5025 = ( _268 ) | ( _64 ) ;
 assign _5026 = ( _771 ) | ( _279 ) ;
 assign _5027 = ( _5025 ) | ( _5024 ) ;
 assign _5028 = ( n_n641 ) | ( _5026 ) ;
 assign _5029 = ( n_n987 ) | ( n_n995 ) ;
 assign _5030 = ( n_n986 ) | ( n_n990 ) ;
 assign _5031 = ( n_n993 ) | ( n_n994 ) ;
 assign _5032 = ( _132 ) | ( _181 ) ;
 assign _5033 = ( _5030 ) | ( _5029 ) ;
 assign _5034 = ( _5032 ) | ( _5031 ) ;
 assign _5035 = ( n_n86  &  (~ i_3_) ) ;
 assign _5036 = ( (~ i_4_)  &  i_3_ ) ;
 assign _5037 = ( _5036  &  _326 ) ;
 assign _5038 = ( _89 ) | ( n_n944 ) ;
 assign _5039 = ( wire4934 ) | ( n_n654 ) ;
 assign _5040 = ( n_n599 ) | ( n_n601 ) ;
 assign _5041 = ( _5039 ) | ( n_n600 ) ;
 assign _5042 = ( _5040 ) | ( wire4935 ) ;
 assign _5043 = ( n_n584 ) | ( _5041 ) ;
 assign _5044 = ( _83 ) | ( _81 ) ;
 assign _5045 = ( _248 ) | ( _231 ) ;
 assign _5046 = ( _112 ) | ( _249 ) ;
 assign _5047 = ( _5044 ) | ( _150 ) ;
 assign _5048 = ( _5046 ) | ( _5045 ) ;
 assign _5049 = ( _131 ) | ( _50 ) ;
 assign _5050 = ( _758 ) | ( _250 ) ;
 assign _5051 = ( _94 ) | ( _759 ) ;
 assign _5052 = ( _5049 ) | ( _165 ) ;
 assign _5053 = ( _5051 ) | ( _5050 ) ;
 assign _5054 = ( _48 ) | ( n_n1267 ) ;
 assign _5055 = ( _183 ) | ( _72 ) ;
 assign _5056 = ( _5054 ) | ( _753 ) ;
 assign _5057 = ( _142 ) | ( _140 ) ;
 assign _5058 = ( _56 ) | ( _749 ) ;
 assign _5059 = ( _748 ) | ( _747 ) ;
 assign _5060 = ( _5058 ) | ( _5057 ) ;
 assign _5061 = ( n_n90  &  n_n64 ) ;
 assign _5062 = ( _74 ) | ( _73 ) ;
 assign _5063 = ( _224 ) | ( _173 ) ;
 assign _5064 = ( _741 ) | ( _740 ) ;
 assign _5065 = ( _5062 ) | ( _70 ) ;
 assign _5066 = ( _5064 ) | ( _5063 ) ;
 assign _5067 = ( n_n1170 ) | ( n_n1176 ) ;
 assign _5068 = ( n_n1174 ) | ( n_n1177 ) ;
 assign _5069 = ( _734 ) | ( _59 ) ;
 assign _5070 = ( _5068 ) | ( _5067 ) ;
 assign _5071 = ( _274 ) | ( n_n1181 ) ;
 assign _5072 = ( _5071 ) | ( _275 ) ;
 assign _5073 = ( n_n590 ) | ( _5072 ) ;
 assign _5074 = ( n_n591 ) | ( wire4977 ) ;
 assign _5075 = ( n_n58  &  _315 ) ;
 assign _5076 = ( _119 ) | ( n_n1281 ) ;
 assign _5077 = ( _5076 ) | ( _180 ) ;
 assign _5078 = ( wire4956 ) | ( _5077 ) ;
 assign _5079 = ( n_n587 ) | ( n_n588 ) ;
 assign _5080 = ( _5079 ) | ( _5078 ) ;
 assign _5081 = ( (~ i_4_)  &  i_3_ ) ;
 assign _5082 = ( n_n95  &  _5081 ) ;
 assign _5083 = ( i_6_  &  i_8_ ) ;
 assign _5084 = ( _5083  &  _35 ) ;
 assign _5085 = ( n_n1095 ) | ( _724 ) ;
 assign _5086 = ( n_n1103 ) | ( n_n1105 ) ;
 assign _5087 = ( _155 ) | ( n_n1101 ) ;
 assign _5088 = ( _245 ) | ( _257 ) ;
 assign _5089 = ( _5086 ) | ( _5085 ) ;
 assign _5090 = ( _5088 ) | ( _5087 ) ;
 assign _5091 = ( _134 ) | ( n_n1156 ) ;
 assign _5092 = ( _164 ) | ( _135 ) ;
 assign _5093 = ( _5091 ) | ( _717 ) ;
 assign _5094 = ( i_3_  &  i_7_ ) ;
 assign _5095 = ( _5094  &  _340 ) ;
 assign _5096 = ( n_n54  &  i_8_ ) ;
 assign _5097 = ( n_n1122 ) | ( _709 ) ;
 assign _5098 = ( _103 ) | ( n_n1118 ) ;
 assign _5099 = ( _199 ) | ( _128 ) ;
 assign _5100 = ( _243 ) | ( _710 ) ;
 assign _5101 = ( _5098 ) | ( _5097 ) ;
 assign _5102 = ( _5100 ) | ( _5099 ) ;
 assign _5103 = ( _80 ) | ( n_n1128 ) ;
 assign _5104 = ( _5103 ) | ( _190 ) ;
 assign _5105 = ( wire4985 ) | ( _5104 ) ;
 assign _5106 = ( n_n594 ) | ( n_n595 ) ;
 assign _5107 = ( _5106 ) | ( _5105 ) ;
 assign _5108 = ( wire5003 ) | ( _5107 ) ;
 assign _5109 = ( n_n953 ) | ( n_n951 ) ;
 assign _5110 = ( n_n960 ) | ( n_n958 ) ;
 assign _5111 = ( n_n959 ) | ( n_n950 ) ;
 assign _5112 = ( _5110 ) | ( _5109 ) ;
 assign _5113 = ( n_n957 ) | ( n_n956 ) ;
 assign _5114 = ( _5113 ) | ( n_n954 ) ;
 assign _5115 = ( n_n962 ) | ( n_n964 ) ;
 assign _5116 = ( n_n961 ) | ( n_n971 ) ;
 assign _5117 = ( _99 ) | ( _287 ) ;
 assign _5118 = ( _5115 ) | ( _209 ) ;
 assign _5119 = ( _5117 ) | ( _5116 ) ;
 assign _5120 = ( _89 ) | ( _178 ) ;
 assign _5121 = ( _282 ) | ( n_n654 ) ;
 assign _5122 = ( _5121 ) | ( _5120 ) ;
 assign _5123 = ( n_n465 ) | ( n_n466 ) ;
 assign _5124 = ( i_4_  &  (~ i_5_) ) ;
 assign _5125 = ( n_n1006 ) | ( n_n1011 ) ;
 assign _5126 = ( n_n1010 ) | ( n_n1001 ) ;
 assign _5127 = ( _702 ) | ( _76 ) ;
 assign _5128 = ( _5126 ) | ( _5125 ) ;
 assign _5129 = ( n_n882 ) | ( _5127 ) ;
 assign _5130 = ( n_n83  &  n_n86 ) ;
 assign _5131 = ( n_n1025 ) | ( n_n1022 ) ;
 assign _5132 = ( _62 ) | ( n_n1026 ) ;
 assign _5133 = ( _696 ) | ( _68 ) ;
 assign _5134 = ( _5132 ) | ( _5131 ) ;
 assign _5135 = ( n_n994 ) | ( n_n991 ) ;
 assign _5136 = ( n_n978 ) | ( n_n989 ) ;
 assign _5137 = ( _5135 ) | ( _132 ) ;
 assign _5138 = ( n_n504 ) | ( _5136 ) ;
 assign _5139 = ( n_n1019 ) | ( n_n1013 ) ;
 assign _5140 = ( _5139 ) | ( _279 ) ;
 assign _5141 = ( wire5079 ) | ( _5140 ) ;
 assign _5142 = ( n_n464 ) | ( n_n463 ) ;
 assign _5143 = ( _5142 ) | ( _5141 ) ;
 assign _5144 = ( _143 ) | ( _75 ) ;
 assign _5145 = ( n_n97  &  n_n70 ) ;
 assign _5146 = ( n_n1055 ) | ( n_n1060 ) ;
 assign _5147 = ( n_n1057 ) | ( n_n1058 ) ;
 assign _5148 = ( _295 ) | ( n_n1059 ) ;
 assign _5149 = ( _5147 ) | ( _5146 ) ;
 assign _5150 = ( n_n421 ) | ( _5148 ) ;
 assign _5151 = ( n_n1074 ) | ( n_n1087 ) ;
 assign _5152 = ( n_n1079 ) | ( n_n1077 ) ;
 assign _5153 = ( _147 ) | ( n_n1070 ) ;
 assign _5154 = ( _5152 ) | ( _5151 ) ;
 assign _5155 = ( n_n1093 ) | ( n_n1100 ) ;
 assign _5156 = ( _5155 ) | ( n_n1101 ) ;
 assign _5157 = ( _304  &  _35 ) ;
 assign _5158 = ( n_n1045 ) | ( _196 ) ;
 assign _5159 = ( n_n1043 ) | ( n_n1046 ) ;
 assign _5160 = ( _687 ) | ( n_n1035 ) ;
 assign _5161 = ( _5159 ) | ( _5158 ) ;
 assign _5162 = ( _61 ) | ( n_n1052 ) ;
 assign _5163 = ( _5162 ) | ( _283 ) ;
 assign _5164 = ( wire5100 ) | ( _5163 ) ;
 assign _5165 = ( n_n459 ) | ( n_n460 ) ;
 assign _5166 = ( _5165 ) | ( _5164 ) ;
 assign _5167 = ( _296  &  (~ i_0_) ) ;
 assign _5168 = ( n_n83  &  _326 ) ;
 assign _5169 = ( n_n96  &  n_n75 ) ;
 assign _5170 = ( n_n1217 ) | ( n_n1216 ) ;
 assign _5171 = ( _192 ) | ( _191 ) ;
 assign _5172 = ( _681 ) | ( _267 ) ;
 assign _5173 = ( _5171 ) | ( _5170 ) ;
 assign _5174 = ( _48 ) | ( n_n1259 ) ;
 assign _5175 = ( _277 ) | ( _276 ) ;
 assign _5176 = ( _676 ) | ( _675 ) ;
 assign _5177 = ( _5175 ) | ( _5174 ) ;
 assign _5178 = ( _26  &  (~ i_1_) ) ;
 assign _5179 = ( _197 ) | ( _74 ) ;
 assign _5180 = ( _5179 ) | ( _671 ) ;
 assign _5181 = ( n_n1184 ) | ( n_n1176 ) ;
 assign _5182 = ( _198 ) | ( n_n1172 ) ;
 assign _5183 = ( _664 ) | ( _274 ) ;
 assign _5184 = ( _5181 ) | ( _238 ) ;
 assign _5185 = ( _5183 ) | ( _5182 ) ;
 assign _5186 = ( _109 ) | ( _108 ) ;
 assign _5187 = ( _658 ) | ( _228 ) ;
 assign _5188 = ( _660 ) | ( _659 ) ;
 assign _5189 = ( _5187 ) | ( _5186 ) ;
 assign _5190 = ( _110 ) | ( n_n1286 ) ;
 assign _5191 = ( _230 ) | ( _122 ) ;
 assign _5192 = ( _288 ) | ( _260 ) ;
 assign _5193 = ( _5191 ) | ( _5190 ) ;
 assign _5194 = ( _5193 ) | ( _5192 ) ;
 assign _5195 = ( _652 ) | ( _66 ) ;
 assign _5196 = ( wire5010 ) | ( _5195 ) ;
 assign _5197 = ( n_n453 ) | ( n_n455 ) ;
 assign _5198 = ( _5196 ) | ( n_n446 ) ;
 assign _5199 = ( n_n94  &  n_n64 ) ;
 assign _5200 = ( n_n93  &  _302 ) ;
 assign _5201 = ( n_n1118 ) | ( n_n1108 ) ;
 assign _5202 = ( _124 ) | ( _85 ) ;
 assign _5203 = ( _202 ) | ( _199 ) ;
 assign _5204 = ( _5202 ) | ( _5201 ) ;
 assign _5205 = ( n_n1125 ) | ( n_n1128 ) ;
 assign _5206 = ( _5205 ) | ( _127 ) ;
 assign _5207 = ( _305  &  n_n70 ) ;
 assign _5208 = ( n_n1145 ) | ( _646 ) ;
 assign _5209 = ( _80 ) | ( n_n1134 ) ;
 assign _5210 = ( _161 ) | ( _135 ) ;
 assign _5211 = ( _5209 ) | ( _5208 ) ;
 assign _5212 = ( n_n1146 ) | ( n_n1164 ) ;
 assign _5213 = ( n_n1153 ) | ( n_n1163 ) ;
 assign _5214 = ( _640 ) | ( n_n1158 ) ;
 assign _5215 = ( _5213 ) | ( _5212 ) ;
 assign _5216 = ( _84 ) | ( n_n1169 ) ;
 assign _5217 = ( _5216 ) | ( _154 ) ;
 assign _5218 = ( n_n1130 ) | ( n_n1132 ) ;
 assign _5219 = ( _5218 ) | ( _190 ) ;
 assign _5220 = ( wire5042 ) | ( _5219 ) ;
 assign _5221 = ( n_n456 ) | ( n_n458 ) ;
 assign _5222 = ( _5221 ) | ( _5220 ) ;
 assign _5223 = ( _5222 ) | ( wire5056 ) ;
 assign _5224 = ( n_n1068 ) | ( n_n1058 ) ;
 assign _5225 = ( _60 ) | ( n_n1057 ) ;
 assign _5226 = ( _143 ) | ( _107 ) ;
 assign _5227 = ( _5225 ) | ( _5224 ) ;
 assign _5228 = ( n_n1095 ) | ( n_n1100 ) ;
 assign _5229 = ( _71 ) | ( n_n1079 ) ;
 assign _5230 = ( _115 ) | ( _111 ) ;
 assign _5231 = ( _5229 ) | ( _5228 ) ;
 assign _5232 = ( n_n1101 ) | ( n_n1103 ) ;
 assign _5233 = ( _5232 ) | ( _114 ) ;
 assign _5234 = ( n_n97  &  _35 ) ;
 assign _5235 = ( n_n1122 ) | ( n_n1132 ) ;
 assign _5236 = ( _80 ) | ( n_n1134 ) ;
 assign _5237 = ( _265 ) | ( _190 ) ;
 assign _5238 = ( _5236 ) | ( _5235 ) ;
 assign _5239 = ( n_n77  &  i_1_ ) ;
 assign _5240 = ( _124 ) | ( n_n1121 ) ;
 assign _5241 = ( _5240 ) | ( _636 ) ;
 assign _5242 = ( n_n1014 ) | ( n_n1013 ) ;
 assign _5243 = ( n_n1021 ) | ( n_n1019 ) ;
 assign _5244 = ( _5242 ) | ( _213 ) ;
 assign _5245 = ( n_n295 ) | ( _5243 ) ;
 assign _5246 = ( n_n1032 ) | ( n_n1047 ) ;
 assign _5247 = ( n_n1028 ) | ( n_n1039 ) ;
 assign _5248 = ( _145 ) | ( _62 ) ;
 assign _5249 = ( _5246 ) | ( _217 ) ;
 assign _5250 = ( _5248 ) | ( _5247 ) ;
 assign _5251 = ( n_n991 ) | ( n_n990 ) ;
 assign _5252 = ( n_n980 ) | ( n_n986 ) ;
 assign _5253 = ( n_n993 ) | ( n_n1001 ) ;
 assign _5254 = ( _132 ) | ( _181 ) ;
 assign _5255 = ( _5252 ) | ( _5251 ) ;
 assign _5256 = ( _5254 ) | ( _5253 ) ;
 assign _5257 = ( n_n953 ) | ( n_n957 ) ;
 assign _5258 = ( n_n950 ) | ( n_n954 ) ;
 assign _5259 = ( _214 ) | ( n_n955 ) ;
 assign _5260 = ( _5257 ) | ( _221 ) ;
 assign _5261 = ( _5259 ) | ( _5258 ) ;
 assign _5262 = ( n_n969 ) | ( n_n964 ) ;
 assign _5263 = ( n_n978 ) | ( n_n977 ) ;
 assign _5264 = ( _58 ) | ( n_n959 ) ;
 assign _5265 = ( _57 ) | ( _624 ) ;
 assign _5266 = ( _5263 ) | ( _5262 ) ;
 assign _5267 = ( _5265 ) | ( _5264 ) ;
 assign _5268 = ( n_n944 ) | ( n_n947 ) ;
 assign _5269 = ( _5268 ) | ( _178 ) ;
 assign _5270 = ( _282 ) | ( n_n654 ) ;
 assign _5271 = ( _5270 ) | ( _5269 ) ;
 assign _5272 = ( n_n532 ) | ( n_n533 ) ;
 assign _5273 = ( n_n529 ) | ( n_n530 ) ;
 assign _5274 = ( _5273 ) | ( n_n531 ) ;
 assign _5275 = ( _283 ) | ( _61 ) ;
 assign _5276 = ( _5275 ) | ( _295 ) ;
 assign _5277 = ( wire5164 ) | ( _5276 ) ;
 assign _5278 = ( n_n526 ) | ( n_n527 ) ;
 assign _5279 = ( _5278 ) | ( _5277 ) ;
 assign _5280 = ( _48 ) | ( n_n1279 ) ;
 assign _5281 = ( _182 ) | ( _72 ) ;
 assign _5282 = ( _616 ) | ( _183 ) ;
 assign _5283 = ( _92 ) | ( _617 ) ;
 assign _5284 = ( _5281 ) | ( _5280 ) ;
 assign _5285 = ( _5283 ) | ( _5282 ) ;
 assign _5286 = ( n_n78  &  _303 ) ;
 assign _5287 = ( _169 ) | ( _156 ) ;
 assign _5288 = ( _293 ) | ( _201 ) ;
 assign _5289 = ( _611 ) | ( _610 ) ;
 assign _5290 = ( _5288 ) | ( _5287 ) ;
 assign _5291 = ( n_n1297 ) | ( n_n1283 ) ;
 assign _5292 = ( _151 ) | ( n_n1312 ) ;
 assign _5293 = ( _230 ) | ( _157 ) ;
 assign _5294 = ( _112 ) | ( _248 ) ;
 assign _5295 = ( _5292 ) | ( _5291 ) ;
 assign _5296 = ( _5294 ) | ( _5293 ) ;
 assign _5297 = ( n_n1193 ) | ( n_n1184 ) ;
 assign _5298 = ( _59 ) | ( n_n1188 ) ;
 assign _5299 = ( _604 ) | ( _186 ) ;
 assign _5300 = ( _5298 ) | ( _5297 ) ;
 assign _5301 = ( n_n71  &  n_n64 ) ;
 assign _5302 = ( n_n1204 ) | ( n_n1216 ) ;
 assign _5303 = ( _123 ) | ( _66 ) ;
 assign _5304 = ( _235 ) | ( _194 ) ;
 assign _5305 = ( _286 ) | ( _596 ) ;
 assign _5306 = ( _5303 ) | ( _5302 ) ;
 assign _5307 = ( _5305 ) | ( _5304 ) ;
 assign _5308 = ( n_n1145 ) | ( n_n1146 ) ;
 assign _5309 = ( n_n1158 ) | ( n_n1156 ) ;
 assign _5310 = ( _5308 ) | ( _218 ) ;
 assign _5311 = ( n_n554 ) | ( _5309 ) ;
 assign _5312 = ( _108 ) | ( _82 ) ;
 assign _5313 = ( _228 ) | ( _117 ) ;
 assign _5314 = ( _590 ) | ( _272 ) ;
 assign _5315 = ( _5313 ) | ( _5312 ) ;
 assign _5316 = ( _297  &  _40 ) ;
 assign _5317 = ( n_n1169 ) | ( _583 ) ;
 assign _5318 = ( _5317 ) | ( _63 ) ;
 assign _5319 = ( wire5108 ) | ( _5318 ) ;
 assign _5320 = ( n_n523 ) | ( n_n519 ) ;
 assign _5321 = ( _5319 ) | ( n_n525 ) ;
 assign _5322 = ( n_n94  &  _303 ) ;
 assign _5323 = ( _193 ) | ( n_n1254 ) ;
 assign _5324 = ( _5323 ) | ( _224 ) ;
 assign _5325 = ( wire5130 ) | ( _5324 ) ;
 assign _5326 = ( n_n520 ) | ( n_n521 ) ;
 assign _5327 = ( _5326 ) | ( _5325 ) ;
 assign _5328 = ( _5327 ) | ( wire5136 ) ;
 assign _5329 = ( _151 ) | ( _113 ) ;
 assign _5330 = ( _232 ) | ( _231 ) ;
 assign _5331 = ( _573 ) | ( _233 ) ;
 assign _5332 = ( _205 ) | ( _574 ) ;
 assign _5333 = ( _5330 ) | ( _5329 ) ;
 assign _5334 = ( _5332 ) | ( _5331 ) ;
 assign _5335 = ( _50 ) | ( n_n1331 ) ;
 assign _5336 = ( _567 ) | ( _288 ) ;
 assign _5337 = ( _569 ) | ( _568 ) ;
 assign _5338 = ( _5336 ) | ( _5335 ) ;
 assign _5339 = ( _173 ) | ( _138 ) ;
 assign _5340 = ( _193 ) | ( _188 ) ;
 assign _5341 = ( _561 ) | ( _194 ) ;
 assign _5342 = ( _5340 ) | ( _5339 ) ;
 assign _5343 = ( _26  &  (~ i_1_) ) ;
 assign _5344 = ( n_n97  &  _297 ) ;
 assign _5345 = ( _182 ) | ( n_n1259 ) ;
 assign _5346 = ( _556 ) | ( _254 ) ;
 assign _5347 = ( _5345 ) | ( _557 ) ;
 assign _5348 = ( _249 ) | ( _79 ) ;
 assign _5349 = ( _5348 ) | ( _277 ) ;
 assign _5350 = ( n_n54  &  n_n70 ) ;
 assign _5351 = ( _269 ) | ( n_n1215 ) ;
 assign _5352 = ( _5351 ) | ( _549 ) ;
 assign _5353 = ( n_n310 ) | ( _5352 ) ;
 assign _5354 = ( n_n311 ) | ( wire5192 ) ;
 assign _5355 = ( _5353 ) | ( n_n312 ) ;
 assign _5356 = ( n_n1193 ) | ( n_n1181 ) ;
 assign _5357 = ( _198 ) | ( n_n1185 ) ;
 assign _5358 = ( _543 ) | ( _274 ) ;
 assign _5359 = ( _5357 ) | ( _5356 ) ;
 assign _5360 = ( _84 ) | ( n_n1172 ) ;
 assign _5361 = ( _5360 ) | ( _154 ) ;
 assign _5362 = ( n_n40  &  n_n70 ) ;
 assign _5363 = ( _192 ) | ( n_n1204 ) ;
 assign _5364 = ( _278 ) | ( _270 ) ;
 assign _5365 = ( _538 ) | ( _537 ) ;
 assign _5366 = ( _5364 ) | ( _5363 ) ;
 assign _5367 = ( _66 ) | ( _51 ) ;
 assign _5368 = ( _5367 ) | ( _186 ) ;
 assign _5369 = ( (~ i_1_)  &  (~ i_4_) ) ;
 assign _5370 = ( _5369  &  _298 ) ;
 assign _5371 = ( n_n1147 ) | ( _531 ) ;
 assign _5372 = ( n_n1144 ) | ( n_n1134 ) ;
 assign _5373 = ( _149 ) | ( _148 ) ;
 assign _5374 = ( _5372 ) | ( _5371 ) ;
 assign _5375 = ( _78 ) | ( n_n1160 ) ;
 assign _5376 = ( _5375 ) | ( _163 ) ;
 assign _5377 = ( wire5214 ) | ( _5376 ) ;
 assign _5378 = ( n_n314 ) | ( n_n315 ) ;
 assign _5379 = ( _5378 ) | ( _5377 ) ;
 assign _5380 = ( n_n970 ) | ( n_n971 ) ;
 assign _5381 = ( n_n939 ) | ( n_n943 ) ;
 assign _5382 = ( n_n944 ) | ( n_n947 ) ;
 assign _5383 = ( n_n949 ) | ( n_n942 ) ;
 assign _5384 = ( _207 ) | ( _178 ) ;
 assign _5385 = ( _5382 ) | ( _5381 ) ;
 assign _5386 = ( _5384 ) | ( _5383 ) ;
 assign _5387 = ( n_n967 ) | ( n_n951 ) ;
 assign _5388 = ( n_n960 ) | ( n_n957 ) ;
 assign _5389 = ( _52 ) | ( _524 ) ;
 assign _5390 = ( _5387 ) | ( _97 ) ;
 assign _5391 = ( _5389 ) | ( _5388 ) ;
 assign _5392 = ( n_n980 ) | ( n_n974 ) ;
 assign _5393 = ( n_n977 ) | ( n_n981 ) ;
 assign _5394 = ( _5392 ) | ( _132 ) ;
 assign _5395 = ( n_n365 ) | ( _5393 ) ;
 assign _5396 = ( _5395 ) | ( _5394 ) ;
 assign _5397 = ( n_n324 ) | ( n_n325 ) ;
 assign _5398 = ( _297  &  n_n73 ) ;
 assign _5399 = ( n_n991 ) | ( n_n990 ) ;
 assign _5400 = ( n_n984 ) | ( n_n994 ) ;
 assign _5401 = ( _98 ) | ( _64 ) ;
 assign _5402 = ( _5399 ) | ( _211 ) ;
 assign _5403 = ( _5401 ) | ( _5400 ) ;
 assign _5404 = ( n_n1022 ) | ( n_n1042 ) ;
 assign _5405 = ( _62 ) | ( n_n1028 ) ;
 assign _5406 = ( _226 ) | ( _268 ) ;
 assign _5407 = ( _5404 ) | ( _227 ) ;
 assign _5408 = ( _5406 ) | ( _5405 ) ;
 assign _5409 = ( n_n1006 ) | ( n_n1009 ) ;
 assign _5410 = ( n_n1014 ) | ( n_n1010 ) ;
 assign _5411 = ( n_n1002 ) | ( n_n1019 ) ;
 assign _5412 = ( _144 ) | ( _77 ) ;
 assign _5413 = ( _5410 ) | ( _5409 ) ;
 assign _5414 = ( _5412 ) | ( _5411 ) ;
 assign _5415 = ( n_n320 ) | ( n_n322 ) ;
 assign _5416 = ( n_n1048 ) | ( n_n1055 ) ;
 assign _5417 = ( _61 ) | ( n_n1057 ) ;
 assign _5418 = ( _107 ) | ( _75 ) ;
 assign _5419 = ( _5417 ) | ( _5416 ) ;
 assign _5420 = ( n_n1070 ) | ( n_n1068 ) ;
 assign _5421 = ( _5420 ) | ( _126 ) ;
 assign _5422 = ( n_n1122 ) | ( n_n1132 ) ;
 assign _5423 = ( n_n1120 ) | ( n_n1130 ) ;
 assign _5424 = ( _127 ) | ( n_n1117 ) ;
 assign _5425 = ( _5423 ) | ( _5422 ) ;
 assign _5426 = ( n_n1077 ) | ( n_n1087 ) ;
 assign _5427 = ( n_n1081 ) | ( n_n1091 ) ;
 assign _5428 = ( _147 ) | ( _71 ) ;
 assign _5429 = ( _245 ) | ( _168 ) ;
 assign _5430 = ( _5427 ) | ( _5426 ) ;
 assign _5431 = ( _5429 ) | ( _5428 ) ;
 assign _5432 = ( n_n66  &  (~ i_7_) ) ;
 assign _5433 = ( _199 ) | ( n_n1108 ) ;
 assign _5434 = ( _5433 ) | ( _513 ) ;
 assign _5435 = ( wire5234 ) | ( _5434 ) ;
 assign _5436 = ( n_n318 ) | ( n_n319 ) ;
 assign _5437 = ( _5436 ) | ( _5435 ) ;
 assign _5438 = ( n_n303 ) | ( n_n309 ) ;
 assign _5439 = ( _304  &  n_n70 ) ;
 assign _5440 = ( n_n1092 ) | ( _507 ) ;
 assign _5441 = ( n_n1095 ) | ( n_n1100 ) ;
 assign _5442 = ( _147 ) | ( n_n1091 ) ;
 assign _5443 = ( _5441 ) | ( _5440 ) ;
 assign _5444 = ( n_n1117 ) | ( n_n1109 ) ;
 assign _5445 = ( _128 ) | ( _124 ) ;
 assign _5446 = ( _202 ) | ( _199 ) ;
 assign _5447 = ( _5445 ) | ( _5444 ) ;
 assign _5448 = ( n_n1108 ) | ( n_n1105 ) ;
 assign _5449 = ( _5448 ) | ( _155 ) ;
 assign _5450 = ( n_n1177 ) | ( n_n1169 ) ;
 assign _5451 = ( _63 ) | ( _59 ) ;
 assign _5452 = ( _502 ) | ( _501 ) ;
 assign _5453 = ( _5451 ) | ( _5450 ) ;
 assign _5454 = ( _84 ) | ( n_n1156 ) ;
 assign _5455 = ( _5454 ) | ( _134 ) ;
 assign _5456 = ( n_n1125 ) | ( n_n1153 ) ;
 assign _5457 = ( _78 ) | ( n_n1121 ) ;
 assign _5458 = ( _163 ) | ( _85 ) ;
 assign _5459 = ( _5457 ) | ( _5456 ) ;
 assign _5460 = ( _265 ) | ( _164 ) ;
 assign _5461 = ( _5460 ) | ( _497 ) ;
 assign _5462 = ( _73 ) | ( n_n1254 ) ;
 assign _5463 = ( _182 ) | ( _174 ) ;
 assign _5464 = ( _276 ) | ( _188 ) ;
 assign _5465 = ( _116 ) | ( _489 ) ;
 assign _5466 = ( _5463 ) | ( _5462 ) ;
 assign _5467 = ( _5465 ) | ( _5464 ) ;
 assign _5468 = ( _109 ) | ( n_n1294 ) ;
 assign _5469 = ( _230 ) | ( _117 ) ;
 assign _5470 = ( _252 ) | ( _232 ) ;
 assign _5471 = ( _5469 ) | ( _5468 ) ;
 assign _5472 = ( n_n1286 ) | ( n_n1283 ) ;
 assign _5473 = ( _119 ) | ( _95 ) ;
 assign _5474 = ( _482 ) | ( _481 ) ;
 assign _5475 = ( _5473 ) | ( _5472 ) ;
 assign _5476 = ( _5475 ) | ( _5474 ) ;
 assign _5477 = ( _5476 ) | ( wire5315 ) ;
 assign _5478 = ( _186 ) | ( _160 ) ;
 assign _5479 = ( _275 ) | ( _191 ) ;
 assign _5480 = ( _476 ) | ( _475 ) ;
 assign _5481 = ( _5479 ) | ( _5478 ) ;
 assign _5482 = ( _198 ) | ( n_n1188 ) ;
 assign _5483 = ( _5482 ) | ( _273 ) ;
 assign _5484 = ( wire5306 ) | ( _5483 ) ;
 assign _5485 = ( n_n385 ) | ( n_n384 ) ;
 assign _5486 = ( n_n374 ) | ( _5484 ) ;
 assign _5487 = ( n_n1074 ) | ( n_n1055 ) ;
 assign _5488 = ( n_n1068 ) | ( n_n1077 ) ;
 assign _5489 = ( n_n1052 ) | ( n_n1047 ) ;
 assign _5490 = ( _5488 ) | ( _5487 ) ;
 assign _5491 = ( n_n421 ) | ( _5489 ) ;
 assign _5492 = ( n_n1088 ) | ( n_n1087 ) ;
 assign _5493 = ( _5492 ) | ( _111 ) ;
 assign _5494 = ( wire5324 ) | ( _5493 ) ;
 assign _5495 = ( n_n388 ) | ( n_n386 ) ;
 assign _5496 = ( _5495 ) | ( _5494 ) ;
 assign _5497 = ( n_n967 ) | ( n_n964 ) ;
 assign _5498 = ( _52 ) | ( n_n961 ) ;
 assign _5499 = ( _209 ) | ( _57 ) ;
 assign _5500 = ( _5498 ) | ( _5497 ) ;
 assign _5501 = ( n_n959 ) | ( n_n953 ) ;
 assign _5502 = ( _221 ) | ( _97 ) ;
 assign _5503 = ( n_n652 ) | ( _5501 ) ;
 assign _5504 = ( _5502 ) | ( n_n654 ) ;
 assign _5505 = ( _5503 ) | ( wire4934 ) ;
 assign _5506 = ( n_n395 ) | ( _5504 ) ;
 assign _5507 = ( n_n1032 ) | ( n_n1022 ) ;
 assign _5508 = ( n_n1026 ) | ( n_n1020 ) ;
 assign _5509 = ( _144 ) | ( _468 ) ;
 assign _5510 = ( _5507 ) | ( _212 ) ;
 assign _5511 = ( _5509 ) | ( _5508 ) ;
 assign _5512 = ( _315  &  _40 ) ;
 assign _5513 = ( n_n1045 ) | ( _153 ) ;
 assign _5514 = ( n_n1043 ) | ( n_n1046 ) ;
 assign _5515 = ( _217 ) | ( _461 ) ;
 assign _5516 = ( _5513 ) | ( _226 ) ;
 assign _5517 = ( _5515 ) | ( _5514 ) ;
 assign _5518 = ( n_n1011 ) | ( n_n1009 ) ;
 assign _5519 = ( n_n1013 ) | ( n_n1006 ) ;
 assign _5520 = ( _76 ) | ( n_n1010 ) ;
 assign _5521 = ( _5519 ) | ( _5518 ) ;
 assign _5522 = ( _329  &  i_1_ ) ;
 assign _5523 = ( n_n999 ) | ( _453 ) ;
 assign _5524 = ( n_n995 ) | ( n_n1004 ) ;
 assign _5525 = ( n_n993 ) | ( n_n994 ) ;
 assign _5526 = ( _454 ) | ( n_n1002 ) ;
 assign _5527 = ( _5524 ) | ( _5523 ) ;
 assign _5528 = ( _5526 ) | ( _5525 ) ;
 assign _5529 = ( n_n986 ) | ( n_n990 ) ;
 assign _5530 = ( n_n983 ) | ( n_n980 ) ;
 assign _5531 = ( _211 ) | ( n_n984 ) ;
 assign _5532 = ( _5529 ) | ( _255 ) ;
 assign _5533 = ( _5531 ) | ( _5530 ) ;
 assign _5534 = ( n_n977 ) | ( n_n974 ) ;
 assign _5535 = ( _264 ) | ( _99 ) ;
 assign _5536 = ( n_n365 ) | ( _5534 ) ;
 assign _5537 = ( _5536 ) | ( _5535 ) ;
 assign _5538 = ( n_n393 ) | ( n_n392 ) ;
 assign _5539 = ( _77 ) | ( n_n1014 ) ;
 assign _5540 = ( _5539 ) | ( _184 ) ;
 assign _5541 = ( wire5268 ) | ( _5540 ) ;
 assign _5542 = ( n_n389 ) | ( n_n390 ) ;
 assign _5543 = ( _5542 ) | ( _5541 ) ;
 assign _5544 = ( wire5290 ) | ( n_n379 ) ;
 assign _5545 = ( n_n1146 ) | ( n_n1147 ) ;
 assign _5546 = ( n_n1122 ) | ( n_n1145 ) ;
 assign _5547 = ( _161 ) | ( n_n1144 ) ;
 assign _5548 = ( _5546 ) | ( _5545 ) ;
 assign _5549 = ( n_n1018 ) | ( _196 ) ;
 assign _5550 = ( n_n1014 ) | ( n_n1010 ) ;
 assign _5551 = ( n_n1020 ) | ( n_n1019 ) ;
 assign _5552 = ( _219 ) | ( _62 ) ;
 assign _5553 = ( _5550 ) | ( _5549 ) ;
 assign _5554 = ( _5552 ) | ( _5551 ) ;
 assign _5555 = ( n_n1092 ) | ( n_n1060 ) ;
 assign _5556 = ( n_n1085 ) | ( n_n1074 ) ;
 assign _5557 = ( _257 ) | ( _75 ) ;
 assign _5558 = ( _5556 ) | ( _5555 ) ;
 assign _5559 = ( n_n1048 ) | ( n_n1045 ) ;
 assign _5560 = ( _5559 ) | ( _61 ) ;
 assign _5561 = ( n_n1120 ) | ( n_n1105 ) ;
 assign _5562 = ( _5561 ) | ( n_n1108 ) ;
 assign _5563 = ( wire5337 ) | ( _5562 ) ;
 assign _5564 = ( n_n204 ) | ( n_n205 ) ;
 assign _5565 = ( n_n1158 ) | ( n_n1169 ) ;
 assign _5566 = ( _148 ) | ( _84 ) ;
 assign _5567 = ( _218 ) | ( _149 ) ;
 assign _5568 = ( _5565 ) | ( _238 ) ;
 assign _5569 = ( _5567 ) | ( _5566 ) ;
 assign _5570 = ( n_n952 ) | ( n_n953 ) ;
 assign _5571 = ( n_n942 ) | ( n_n958 ) ;
 assign _5572 = ( _89 ) | ( _178 ) ;
 assign _5573 = ( _5570 ) | ( _222 ) ;
 assign _5574 = ( _5572 ) | ( _5571 ) ;
 assign _5575 = ( n_n994 ) | ( n_n991 ) ;
 assign _5576 = ( n_n980 ) | ( n_n974 ) ;
 assign _5577 = ( n_n984 ) | ( n_n981 ) ;
 assign _5578 = ( _98 ) | ( _58 ) ;
 assign _5579 = ( _5576 ) | ( _5575 ) ;
 assign _5580 = ( _5578 ) | ( _5577 ) ;
 assign _5581 = ( n_n967 ) | ( n_n964 ) ;
 assign _5582 = ( n_n970 ) | ( n_n971 ) ;
 assign _5583 = ( _5581 ) | ( _52 ) ;
 assign _5584 = ( _57 ) | ( n_n961 ) ;
 assign _5585 = ( wire5365 ) | ( _5584 ) ;
 assign _5586 = ( n_n206 ) | ( n_n208 ) ;
 assign _5587 = ( _180 ) | ( n_n1267 ) ;
 assign _5588 = ( _254 ) | ( _194 ) ;
 assign _5589 = ( _447 ) | ( _269 ) ;
 assign _5590 = ( _5588 ) | ( _5587 ) ;
 assign _5591 = ( n_n1177 ) | ( n_n1216 ) ;
 assign _5592 = ( _67 ) | ( n_n1174 ) ;
 assign _5593 = ( _198 ) | ( _142 ) ;
 assign _5594 = ( _236 ) | ( _216 ) ;
 assign _5595 = ( _5592 ) | ( _5591 ) ;
 assign _5596 = ( _5594 ) | ( _5593 ) ;
 assign _5597 = ( _197 ) | ( _173 ) ;
 assign _5598 = ( _5597 ) | ( _437 ) ;
 assign _5599 = ( wire5350 ) | ( _5598 ) ;
 assign _5600 = ( n_n201 ) | ( n_n202 ) ;
 assign _5601 = ( _5600 ) | ( _5599 ) ;
 assign _5602 = ( n_n196 ) | ( n_n195 ) ;
 assign _5603 = ( _108 ) | ( _82 ) ;
 assign _5604 = ( _430 ) | ( _228 ) ;
 assign _5605 = ( _165 ) | ( _431 ) ;
 assign _5606 = ( _5603 ) | ( _205 ) ;
 assign _5607 = ( _5605 ) | ( _5604 ) ;
 assign _5608 = ( n_n40  &  n_n75 ) ;
 assign _5609 = ( _113 ) | ( _83 ) ;
 assign _5610 = ( _159 ) | ( _151 ) ;
 assign _5611 = ( _424 ) | ( _237 ) ;
 assign _5612 = ( _5610 ) | ( _5609 ) ;
 assign _5613 = ( _158 ) | ( n_n1286 ) ;
 assign _5614 = ( _5613 ) | ( _249 ) ;
 assign _5615 = ( n_n58  &  _303 ) ;
 assign _5616 = ( _416 ) | ( _262 ) ;
 assign _5617 = ( _5616 ) | ( _86 ) ;
 assign _5618 = ( n_n198 ) | ( _5617 ) ;
 assign _5619 = ( _5618 ) | ( n_n199 ) ;
 assign _5620 = ( n_n1100 ) | ( n_n1092 ) ;
 assign _5621 = ( n_n1105 ) | ( n_n1088 ) ;
 assign _5622 = ( _115 ) | ( _114 ) ;
 assign _5623 = ( _136 ) | ( _155 ) ;
 assign _5624 = ( _5621 ) | ( _5620 ) ;
 assign _5625 = ( _5623 ) | ( _5622 ) ;
 assign _5626 = ( n_n78  &  i_2_ ) ;
 assign _5627 = ( n_n1128 ) | ( n_n1147 ) ;
 assign _5628 = ( _164 ) | ( _148 ) ;
 assign _5629 = ( _411 ) | ( _410 ) ;
 assign _5630 = ( _5628 ) | ( _5627 ) ;
 assign _5631 = ( n_n1120 ) | ( n_n1122 ) ;
 assign _5632 = ( _5631 ) | ( _103 ) ;
 assign _5633 = ( (~ i_0_)  &  (~ i_4_) ) ;
 assign _5634 = ( _5633  &  _26 ) ;
 assign _5635 = ( n_n1164 ) | ( _404 ) ;
 assign _5636 = ( _78 ) | ( n_n1156 ) ;
 assign _5637 = ( _154 ) | ( _149 ) ;
 assign _5638 = ( _5636 ) | ( _5635 ) ;
 assign _5639 = ( n_n1043 ) | ( _153 ) ;
 assign _5640 = ( _68 ) | ( n_n1048 ) ;
 assign _5641 = ( _212 ) | ( _195 ) ;
 assign _5642 = ( _5639 ) | ( _226 ) ;
 assign _5643 = ( _5641 ) | ( _5640 ) ;
 assign _5644 = ( n_n1068 ) | ( n_n1087 ) ;
 assign _5645 = ( n_n1057 ) | ( n_n1079 ) ;
 assign _5646 = ( _283 ) | ( _60 ) ;
 assign _5647 = ( _245 ) | ( _295 ) ;
 assign _5648 = ( _5645 ) | ( _5644 ) ;
 assign _5649 = ( _5647 ) | ( _5646 ) ;
 assign _5650 = ( _77 ) | ( n_n1014 ) ;
 assign _5651 = ( _219 ) | ( _144 ) ;
 assign _5652 = ( n_n295 ) | ( _5650 ) ;
 assign _5653 = ( _5652 ) | ( _5651 ) ;
 assign _5654 = ( n_n258 ) | ( n_n259 ) ;
 assign _5655 = ( n_n1184 ) | ( n_n1176 ) ;
 assign _5656 = ( _5655 ) | ( n_n1173 ) ;
 assign _5657 = ( wire5420 ) | ( _5656 ) ;
 assign _5658 = ( n_n256 ) | ( n_n257 ) ;
 assign _5659 = ( _5658 ) | ( _5657 ) ;
 assign _5660 = ( n_n953 ) | ( n_n969 ) ;
 assign _5661 = ( n_n962 ) | ( n_n958 ) ;
 assign _5662 = ( n_n966 ) | ( n_n970 ) ;
 assign _5663 = ( _5661 ) | ( _5660 ) ;
 assign _5664 = ( n_n974 ) | ( n_n975 ) ;
 assign _5665 = ( _5664 ) | ( n_n977 ) ;
 assign _5666 = ( n_n990 ) | ( n_n995 ) ;
 assign _5667 = ( n_n978 ) | ( n_n994 ) ;
 assign _5668 = ( _98 ) | ( _64 ) ;
 assign _5669 = ( _5666 ) | ( _255 ) ;
 assign _5670 = ( _5668 ) | ( _5667 ) ;
 assign _5671 = ( _96 ) | ( n_n944 ) ;
 assign _5672 = ( n_n654 ) | ( n_n652 ) ;
 assign _5673 = ( _5672 ) | ( _5671 ) ;
 assign _5674 = ( n_n261 ) | ( n_n262 ) ;
 assign _5675 = ( _5674 ) | ( _5673 ) ;
 assign _5676 = ( _246 ) | ( _223 ) ;
 assign _5677 = ( _284 ) | ( _277 ) ;
 assign _5678 = ( _399 ) | ( _398 ) ;
 assign _5679 = ( _5677 ) | ( _5676 ) ;
 assign _5680 = ( n_n1297 ) | ( n_n1294 ) ;
 assign _5681 = ( _113 ) | ( _110 ) ;
 assign _5682 = ( _237 ) | ( _157 ) ;
 assign _5683 = ( _5681 ) | ( _5680 ) ;
 assign _5684 = ( _158 ) | ( n_n1283 ) ;
 assign _5685 = ( _5684 ) | ( _159 ) ;
 assign _5686 = ( n_n1188 ) | ( n_n1193 ) ;
 assign _5687 = ( _142 ) | ( n_n1215 ) ;
 assign _5688 = ( _267 ) | ( _160 ) ;
 assign _5689 = ( _236 ) | ( _278 ) ;
 assign _5690 = ( _5687 ) | ( _5686 ) ;
 assign _5691 = ( _5689 ) | ( _5688 ) ;
 assign _5692 = ( _235 ) | ( _156 ) ;
 assign _5693 = ( _5692 ) | ( _392 ) ;
 assign _5694 = ( wire5389 ) | ( _5693 ) ;
 assign _5695 = ( n_n254 ) | ( n_n252 ) ;
 assign _5696 = ( _388 ) | ( _260 ) ;
 assign _5697 = ( _86 ) | ( _389 ) ;
 assign _5698 = ( _5696 ) | ( _387 ) ;
 assign _5699 = ( _121 ) | ( _109 ) ;
 assign _5700 = ( _291 ) | ( _263 ) ;
 assign _5701 = ( _382 ) | ( _381 ) ;
 assign _5702 = ( _5700 ) | ( _5699 ) ;
 assign _5703 = ( _271 ) | ( _248 ) ;
 assign _5704 = ( _5703 ) | ( _374 ) ;
 assign _5705 = ( n_n250 ) | ( _5704 ) ;
 assign _5706 = ( _5705 ) | ( wire5405 ) ;
 assign _5707 = ( n_n246 ) | ( _5706 ) ;


endmodule

