module k2 (
	Pz, Py, Px, Pw, Pv, Pu, Pt, Ps0, 
	Ps, Pr0, Pr, Pq0, Pq, Pp0, Pp, Po0, Po, Pn0, 
	Pn, Pm0, Pm, Pl0, Pl, Pk0, Pk, Pj0, Pj, Pi0, 
	Pi, Ph0, Ph, Pg0, Pg, Pf0, Pf, Pe0, Pe, Pd0, 
	Pd, Pc0, Pc, Pb0, Pb, Pa0, Pa, Pz1, Pz0, Py1, 
	Py0, Px1, Px0, Pw1, Pw0, Pv1, Pv0, Pu1, Pu0, Pt1, 
	Pt0, Ps1, Pr1, Pq1, Pp1, Po1, Pn1, Pm1, Pl2, Pl1, 
	Pk2, Pk1, Pj2, Pj1, Pi2, Pi1, Ph2, Ph1, Pg2, Pg1, 
	Pf2, Pf1, Pe2, Pe1, Pd2, Pd1, Pc2, Pc1, Pb2, Pb1, 
	Pa2, Pa1);

input Pz, Py, Px, Pw, Pv, Pu, Pt, Ps0, Ps, Pr0, Pr, Pq0, Pq, Pp0, Pp, Po0, Po, Pn0, Pn, Pm0, Pm, Pl0, Pl, Pk0, Pk, Pj0, Pj, Pi0, Pi, Ph0, Ph, Pg0, Pg, Pf0, Pf, Pe0, Pe, Pd0, Pd, Pc0, Pc, Pb0, Pb, Pa0, Pa;

output Pz1, Pz0, Py1, Py0, Px1, Px0, Pw1, Pw0, Pv1, Pv0, Pu1, Pu0, Pt1, Pt0, Ps1, Pr1, Pq1, Pp1, Po1, Pn1, Pm1, Pl2, Pl1, Pk2, Pk1, Pj2, Pj1, Pi2, Pi1, Ph2, Ph1, Pg2, Pg1, Pf2, Pf1, Pe2, Pe1, Pd2, Pd1, Pc2, Pc1, Pb2, Pb1, Pa2, Pa1;

wire n7, n8, n9, n10, n6, n12, n11, n14, n13, n15, n17, n18, n19, n20, n16, n22, n23, n24, n21, n26, n27, n25, n29, n30, n31, n28, n32, n34, n35, n33, n37, n38, n39, n40, n36, n42, n43, n44, n45, n41, n47, n48, n49, n46, n51, n52, n50, n54, n53, n57, n58, n56, n60, n61, n62, n59, n66, n67, n68, n69, n70, n63, n72, n73, n74, n75, n71, n77, n78, n79, n80, n81, n76, n83, n84, n85, n86, n87, n88, n89, n82, n91, n92, n93, n90, n95, n96, n97, n98, n99, n100, n101, n94, n103, n104, n105, n106, n108, n102, n110, n111, n112, n109, n114, n115, n116, n117, n118, n119, n113, n121, n122, n123, n124, n120, n126, n127, n128, n125, n130, n131, n132, n133, n134, n129, n136, n135, n138, n139, n137, n141, n140, n143, n144, n146, n147, n148, n149, n142, n151, n152, n153, n154, n155, n150, n158, n156, n160, n161, n162, n159, n165, n166, n167, n168, n170, n169, n173, n176, n180, n187, n184, n190, n191, n192, n188, n194, n193, n196, n197, n198, n199, n200, n201, n195, n203, n202, n205, n204, n210, n207, n211, n214, n213, n217, n218, n219, n221, n222, n226, n225, n223, n228, n227, n232, n233, n235, n236, n234, n239, n238, n237, n240, n241, n242, n245, n243, n246, n247, n251, n250, n248, n252, n255, n256, n257, n258, n259, n262, n263, n264, n266, n267, n269, n271, n277, n274, n275, n273, n279, n280, n281, n282, n278, n283, n286, n284, n288, n287, n290, n291, n289, n293, n292, n302, n299, n304, n303, n307, n306, n305, n308, n312, n311, n314, n313, n319, n317, n318, n320, n321, n323, n326, n327, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n349, n351, n353, n354, n355, n356, n357, n359, n360, n361, n362, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n377, n379, n380, n381, n383, n384, n385, n386, n387, n388, n390, n391, n392, n393, n394, n395, n397, n398, n399, n400, n401, n403, n402, n405, n406, n404, n407, n410, n414, n415, n418, n417, n419, n421, n422, n423, n425, n426, n428, n438, n446;

assign Pz1 = ( (~ n414) ) ;
 assign Pz0 = ( (~ n56) ) ;
 assign Py1 = ( (~ n36) ) ;
 assign Py0 = ( (~ n16) ) ;
 assign Px1 = ( (~ n33) ) ;
 assign Px0 = ( (~ n8) ) ;
 assign Pw1 = ( (~ n140) ) ;
 assign Pw0 = ( (~ n13) ) ;
 assign Pv1 = ( (~ n137) ) ;
 assign Pv0 =((~ Pz) & Pz);
 assign Pu1 = ( (~ n135) ) ;
 assign Pu0 = ( (~ n11) ) ;
 assign Pt1 = ( (~ n234) ) ;
 assign Pt0 = ( (~ n6) ) ;
 assign Ps1 = ( (~ n129) ) ;
 assign Pr1 = ( (~ n52) ) ;
 assign Pq1 = ( (~ n32) ) ;
 assign Pp1 = ( (~ n125) ) ;
 assign Po1 = ( (~ n256) ) ;
 assign Pn1 = ( (~ n257) ) ;
 assign Pm1 = ( (~ n120) ) ;
 assign Pl2 = ( (~ n52) ) ;
 assign Pl1 = ( (~ n113) ) ;
 assign Pk2 = ( (~ n50) ) ;
 assign Pk1 = ( (~ n109) ) ;
 assign Pj2 =((~ Pz) & Pz);
 assign Pj1 = ( (~ n102) ) ;
 assign Pi2 = ( (~ n351) ) ;
 assign Pi1 = ( (~ n94) ) ;
 assign Ph2 = ( (~ n46) ) ;
 assign Ph1 = ( (~ n90) ) ;
 assign Pg2 = ( (~ n100) ) ;
 assign Pg1 = ( (~ n82) ) ;
 assign Pf2 = ( (~ n7) ) | ( (~ n11) ) | ( (~ n40) ) | ( n165 ) | ( n166 ) ;
 assign Pf1 = ( (~ n76) ) ;
 assign Pe2 = ( (~ n159) ) ;
 assign Pe1 = ( (~ n71) ) ;
 assign Pd2 = ( (~ n156) ) ;
 assign Pd1 = ( (~ n63) ) ;
 assign Pc2 = ( (~ n150) ) ;
 assign Pc1 = ( (~ n28) ) ;
 assign Pb2 = ( (~ n142) ) ;
 assign Pb1 = ( (~ n59) ) ;
 assign Pa2 = ( (~ n41) ) ;
 assign Pa1 = ( (~ n21) ) ;
 assign n7 = ( Pa ) | ( n332 ) | ( n345 ) ;
 assign n8 = ( n15  &  n14  &  n12 ) ;
 assign n9 = ( (~ Py) ) | ( Pa ) | ( n286 ) ;
 assign n10 = ( n201 ) | ( (~ n339) ) ;
 assign n6 = ( n7  &  n8  &  n9  &  n10 ) ;
 assign n12 = ( (~ Py) ) | ( Pd0 ) | ( Pa ) | ( n217 ) ;
 assign n11 = ( n12  &  n9 ) ;
 assign n14 = ( (~ Pa0) ) | ( n201 ) ;
 assign n13 = ( n14  &  n10 ) ;
 assign n15 = ( (~ Py) ) | ( n201 ) ;
 assign n17 = ( (~ Pa) ) | ( n332 ) | ( n345 ) ;
 assign n18 = ( Pd0 ) | ( (~ Pa) ) | ( n217 ) ;
 assign n19 = ( (~ Py) ) | ( n344 ) ;
 assign n20 = ( n329 ) | ( n331 ) | ( n361 ) ;
 assign n16 = ( n17  &  n18  &  n19  &  n20 ) ;
 assign n22 = ( (~ n339) ) | ( n344 ) ;
 assign n23 = ( n200 ) | ( (~ n339) ) ;
 assign n24 = ( n27 ) | ( (~ n339) ) ;
 assign n21 = ( n22  &  n23  &  n24 ) ;
 assign n26 = ( Pl ) | ( (~ n339) ) ;
 assign n27 = ( (~ Pa) ) | ( (~ n205) ) | ( n240 ) ;
 assign n25 = ( n26 ) | ( n27 ) ;
 assign n29 = ( n332 ) | ( n302 ) | ( n330 ) | ( n331 ) ;
 assign n30 = ( (~ Pa) ) | ( n336 ) | ( n337 ) ;
 assign n31 = ( (~ Pd) ) | ( (~ Pa) ) | ( n320 ) | ( (~ n338) ) ;
 assign n28 = ( n29  &  n30  &  n31 ) ;
 assign n32 = ( n251  &  n250 ) | ( (~ n187)  &  n251  &  n248 ) ;
 assign n34 = ( (~ Pa) ) | ( n241 ) | ( n337 ) ;
 assign n35 = ( n354  &  n40  &  n25  &  n39 ) ;
 assign n33 = ( n24  &  n34  &  n35 ) ;
 assign n37 = ( n331 ) | ( n341 ) ;
 assign n38 = ( n331 ) | ( n342 ) ;
 assign n39 = ( n331 ) | ( n192 ) ;
 assign n40 = ( Pa ) | ( Pe ) | ( n353 ) ;
 assign n36 = ( n37  &  n38  &  n39  &  n40 ) ;
 assign n42 = ( (~ Pf) ) | ( Pc0 ) | ( n288 ) ;
 assign n43 = ( (~ Pe) ) | ( n353 ) ;
 assign n44 = ( (~ Pc0) ) | ( n288 ) ;
 assign n45 = ( n329 ) | ( (~ n338) ) ;
 assign n41 = ( n31  &  n42  &  n43  &  n44  &  n45 ) ;
 assign n47 = ( (~ Pf) ) | ( Pc0 ) | ( n192 ) ;
 assign n48 = ( (~ Pf)  &  n196 ) | ( (~ Pf)  &  n218 ) | ( n196  &  n219 ) | ( n218  &  n219 ) ;
 assign n49 = ( n42  &  n227 ) | ( n42  &  (~ n307) ) ;
 assign n46 = ( n47  &  n48  &  n49 ) ;
 assign n51 = ( (~ Py) ) | ( n222 ) ;
 assign n52 = ( (~ Pw) ) | ( n222 ) ;
 assign n50 = ( n51  &  n52 ) ;
 assign n54 = ( n343 ) | ( n369 ) ;
 assign n53 = ( (~ Pa0) ) | ( n54 ) ;
 assign n57 = ( Pc0 ) | ( n288 ) | ( n191 ) ;
 assign n58 = ( n38  &  n59  &  n141  &  n24  &  n34  &  n37 ) ;
 assign n56 = ( n28  &  n57  &  n58 ) ;
 assign n60 = ( n232  &  n160  &  n355  &  n356 ) ;
 assign n61 = ( n342 ) | ( n331 ) | ( Pl ) ;
 assign n62 = ( (~ Pl) ) | ( n331 ) | ( n341 ) ;
 assign n59 = ( n35  &  n60  &  n61  &  n62 ) ;
 assign n66 = ( (~ Pm0) ) | ( n370 ) ;
 assign n67 = ( (~ Pq0) ) | ( Pn0 ) | ( n371 ) ;
 assign n68 = ( n106  &  n73  &  n84  &  n53  &  n391  &  n377 ) ;
 assign n69 = ( n151  &  n86  &  n32  &  n101 ) ;
 assign n70 = ( n397  &  n77 ) ;
 assign n63 = ( n66  &  n67  &  n68  &  n69  &  n70  &  (~ n169)  &  (~ n438) ) ;
 assign n72 = ( Pd ) | ( n320 ) | ( (~ n338) ) ;
 assign n73 = ( (~ Px) ) | ( (~ Pb) ) | ( n238 ) | ( n293 ) ;
 assign n74 = ( n32  &  n101  &  n144 ) ;
 assign n75 = ( n138  &  (~ n169)  &  n375  &  n402  &  n404 ) ;
 assign n71 = ( n72  &  n73  &  n70  &  n74  &  n75 ) ;
 assign n77 = ( n45  &  n95  &  n168  &  (~ n395) ) ;
 assign n78 = ( n44  &  n390  &  n167 ) ;
 assign n79 = ( Pr0 ) | ( n372 ) ;
 assign n80 = ( (~ Pd0)  &  n199 ) | ( n199  &  n217 ) | ( (~ Pd0)  &  (~ n339) ) | ( n217  &  (~ n339) ) ;
 assign n81 = ( (~ Pa0) ) | ( n199 ) ;
 assign n76 = ( n77  &  n75  &  n78  &  n69  &  n79  &  n80  &  n72  &  n81 ) ;
 assign n83 = ( n116  &  (~ n176) ) ;
 assign n84 = ( n143  &  n78 ) ;
 assign n85 = ( (~ Pn) ) | ( n262 ) | ( n321 ) ;
 assign n86 = ( (~ Ps0) ) | ( Pr0 ) | ( Po0 ) | ( n267 ) ;
 assign n87 = ( n72  &  (~ n173)  &  n392  &  n393 ) ;
 assign n88 = ( n67  &  n131  &  n394  &  (~ n438) ) ;
 assign n89 = ( n123  &  n132  &  n81  &  n80  &  n400 ) ;
 assign n82 = ( n83  &  n84  &  n85  &  n86  &  n87  &  n88  &  n89 ) ;
 assign n91 = ( (~ Po0)  &  (~ Ph0) ) | ( (~ Po0)  &  n266 ) | ( (~ Ph0)  &  n267 ) | ( n266  &  n267 ) ;
 assign n92 = ( (~ Pc0) ) | ( n280 ) | ( n361 ) ;
 assign n93 = ( n349 ) | ( n280 ) ;
 assign n90 = ( n91  &  n68  &  n87  &  n92  &  n81  &  n93 ) ;
 assign n95 = ( n194  &  n283  &  Pc0 ) | ( n194  &  n283  &  n278 ) ;
 assign n96 = ( n118  &  n124  &  n144  &  (~ n176)  &  n383  &  n390  &  n399  &  n407 ) ;
 assign n97 = ( n373  &  n213  &  n121  &  n114 ) ;
 assign n98 = ( n31  &  n29  &  n232  &  n233 ) ;
 assign n99 = ( (~ n274) ) | ( n304 ) | ( (~ n306) ) ;
 assign n100 = ( n47  &  n136  &  n152  &  n167  &  n168  &  (~ n169) ) ;
 assign n101 = ( n326 ) | ( n304 ) ;
 assign n94 = ( n95  &  n96  &  n97  &  n98  &  n99  &  n100  &  n17  &  n101 ) ;
 assign n103 = ( n88  &  n69  &  n66  &  n135  &  n398  &  n130  &  n132  &  n399 ) ;
 assign n104 = ( n52  &  n401  &  n87 ) ;
 assign n105 = ( n237  &  n241 ) | ( n240  &  n241 ) | ( n237  &  n242 ) | ( n240  &  n242 ) ;
 assign n106 = ( (~ Pp0) ) | ( Pm0 ) | ( n370 ) ;
 assign n108 = ( Pc0 ) | ( n326 ) | ( n329 ) ;
 assign n102 = ( n84  &  n85  &  n103  &  n104  &  n105  &  n106  &  n108  &  (~ n176) ) ;
 assign n110 = ( n115  &  n211  &  n374  &  n79 ) ;
 assign n111 = ( n255  &  n256  &  n257  &  n258 ) ;
 assign n112 = ( (~ n173)  &  n251  &  n398 ) ;
 assign n109 = ( n91  &  n77  &  n89  &  n96  &  n75  &  n110  &  n111  &  n112 ) ;
 assign n114 = ( (~ Pi0) ) | ( n366 ) ;
 assign n115 = ( (~ Pk0) ) | ( n367 ) ;
 assign n116 = ( n243  &  n105  &  n234  &  n383 ) ;
 assign n117 = ( n17  &  n77  &  (~ n169)  &  n373  &  n386  &  n399  &  n400 ) ;
 assign n118 = ( n85  &  n379  &  n51  &  n394 ) ;
 assign n119 = ( n374  &  n387  &  n131  &  n132  &  n203  &  n72 ) ;
 assign n113 = ( n114  &  n115  &  n116  &  n117  &  n118  &  n119 ) ;
 assign n121 = ( (~ Pg0) ) | ( Pf0 ) | ( n214 ) ;
 assign n122 = ( (~ Ph0) ) | ( n365 ) ;
 assign n123 = ( (~ Px) ) | ( (~ Pu) ) | ( n368 ) ;
 assign n124 = ( (~ Pw) ) | ( (~ Pe0) ) | ( (~ Pc0) ) | ( (~ n306) ) | ( n343 ) ;
 assign n120 = ( n104  &  n117  &  n83  &  n74  &  n121  &  n122  &  n123  &  n124 ) ;
 assign n126 = ( n375  &  n133  &  n97  &  n110  &  n122  &  n80  &  n379  &  n380 ) ;
 assign n127 = ( n123  &  n50  &  n246  &  n247 ) ;
 assign n128 = ( n405  &  n403  &  n144  &  n17  &  n406  &  n99 ) ;
 assign n125 = ( n90  &  n126  &  n127  &  n70  &  n103  &  n128 ) ;
 assign n130 = ( (~ n275) ) | ( n329 ) | ( n336 ) ;
 assign n131 = ( (~ Pa0) ) | ( (~ n275) ) | ( n329 ) | ( n335 ) ;
 assign n132 = ( (~ Pw) ) | ( (~ Pu) ) | ( n368 ) ;
 assign n133 = ( n203  &  n195 ) | ( n203  &  n202 ) ;
 assign n134 = ( (~ Pw)  &  (~ Pa0) ) | ( (~ Pa0)  &  n221 ) | ( (~ Pw)  &  n222 ) | ( n221  &  n222 ) ;
 assign n129 = ( n130  &  n131  &  n132  &  n85  &  n133  &  n134  &  n127 ) ;
 assign n136 = ( n330 ) | ( n381 ) ;
 assign n135 = ( n136  &  n98  &  n43  &  n47 ) ;
 assign n138 = ( n92  &  n377 ) ;
 assign n139 = ( n48  &  n134  &  (~ n223)  &  n367 ) ;
 assign n137 = ( n52  &  n81  &  n138  &  n139  &  n126 ) ;
 assign n141 = ( n22  &  n23  &  n359  &  n360  &  n193 ) ;
 assign n140 = ( n16  &  n28  &  n57  &  n60  &  n141 ) ;
 assign n143 = ( (~ n259)  &  n262 ) | ( (~ n259)  &  n263 ) | ( (~ n259)  &  n264 ) ;
 assign n144 = ( (~ Pr0) ) | ( n372 ) ;
 assign n146 = ( n20  &  n36  &  n410  &  n57  &  n266 ) ;
 assign n147 = ( n91  &  n402  &  n101  &  n99 ) ;
 assign n148 = ( n404  &  n303 ) ;
 assign n149 = ( n67  &  n86  &  n66  &  n106  &  n168  &  n232  &  n29  &  n418 ) ;
 assign n142 = ( n95  &  n143  &  n144  &  n146  &  n147  &  n148  &  n149  &  (~ n173) ) ;
 assign n151 = ( Pj ) | ( n388 ) ;
 assign n152 = ( n32  &  n43  &  n45  &  n73  &  (~ n395)  &  n397 ) ;
 assign n153 = ( n319  &  Pg ) | ( n319  &  n317  &  n318 ) ;
 assign n154 = ( n72  &  n255  &  n398  &  (~ n438) ) ;
 assign n155 = ( n410  &  n390  &  n51  &  n246  &  n30  &  n42  &  n16  &  n29 ) ;
 assign n150 = ( n58  &  n83  &  n151  &  n152  &  n153  &  n154  &  n155  &  (~ n173) ) ;
 assign n158 = ( n30  &  n193  &  n303  &  (~ n308)  &  (~ n311)  &  (~ n313)  &  n355  &  n414 ) ;
 assign n156 = ( n31  &  n32  &  n33  &  n147  &  n154  &  n158  &  (~ n395) ) ;
 assign n160 = ( (~ n184)  &  n351 ) ;
 assign n161 = ( (~ Pa0) ) | ( n217 ) ;
 assign n162 = ( n360  &  n125  &  n354  &  n359  &  n21  &  n34  &  n19  &  n18 ) ;
 assign n159 = ( n139  &  n146  &  n153  &  n158  &  n160  &  n161  &  n162  &  (~ n169) ) ;
 assign n165 = ( Px  &  (~ Pb)  &  (~ n292) ) | ( Pw  &  (~ Pb)  &  (~ n292) ) ;
 assign n166 = ( (~ Pa)  &  (~ n415) ) | ( (~ Pa)  &  (~ n425) ) | ( (~ Pa)  &  (~ n426) ) ;
 assign n167 = ( n386  &  n387  &  n111 ) ;
 assign n168 = ( n335 ) | ( n369 ) ;
 assign n170 = ( (~ Pt)  &  (~ Ps)  &  n205 ) ;
 assign n169 = ( Pc0  &  (~ n364) ) | ( (~ Pv)  &  Pc0  &  n170 ) ;
 assign n173 = ( Pd  &  (~ n381) ) | ( (~ Pc)  &  (~ n381) ) ;
 assign n176 = ( (~ Pc0)  &  (~ n342) ) | ( Pr  &  (~ Pc0)  &  (~ n341) ) ;
 assign n180 = ( (~ Ph0)  &  (~ Pf0)  &  (~ n266) ) ;
 assign n187 = ( (~ Pl)  &  Pa0 ) ;
 assign n184 = ( Pw  &  (~ n200) ) | ( n187  &  (~ n200) ) | ( Pw  &  (~ n344) ) | ( n187  &  (~ n344) ) ;
 assign n190 = ( (~ n205) ) | ( n281 ) ;
 assign n191 = ( Pf ) | ( (~ Pa) ) ;
 assign n192 = ( (~ n277) ) | ( n279 ) ;
 assign n188 = ( (~ Pa)  &  n191 ) | ( n190  &  n191 ) | ( (~ Pa)  &  n192 ) | ( n190  &  n192 ) ;
 assign n194 = ( (~ Pr) ) | ( Pc0 ) | ( n357 ) ;
 assign n193 = ( Pc0  &  (~ Pa) ) | ( (~ Pa)  &  n188 ) | ( Pc0  &  n194 ) | ( n188  &  n194 ) ;
 assign n196 = ( (~ Pf) ) | ( n290 ) ;
 assign n197 = ( Pu ) | ( n368 ) ;
 assign n198 = ( (~ n333) ) | ( n343 ) ;
 assign n199 = ( Pu ) | ( n362 ) ;
 assign n200 = ( Pp ) | ( n191 ) | ( n290 ) ;
 assign n201 = ( n329 ) | ( n293 ) ;
 assign n195 = ( n196  &  n197  &  n198  &  n199  &  n200  &  n201 ) ;
 assign n203 = ( n197 ) | ( (~ n339) ) ;
 assign n202 = ( (~ Pz) ) | ( Pk ) ;
 assign n205 = ( (~ Pu)  &  n277 ) ;
 assign n204 = ( Px  &  n205  &  (~ n293) ) | ( Pw  &  n205  &  (~ n293) ) ;
 assign n210 = ( n345 ) | ( n369 ) ;
 assign n207 = ( (~ Pz) ) | ( (~ Pl) ) | ( n210 ) ;
 assign n211 = ( (~ Pw) ) | ( n199 ) ;
 assign n214 = ( (~ Px) ) | ( (~ Pv) ) | ( (~ n170) ) ;
 assign n213 = ( (~ Pf0) ) | ( n214 ) ;
 assign n217 = ( (~ Pu) ) | ( n362 ) ;
 assign n218 = ( Pz  &  (~ n339) ) ;
 assign n219 = ( n329 ) | ( n349 ) ;
 assign n221 = ( n217  &  n197 ) ;
 assign n222 = ( n302 ) | ( n242 ) ;
 assign n226 = ( Pq  &  Pi ) | ( (~ Pq)  &  Ph ) | ( Pi  &  Ph ) ;
 assign n225 = ( Pc0  &  n333  &  n274 ) ;
 assign n223 = ( n226  &  n225 ) | ( n226  &  (~ n446) ) ;
 assign n228 = ( Pd ) | ( (~ n170) ) ;
 assign n227 = ( (~ Pf)  &  (~ Pd) ) | ( (~ Pf)  &  (~ n170) ) | ( (~ Pd)  &  n228 ) | ( (~ n170)  &  n228 ) ;
 assign n232 = ( (~ Pa) ) | ( n318 ) ;
 assign n233 = ( (~ Pg)  &  n49 ) | ( n49  &  n317  &  n318 ) ;
 assign n235 = ( Pc0 ) | ( n329 ) | ( n279 ) ;
 assign n236 = ( n336  &  n332 ) | ( n242  &  n332 ) | ( n336  &  n335 ) | ( n242  &  n335 ) ;
 assign n234 = ( n235  &  n108  &  n236 ) ;
 assign n239 = ( (~ Pw) ) | ( n238 ) ;
 assign n238 = ( Pu ) | ( n329 ) ;
 assign n237 = ( n239  &  n238 ) | ( n239  &  (~ n339) ) ;
 assign n240 = ( (~ Pt) ) | ( n323 ) ;
 assign n241 = ( Pc0 ) | ( Pr ) | ( n340 ) ;
 assign n242 = ( n329 ) | ( (~ n333) ) ;
 assign n245 = ( (~ Pt) ) | ( n302 ) ;
 assign n243 = ( (~ Px) ) | ( n238 ) | ( n245 ) ;
 assign n246 = ( (~ Px) ) | ( n332 ) | ( n343 ) ;
 assign n247 = ( n83  &  n240 ) | ( n83  &  n238 ) | ( n83  &  n202 ) ;
 assign n251 = ( (~ Pa0) ) | ( n384 ) ;
 assign n250 = ( n337 ) | ( n345 ) ;
 assign n248 = ( (~ Pl) ) | ( (~ Pa0) ) ;
 assign n252 = ( Pz  &  (~ n240)  &  (~ n282) ) | ( Pw  &  (~ n240)  &  (~ n282) ) ;
 assign n255 = ( (~ Pz) ) | ( (~ Pl) ) | ( n250 ) ;
 assign n256 = ( (~ Pc0) ) | ( n357 ) ;
 assign n257 = ( n241 ) | ( n369 ) ;
 assign n258 = ( (~ Pc0)  &  (~ n252) ) | ( n190  &  (~ n252) ) ;
 assign n259 = ( Pn0  &  n180 ) | ( (~ Pq0)  &  Pn0  &  (~ n371) ) ;
 assign n262 = ( (~ Pv) ) | ( Pc0 ) ;
 assign n263 = ( (~ Pw) ) | ( Ps ) ;
 assign n264 = ( Pt ) | ( n282 ) ;
 assign n266 = ( (~ Pj) ) | ( n388 ) ;
 assign n267 = ( Pn0 ) | ( Pq0 ) | ( n371 ) ;
 assign n269 = ( Py  &  (~ n384) ) | ( (~ Pa0)  &  (~ n384) ) ;
 assign n271 = ( Pw  &  (~ n250) ) | ( Pz  &  (~ Pl)  &  (~ n250) ) ;
 assign n277 = ( (~ Pe0)  &  Pd0 ) ;
 assign n274 = ( Pv  &  Ps ) ;
 assign n275 = ( Pt  &  Pu ) ;
 assign n273 = ( n277  &  (~ n349) ) | ( n277  &  n274  &  n275 ) ;
 assign n279 = ( Pv ) | ( n347 ) ;
 assign n280 = ( (~ Pe0) ) | ( (~ Pd0) ) ;
 assign n281 = ( (~ Pa0) ) | ( n240 ) ;
 assign n282 = ( Pu ) | ( n280 ) ;
 assign n278 = ( n279  &  n281 ) | ( n280  &  n281 ) | ( n279  &  n282 ) | ( n280  &  n282 ) ;
 assign n283 = ( n335 ) | ( n264 ) ;
 assign n286 = ( n242 ) | ( n343 ) ;
 assign n284 = ( (~ n205)  &  n286 ) | ( n240  &  n286 ) ;
 assign n288 = ( (~ Pe0) ) | ( n327 ) ;
 assign n287 = ( n288  &  Pv ) | ( n288  &  n228 ) ;
 assign n290 = ( n242 ) | ( n345 ) ;
 assign n291 = ( (~ Pw) ) | ( (~ Pu) ) | ( n329 ) | ( n343 ) ;
 assign n289 = ( n192  &  Pp ) | ( n192  &  n290  &  n291 ) ;
 assign n293 = ( (~ Pt) ) | ( Ps ) | ( n262 ) ;
 assign n292 = ( (~ n205)  &  n238 ) | ( n238  &  n245 ) | ( (~ n205)  &  n293 ) | ( n245  &  n293 ) ;
 assign n302 = ( Ps ) | ( Pv ) ;
 assign n299 = ( n279  &  n302 ) | ( n279  &  (~ n306)  &  (~ n333) ) ;
 assign n304 = ( (~ Pc0) ) | ( n320 ) ;
 assign n303 = ( n13  &  n15  &  n299 ) | ( n13  &  n15  &  n304 ) ;
 assign n307 = ( (~ Pv)  &  (~ Pc0) ) ;
 assign n306 = ( (~ Pu)  &  (~ Pt) ) ;
 assign n305 = ( n307  &  Pn ) | ( n307  &  n306  &  Ps ) ;
 assign n308 = ( Pp  &  (~ Pf)  &  (~ n219) ) | ( Pp  &  (~ Pf)  &  (~ n290) ) ;
 assign n312 = ( Pq  &  (~ Pi) ) | ( (~ Pq)  &  (~ Ph) ) | ( (~ Pi)  &  (~ Ph) ) ;
 assign n311 = ( n225  &  n312 ) | ( n312  &  (~ n446) ) ;
 assign n314 = ( (~ Px)  &  n333 ) ;
 assign n313 = ( n305  &  (~ n321) ) | ( n314  &  (~ n321)  &  (~ n335) ) ;
 assign n319 = ( n332 ) | ( n346 ) ;
 assign n317 = ( (~ Pd) ) | ( (~ Pc0) ) | ( n222 ) ;
 assign n318 = ( n242 ) | ( n346 ) ;
 assign n320 = ( Pd0 ) | ( Pe0 ) ;
 assign n321 = ( Pb0 ) | ( Po ) | ( n320 ) ;
 assign n323 = ( Pv ) | ( (~ Ps) ) ;
 assign n326 = ( (~ Pu) ) | ( Pb0 ) | ( n240 ) ;
 assign n327 = ( (~ Pd0) ) | ( n326 ) ;
 assign n329 = ( (~ Pe0) ) | ( Pd0 ) ;
 assign n330 = ( Pd ) | ( (~ Pc) ) ;
 assign n331 = ( (~ Pc0) ) | ( (~ Pa) ) ;
 assign n332 = ( Pt ) | ( n238 ) ;
 assign n333 = ( Pu  &  (~ Pt) ) ;
 assign n334 = ( (~ Pd0) ) | ( (~ n333) ) ;
 assign n335 = ( Pc0 ) | ( n302 ) ;
 assign n336 = ( (~ Px) ) | ( n335 ) ;
 assign n337 = ( Pe0 ) | ( n334 ) ;
 assign n338 = ( Pu  &  Pb0  &  (~ n240) ) ;
 assign n339 = ( Pk  &  Pz ) ;
 assign n340 = ( (~ Pa0) ) | ( n323 ) ;
 assign n341 = ( n340 ) | ( n242 ) ;
 assign n342 = ( n238 ) | ( n281 ) ;
 assign n343 = ( (~ Pv) ) | ( Ps ) ;
 assign n344 = ( (~ Pa) ) | ( n286 ) ;
 assign n345 = ( (~ Ps) ) | ( n262 ) ;
 assign n346 = ( Pd ) | ( (~ Pc0) ) | ( Pc ) | ( n302 ) ;
 assign n347 = ( n263 ) | ( (~ n275) ) ;
 assign n349 = ( n262 ) | ( n347 ) ;
 assign n351 = ( Pp ) | ( n191 ) | ( n219 ) ;
 assign n353 = ( Pe0 ) | ( (~ Pc0) ) | ( n327 ) ;
 assign n354 = ( (~ Pw) ) | ( n27 ) ;
 assign n355 = ( n191 ) | ( n228 ) | ( (~ n307) ) ;
 assign n356 = ( n26 ) | ( n200  &  n344 ) ;
 assign n357 = ( n337 ) | ( n340 ) ;
 assign n359 = ( n200 ) | ( n248 ) ;
 assign n360 = ( n344 ) | ( n248 ) ;
 assign n361 = ( (~ Pt) ) | ( n343 ) ;
 assign n362 = ( (~ Pt) ) | ( (~ Pe0) ) | ( (~ n274) ) ;
 assign n364 = ( n302 ) | ( n337 ) ;
 assign n365 = ( Pf0 ) | ( Pg0 ) | ( n214 ) ;
 assign n366 = ( Ph0 ) | ( n365 ) ;
 assign n367 = ( Pi0 ) | ( Pj0 ) | ( n366 ) ;
 assign n368 = ( Pt ) | ( (~ Pe0) ) | ( n323 ) ;
 assign n369 = ( (~ Pe0) ) | ( n334 ) ;
 assign n370 = ( (~ Pw) ) | ( Pj ) | ( (~ n170) ) | ( n262 ) ;
 assign n371 = ( Pm0 ) | ( Pp0 ) | ( n370 ) ;
 assign n372 = ( Ps0 ) | ( Po0 ) | ( n267 ) ;
 assign n373 = ( (~ Pj0) ) | ( Pi0 ) | ( n366 ) ;
 assign n374 = ( (~ Pc0) ) | ( (~ n274) ) | ( n332 ) ;
 assign n375 = ( n54  &  (~ n204)  &  n207 ) ;
 assign n377 = ( n248 ) | ( n210 ) ;
 assign n379 = ( (~ Pl0) ) | ( Pk0 ) | ( n367 ) ;
 assign n380 = ( n124  &  n401 ) ;
 assign n381 = ( (~ Pc0) ) | ( n279 ) | ( n329 ) ;
 assign n383 = ( n239 ) | ( n245 ) ;
 assign n384 = ( n337 ) | ( n343 ) ;
 assign n385 = ( (~ Pb) ) | ( (~ n205) ) | ( n245 ) ;
 assign n386 = ( (~ Px) ) | ( n385 ) ;
 assign n387 = ( (~ Pw) ) | ( n385 ) ;
 assign n388 = ( n262 ) | ( n332 ) | ( n263 ) ;
 assign n390 = ( (~ Pc0) ) | ( n279 ) | ( n280 ) ;
 assign n391 = ( (~ n187) ) | ( n210 ) ;
 assign n392 = ( (~ Pr) ) | ( n304 ) | ( (~ n333) ) | ( n340 ) ;
 assign n393 = ( Pu ) | ( n281 ) | ( n304 ) ;
 assign n394 = ( (~ Po) ) | ( Pc0 ) | ( Pb0 ) | ( n320 ) ;
 assign n395 = ( n269 ) | ( n271 ) | ( n273 ) | ( (~ n417) ) ;
 assign n397 = ( (~ Pb) ) | ( n239 ) | ( n293 ) ;
 assign n398 = ( Pc0 ) | ( Pe0 ) | ( n327 ) ;
 assign n399 = ( Pc0 ) | ( (~ n277) ) | ( (~ n338) ) ;
 assign n400 = ( n130  &  n397  &  n73 ) ;
 assign n401 = ( (~ Py) ) | ( n364 ) ;
 assign n403 = ( (~ Pz) ) | ( Pl ) | ( n210 ) ;
 assign n402 = ( n393  &  n403  &  n392 ) ;
 assign n405 = ( (~ Pw) ) | ( n210 ) ;
 assign n406 = ( n345 ) | ( n264 ) ;
 assign n404 = ( n405  &  n391  &  n93  &  n406 ) ;
 assign n407 = ( n44  &  n246 ) ;
 assign n410 = ( (~ Pc0) ) | ( n326 ) | ( n329 ) ;
 assign n414 = ( n321 ) | ( n262 ) | ( Pn ) | ( Pm ) ;
 assign n415 = ( (~ Pc0)  &  (~ n428) ) | ( n421  &  n422  &  (~ n428) ) ;
 assign n418 = ( (~ Pc0) ) | ( (~ n277) ) | ( n361 ) ;
 assign n417 = ( Pt  &  n418 ) | ( (~ n205)  &  n418 ) | ( n345  &  n418 ) ;
 assign n419 = ( (~ Px)  &  Pf ) | ( (~ Px)  &  n287 ) | ( Pf  &  n364 ) | ( n287  &  n364 ) ;
 assign n421 = ( n342  &  n192  &  n330 ) | ( n342  &  n192  &  n222 ) ;
 assign n422 = ( (~ Pl)  &  n329 ) | ( n329  &  n341 ) | ( (~ Pl)  &  n361 ) | ( n341  &  n361 ) ;
 assign n423 = ( Pd0  &  n319 ) | ( (~ Pd)  &  n319 ) | ( n319  &  (~ n338) ) ;
 assign n425 = ( n284  &  n423 ) | ( (~ Pz)  &  (~ Pw)  &  n423 ) ;
 assign n426 = ( Pf  &  (~ Pa0) ) | ( Pf  &  n286 ) | ( (~ Pa0)  &  n289 ) | ( n286  &  n289 ) ;
 assign n428 = ( (~ Pc0)  &  (~ n190) ) | ( (~ Pc0)  &  (~ n357) ) | ( (~ Pc0)  &  (~ n419) ) ;
 assign n438 = ( Pq0  &  Pn0  &  (~ n371) ) ;
 assign n446 = ( (~ Pv) ) | ( n304 ) | ( n347 ) ;


endmodule

