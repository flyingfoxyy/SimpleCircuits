module x4 (
	a, b, g, h, i, k, l, m, 
	n, o, p, q, r, s, t, u, v, w, 
	x, y, z, a0, b0, c0, d0, e0, f0, g0, 
	h0, i0, k0, l0, m0, n0, o0, p0, q0, r0, 
	s0, t0, u0, v0, w0, x0, y0, z0, a1, b1, 
	c1, d1, e1, f1, g1, h1, i1, j1, k1, l1, 
	m1, n1, o1, p1, q1, r1, s1, t1, u1, v1, 
	w1, x1, y1, z1, a2, b2, c2, d2, e2, f2, 
	g2, h2, i2, j2, k2, l2, m2, n2, o2, p2, 
	q2, r2, s2, t2, u2, v2, w2, x2, y2, z2, 
	a3, b3, c3, d3, e3, f3, g3, h3, i3, j3, 
	k3, l3, m3, n3, o3, p3, q3, r3, s3, t3, 
	u3, v3, w3, x3, y3, z3, a4, b4, c4, d4, 
	e4, f4, g4, h4, i4, j4, k4, l4, m4, n4, 
	o4, p4, q4, r4, s4, t4, u4, v4, w4, x4, 
	y4, z4, a5, b5, c5, d5, e5, f5, g5, h5, 
	i5, j5, k5, l5, m5, n5, o5);

input a, b, g, h, i, k, l, m, n, o, p, q, r, s, t, u, v, w, x, y, z, a0, b0, c0, d0, e0, f0, g0, h0, i0, k0, l0, m0, n0, o0, p0, q0, r0, s0, t0, u0, v0, w0, x0, y0, z0, a1, b1, c1, d1, e1, f1, g1, h1, i1, j1, k1, l1, m1, n1, o1, p1, q1, r1, s1, t1, u1, v1, w1, x1, y1, z1, a2, b2, c2, d2, e2, f2, g2, h2, i2, j2, k2, l2, m2, n2, o2, p2, q2, r2, s2, t2, u2, v2;

output w2, x2, y2, z2, a3, b3, c3, d3, e3, f3, g3, h3, i3, j3, k3, l3, m3, n3, o3, p3, q3, r3, s3, t3, u3, v3, w3, x3, y3, z3, a4, b4, c4, d4, e4, f4, g4, h4, i4, j4, k4, l4, m4, n4, o4, p4, q4, r4, s4, t4, u4, v4, w4, x4, y4, z4, a5, b5, c5, d5, e5, f5, g5, h5, i5, j5, k5, l5, m5, n5, o5;

wire j8, k8, m8, o8, w8, x8, f9, i9, k9, l9, d10, e10, f10, g10, l10, n10, u10, v10, x10, y10, z10, a11, c11, e11, f11, i11, j11, k11, l11, n11, q11, t11, w11, z11, c12, f12, i12, l12, o12, r12, u12, x12, a13, d13, g13, j13, m13, p13, u13, v13, w13, x13, y13, z13, a14, b14, c14, d14, e14, f14, g14, h14, j14, k14, l14;

assign w2 = ( (~ f1) ) ;
 assign x2 = ( (~ g1) ) ;
 assign y2 = ( (~ h1) ) ;
 assign z2 = ( (~ i1) ) ;
 assign a3 = ( (~ j1) ) ;
 assign b3 = ( (~ k1) ) ;
 assign c3 = ( (~ i0)  &  s2  &  (~ m8) ) | ( (~ i0)  &  e1  &  (~ j8)  &  (~ k8) ) ;
 assign d3 = ( (~ x8) ) | ( v2  &  (~ c1)  &  g0  &  (~ w8) ) ;
 assign e3 = ( (~ c1)  &  l0 ) | ( (~ c1)  &  e1  &  n2  &  (~ f9) ) ;
 assign f3 = ( (~ i9) ) | ( v2  &  g0  &  (~ w8) ) ;
 assign g3 = ( (~ c1)  &  (~ i0)  &  (~ k9) ) ;
 assign h3 = ( (~ c1)  &  o0  &  (~ i0) ) ;
 assign i3 = ( (~ c1)  &  p0  &  (~ i0) ) ;
 assign j3 = ( (~ c1)  &  q0  &  (~ i0) ) ;
 assign k3 = ( (~ c1)  &  r0  &  (~ i0) ) ;
 assign l3 = ( (~ c1)  &  s0  &  (~ i0) ) ;
 assign m3 = ( (~ c1)  &  t0  &  (~ i0) ) ;
 assign n3 = ( (~ i0)  &  b ) ;
 assign o3 = ( (~ i0)  &  a ) ;
 assign p3 = ( v0  &  (~ i0) ) ;
 assign q3 = ( w0  &  (~ i0) ) ;
 assign r3 = ( x0  &  (~ i0) ) ;
 assign s3 = ( y0  &  (~ i0) ) ;
 assign t3 = ( z0  &  (~ i0) ) ;
 assign u3 = ( a1  &  (~ i0) ) ;
 assign v3 = ( (~ f10) ) | ( v2  &  g0  &  (~ w8) ) | ( n2  &  e1  &  (~ d10)  &  (~ e10) ) ;
 assign w3 = ( v2  &  (~ g10) ) ;
 assign x3 = ( (~ c1)  &  e1 ) | ( (~ c1)  &  d1 ) | ( (~ c1)  &  (~ k2)  &  l2  &  m2 ) ;
 assign y3 = ( n2  &  f1  &  (~ c1) ) | ( (~ e1)  &  f1  &  (~ c1) ) | ( o0  &  f1  &  (~ c1) ) | ( (~ l10)  &  f1  &  (~ c1) ) | ( n2  &  (~ n10)  &  (~ c1) ) | ( (~ e1)  &  (~ n10)  &  (~ c1) ) | ( o0  &  (~ n10)  &  (~ c1) ) | ( (~ l10)  &  (~ n10)  &  (~ c1) ) ;
 assign z3 = ( n2  &  g1  &  (~ c1) ) | ( (~ e1)  &  g1  &  (~ c1) ) | ( p0  &  g1  &  (~ c1) ) | ( (~ l10)  &  g1  &  (~ c1) ) | ( n2  &  (~ n10)  &  (~ c1) ) | ( (~ e1)  &  (~ n10)  &  (~ c1) ) | ( p0  &  (~ n10)  &  (~ c1) ) | ( (~ l10)  &  (~ n10)  &  (~ c1) ) ;
 assign a4 = ( n2  &  h1  &  (~ c1) ) | ( (~ e1)  &  h1  &  (~ c1) ) | ( q0  &  h1  &  (~ c1) ) | ( (~ l10)  &  h1  &  (~ c1) ) | ( n2  &  (~ n10)  &  (~ c1) ) | ( (~ e1)  &  (~ n10)  &  (~ c1) ) | ( q0  &  (~ n10)  &  (~ c1) ) | ( (~ l10)  &  (~ n10)  &  (~ c1) ) ;
 assign b4 = ( n2  &  i1  &  (~ c1) ) | ( (~ e1)  &  i1  &  (~ c1) ) | ( r0  &  i1  &  (~ c1) ) | ( (~ l10)  &  i1  &  (~ c1) ) | ( n2  &  (~ n10)  &  (~ c1) ) | ( (~ e1)  &  (~ n10)  &  (~ c1) ) | ( r0  &  (~ n10)  &  (~ c1) ) | ( (~ l10)  &  (~ n10)  &  (~ c1) ) ;
 assign c4 = ( n2  &  j1  &  (~ c1) ) | ( (~ e1)  &  j1  &  (~ c1) ) | ( s0  &  j1  &  (~ c1) ) | ( (~ l10)  &  j1  &  (~ c1) ) | ( n2  &  (~ n10)  &  (~ c1) ) | ( (~ e1)  &  (~ n10)  &  (~ c1) ) | ( s0  &  (~ n10)  &  (~ c1) ) | ( (~ l10)  &  (~ n10)  &  (~ c1) ) ;
 assign d4 = ( n2  &  k1  &  (~ c1) ) | ( (~ e1)  &  k1  &  (~ c1) ) | ( t0  &  k1  &  (~ c1) ) | ( (~ l10)  &  k1  &  (~ c1) ) | ( n2  &  (~ n10)  &  (~ c1) ) | ( (~ e1)  &  (~ n10)  &  (~ c1) ) | ( t0  &  (~ n10)  &  (~ c1) ) | ( (~ l10)  &  (~ n10)  &  (~ c1) ) ;
 assign e4 = ( (~ c1)  &  l1 ) | ( (~ c1)  &  e1  &  n2  &  (~ f9) ) ;
 assign f4 = ( m1  &  (~ v10) ) | ( (~ u10)  &  (~ v10) ) ;
 assign g4 = ( (~ i0)  &  n1  &  (~ c11) ) | ( (~ i0)  &  (~ m0)  &  (~ y10)  &  (~ z10) ) | ( (~ i0)  &  g0  &  i  &  (~ a11) ) ;
 assign h4 = ( (~ f11) ) | ( v2  &  m1  &  g0  &  (~ e11) ) ;
 assign i4 = ( (~ i0)  &  p1  &  (~ l11) ) | ( g0  &  (~ e11)  &  k  &  (~ i11) ) | ( (~ i0)  &  (~ m0)  &  (~ j11)  &  (~ k11) ) ;
 assign j4 = ( (~ i0)  &  (~ l11)  &  q1 ) | ( g0  &  (~ e11)  &  (~ i11)  &  l ) | ( (~ i0)  &  (~ m0)  &  (~ k11)  &  (~ n11) ) ;
 assign k4 = ( (~ i0)  &  (~ l11)  &  r1 ) | ( g0  &  (~ e11)  &  (~ i11)  &  m ) | ( (~ i0)  &  (~ m0)  &  (~ k11)  &  (~ q11) ) ;
 assign l4 = ( (~ i0)  &  (~ l11)  &  s1 ) | ( g0  &  (~ e11)  &  (~ i11)  &  n ) | ( (~ i0)  &  (~ m0)  &  (~ k11)  &  (~ t11) ) ;
 assign m4 = ( (~ i0)  &  (~ l11)  &  t1 ) | ( g0  &  (~ e11)  &  (~ i11)  &  o ) | ( (~ i0)  &  (~ m0)  &  (~ k11)  &  (~ w11) ) ;
 assign n4 = ( (~ i0)  &  (~ l11)  &  u1 ) | ( g0  &  (~ e11)  &  (~ i11)  &  p ) | ( (~ i0)  &  (~ m0)  &  (~ k11)  &  (~ z11) ) ;
 assign o4 = ( (~ i0)  &  (~ l11)  &  v1 ) | ( g0  &  (~ e11)  &  (~ i11)  &  q ) | ( (~ i0)  &  (~ m0)  &  (~ k11)  &  (~ c12) ) ;
 assign p4 = ( (~ i0)  &  (~ l11)  &  w1 ) | ( g0  &  (~ e11)  &  (~ i11)  &  r ) | ( (~ i0)  &  (~ m0)  &  (~ k11)  &  (~ f12) ) ;
 assign q4 = ( (~ i0)  &  (~ l11)  &  x1 ) | ( g0  &  (~ e11)  &  (~ i11)  &  s ) | ( (~ i0)  &  (~ m0)  &  (~ k11)  &  (~ i12) ) ;
 assign r4 = ( (~ i0)  &  (~ l11)  &  y1 ) | ( g0  &  (~ e11)  &  (~ i11)  &  t ) | ( (~ i0)  &  (~ m0)  &  (~ k11)  &  (~ l12) ) ;
 assign s4 = ( (~ i0)  &  (~ l11)  &  z1 ) | ( g0  &  (~ e11)  &  (~ i11)  &  u ) | ( (~ i0)  &  (~ m0)  &  (~ k11)  &  (~ o12) ) ;
 assign t4 = ( (~ i0)  &  (~ l11)  &  a2 ) | ( g0  &  (~ e11)  &  (~ i11)  &  v ) | ( (~ i0)  &  (~ m0)  &  (~ k11)  &  (~ r12) ) ;
 assign u4 = ( (~ i0)  &  (~ l11)  &  b2 ) | ( g0  &  (~ e11)  &  (~ i11)  &  w ) | ( (~ i0)  &  (~ m0)  &  (~ k11)  &  (~ u12) ) ;
 assign v4 = ( (~ i0)  &  (~ l11)  &  c2 ) | ( g0  &  (~ e11)  &  (~ i11)  &  x ) | ( (~ i0)  &  (~ m0)  &  (~ k11)  &  (~ x12) ) ;
 assign w4 = ( (~ i0)  &  (~ l11)  &  d2 ) | ( g0  &  (~ e11)  &  (~ i11)  &  y ) | ( (~ i0)  &  (~ m0)  &  (~ k11)  &  (~ a13) ) ;
 assign x4 = ( (~ i0)  &  (~ l11)  &  e2 ) | ( g0  &  (~ e11)  &  (~ i11)  &  z ) | ( (~ i0)  &  (~ m0)  &  (~ k11)  &  (~ d13) ) ;
 assign y4 = ( (~ i0)  &  (~ l11)  &  f2 ) | ( g0  &  (~ e11)  &  (~ i11)  &  a0 ) | ( (~ i0)  &  (~ m0)  &  (~ k11)  &  (~ g13) ) ;
 assign z4 = ( (~ i0)  &  (~ l11)  &  g2 ) | ( g0  &  (~ e11)  &  (~ i11)  &  b0 ) | ( (~ i0)  &  (~ m0)  &  (~ k11)  &  (~ j13) ) ;
 assign a5 = ( (~ i0)  &  (~ l11)  &  h2 ) | ( g0  &  (~ e11)  &  (~ i11)  &  c0 ) | ( (~ i0)  &  (~ m0)  &  (~ k11)  &  (~ m13) ) ;
 assign b5 = ( (~ i0)  &  (~ l11)  &  i2 ) | ( g0  &  (~ e11)  &  (~ i11)  &  d0 ) | ( (~ i0)  &  (~ m0)  &  (~ k11)  &  (~ p13) ) ;
 assign c5 = ( j2  &  (~ i0)  &  (~ l11) ) | ( g0  &  e0  &  (~ i11)  &  (~ e11) ) ;
 assign d5 = ( u2  &  (~ v13) ) | ( k2  &  (~ v13) ) | ( (~ u13)  &  (~ v13) ) ;
 assign e5 = ( (~ k2)  &  l2  &  (~ x13) ) | ( (~ k2)  &  u2  &  (~ x13) ) | ( (~ l2)  &  u2  &  (~ x13) ) | ( (~ k2)  &  (~ u13)  &  (~ x13) ) | ( (~ l2)  &  (~ u13)  &  (~ x13) ) | ( l2  &  (~ w13)  &  (~ x13) ) | ( u2  &  (~ w13)  &  (~ x13) ) | ( (~ u13)  &  (~ w13)  &  (~ x13) ) ;
 assign f5 = ( (~ l2)  &  m2  &  (~ y13) ) | ( (~ l2)  &  u2  &  (~ y13) ) | ( (~ m2)  &  u2  &  (~ y13) ) | ( (~ l2)  &  (~ u13)  &  (~ y13) ) | ( (~ m2)  &  (~ u13)  &  (~ y13) ) | ( m2  &  (~ w13)  &  (~ y13) ) | ( u2  &  (~ w13)  &  (~ y13) ) | ( (~ u13)  &  (~ w13)  &  (~ y13) ) ;
 assign g5 = ( n2  &  (~ a14) ) | ( e1  &  (~ a14) ) | ( d1  &  (~ a14) ) | ( (~ z13)  &  (~ a14) ) ;
 assign h5 = ( (~ n2)  &  o2  &  (~ c14) ) | ( (~ n2)  &  e1  &  (~ c14) ) | ( (~ o2)  &  e1  &  (~ c14) ) | ( (~ n2)  &  d1  &  (~ c14) ) | ( (~ o2)  &  d1  &  (~ c14) ) | ( (~ n2)  &  (~ z13)  &  (~ c14) ) | ( (~ o2)  &  (~ z13)  &  (~ c14) ) | ( o2  &  (~ b14)  &  (~ c14) ) | ( e1  &  (~ b14)  &  (~ c14) ) | ( d1  &  (~ b14)  &  (~ c14) ) | ( (~ z13)  &  (~ b14)  &  (~ c14) ) ;
 assign i5 = ( (~ n2)  &  p2  &  (~ d14) ) | ( (~ o2)  &  p2  &  (~ d14) ) | ( (~ n2)  &  e1  &  (~ d14) ) | ( (~ o2)  &  e1  &  (~ d14) ) | ( (~ p2)  &  e1  &  (~ d14) ) | ( (~ n2)  &  d1  &  (~ d14) ) | ( (~ o2)  &  d1  &  (~ d14) ) | ( (~ p2)  &  d1  &  (~ d14) ) | ( (~ n2)  &  (~ z13)  &  (~ d14) ) | ( (~ o2)  &  (~ z13)  &  (~ d14) ) | ( (~ p2)  &  (~ z13)  &  (~ d14) ) | ( p2  &  (~ b14)  &  (~ d14) ) | ( e1  &  (~ b14)  &  (~ d14) ) | ( d1  &  (~ b14)  &  (~ d14) ) | ( (~ z13)  &  (~ b14)  &  (~ d14) ) ;
 assign j5 = ( (~ o2)  &  q2  &  (~ f14) ) | ( (~ n2)  &  q2  &  (~ f14) ) | ( (~ e14)  &  q2  &  (~ f14) ) | ( (~ b14)  &  q2  &  (~ f14) ) | ( (~ o2)  &  e1  &  (~ f14) ) | ( (~ n2)  &  e1  &  (~ f14) ) | ( (~ e14)  &  e1  &  (~ f14) ) | ( (~ b14)  &  e1  &  (~ f14) ) | ( (~ o2)  &  d1  &  (~ f14) ) | ( (~ n2)  &  d1  &  (~ f14) ) | ( (~ e14)  &  d1  &  (~ f14) ) | ( (~ b14)  &  d1  &  (~ f14) ) | ( (~ o2)  &  (~ z13)  &  (~ f14) ) | ( (~ n2)  &  (~ z13)  &  (~ f14) ) | ( (~ e14)  &  (~ z13)  &  (~ f14) ) | ( (~ b14)  &  (~ z13)  &  (~ f14) ) ;
 assign k5 = ( (~ n2)  &  r2  &  (~ c1) ) | ( (~ o2)  &  r2  &  (~ c1) ) | ( r2  &  (~ b14)  &  (~ c1) ) | ( r2  &  (~ g14)  &  (~ c1) ) | ( (~ n2)  &  e1  &  (~ h14)  &  (~ c1) ) | ( (~ o2)  &  e1  &  (~ h14)  &  (~ c1) ) | ( (~ n2)  &  d1  &  (~ h14)  &  (~ c1) ) | ( (~ o2)  &  d1  &  (~ h14)  &  (~ c1) ) | ( (~ n2)  &  (~ z13)  &  (~ h14)  &  (~ c1) ) | ( (~ o2)  &  (~ z13)  &  (~ h14)  &  (~ c1) ) | ( e1  &  (~ b14)  &  (~ h14)  &  (~ c1) ) | ( d1  &  (~ b14)  &  (~ h14)  &  (~ c1) ) | ( (~ z13)  &  (~ b14)  &  (~ h14)  &  (~ c1) ) | ( e1  &  (~ g14)  &  (~ h14)  &  (~ c1) ) | ( d1  &  (~ g14)  &  (~ h14)  &  (~ c1) ) | ( (~ z13)  &  (~ g14)  &  (~ h14)  &  (~ c1) ) ;
 assign l5 = ( (~ i0)  &  m0  &  b1 ) | ( (~ i0)  &  (~ e1)  &  b1 ) | ( (~ i0)  &  b1  &  n1 ) | ( (~ i0)  &  (~ m0)  &  e1  &  n1 ) ;
 assign m5 = ( (~ c1)  &  (~ l1)  &  t2 ) | ( (~ c1)  &  (~ s2)  &  t2 ) | ( (~ c1)  &  l1  &  s2  &  (~ t2) ) ;
 assign n5 = ( (~ m2)  &  (~ j14) ) | ( (~ l2)  &  (~ j14) ) | ( k2  &  (~ j14) ) | ( (~ u13)  &  (~ j14) ) ;
 assign o5 = ( (~ v10)  &  (~ k14) ) | ( (~ f0)  &  v2  &  (~ v10) ) ;
 assign j8 = ( (~ r2) ) | ( p2 ) | ( o2 ) | ( (~ n2) ) ;
 assign k8 = ( (~ i)  &  (~ q2) ) | ( (~ h0)  &  t2 ) | ( h0  &  (~ t2) ) ;
 assign m8 = ( (~ p2)  &  r2  &  (~ o8) ) ;
 assign o8 = ( (~ n2) ) | ( (~ e1) ) | ( o2 ) | ( (~ i)  &  (~ q2) ) ;
 assign w8 = ( g  &  m1 ) | ( h  &  m1 ) | ( i  &  m1 ) | ( (~ h0)  &  m1 ) ;
 assign x8 = ( c1 ) | ( (~ f0)  &  (~ k0) ) | ( (~ k0)  &  (~ v2) ) ;
 assign f9 = ( r2 ) | ( q2 ) | ( p2 ) | ( o2 ) ;
 assign i9 = ( (~ i0)  &  (~ m0) ) | ( (~ i0)  &  v2  &  g0 ) ;
 assign k9 = ( o2  &  (~ n0) ) | ( (~ n2)  &  (~ n0) ) | ( (~ e1)  &  (~ n0) ) | ( (~ l9)  &  (~ n0) ) ;
 assign l9 = ( (~ r2)  &  (~ q2)  &  (~ p2) ) ;
 assign d10 = ( (~ r2) ) | ( p2 ) | ( o2 ) ;
 assign e10 = ( (~ q2)  &  (~ i) ) ;
 assign f10 = ( (~ f0)  &  (~ i0) ) | ( (~ i0)  &  (~ v2) ) ;
 assign g10 = ( (~ i0) ) | ( g0 ) | ( m1 ) | ( (~ g)  &  (~ h)  &  (~ i)  &  h0 ) ;
 assign l10 = ( (~ r2)  &  (~ q2)  &  (~ p2)  &  o2 ) ;
 assign n10 = ( (~ o2) ) | ( n2 ) | ( (~ e1) ) | ( (~ l9) ) ;
 assign u10 = ( k2 ) | ( h ) | ( g ) | ( (~ x10) ) ;
 assign v10 = ( i0 ) | ( v2  &  g0 ) ;
 assign x10 = ( m2  &  l2 ) ;
 assign y10 = ( o1 ) | ( (~ e1) ) ;
 assign z10 = ( g  &  g0  &  v2  &  m1 ) | ( h  &  g0  &  v2  &  m1 ) | ( (~ h0)  &  g0  &  v2  &  m1 ) ;
 assign a11 = ( (~ v2) ) | ( (~ m1) ) ;
 assign c11 = ( (~ m0)  &  e1 ) | ( (~ h0)  &  v2  &  g0  &  m1 ) | ( v2  &  g0  &  g  &  m1 ) | ( v2  &  g0  &  h  &  m1 ) ;
 assign e11 = ( h0  &  (~ i)  &  (~ h)  &  (~ g) ) ;
 assign f11 = ( (~ i0)  &  m0  &  (~ o1) ) | ( (~ i0)  &  (~ e1)  &  (~ o1) ) | ( (~ i0)  &  (~ o1)  &  p1 ) | ( (~ i0)  &  (~ m0)  &  e1  &  p1 ) ;
 assign i11 = ( (~ v2) ) | ( (~ m1) ) | ( i0 ) ;
 assign j11 = ( (~ q1) ) | ( (~ e1) ) ;
 assign k11 = ( g  &  g0  &  v2  &  m1 ) | ( h  &  g0  &  v2  &  m1 ) | ( i  &  g0  &  v2  &  m1 ) | ( (~ h0)  &  g0  &  v2  &  m1 ) ;
 assign l11 = ( e1  &  (~ m0) ) | ( v2  &  m1  &  g0  &  (~ e11) ) ;
 assign n11 = ( (~ r1) ) | ( (~ e1) ) ;
 assign q11 = ( (~ s1) ) | ( (~ e1) ) ;
 assign t11 = ( (~ t1) ) | ( (~ e1) ) ;
 assign w11 = ( (~ u1) ) | ( (~ e1) ) ;
 assign z11 = ( (~ v1) ) | ( (~ e1) ) ;
 assign c12 = ( (~ w1) ) | ( (~ e1) ) ;
 assign f12 = ( (~ x1) ) | ( (~ e1) ) ;
 assign i12 = ( (~ y1) ) | ( (~ e1) ) ;
 assign l12 = ( (~ z1) ) | ( (~ e1) ) ;
 assign o12 = ( (~ a2) ) | ( (~ e1) ) ;
 assign r12 = ( (~ b2) ) | ( (~ e1) ) ;
 assign u12 = ( (~ c2) ) | ( (~ e1) ) ;
 assign x12 = ( (~ d2) ) | ( (~ e1) ) ;
 assign a13 = ( (~ e2) ) | ( (~ e1) ) ;
 assign d13 = ( (~ f2) ) | ( (~ e1) ) ;
 assign g13 = ( (~ g2) ) | ( (~ e1) ) ;
 assign j13 = ( (~ h2) ) | ( (~ e1) ) ;
 assign m13 = ( (~ i2) ) | ( (~ e1) ) ;
 assign p13 = ( (~ j2) ) | ( (~ e1) ) ;
 assign u13 = ( u0 ) | ( (~ b) ) ;
 assign v13 = ( c1 ) | ( k2  &  u2 ) | ( (~ u0)  &  b  &  k2 ) ;
 assign w13 = ( u2 ) | ( (~ u0)  &  b ) ;
 assign x13 = ( c1 ) | ( (~ k2)  &  (~ l2) ) | ( (~ k2)  &  m2 ) ;
 assign y13 = ( c1 ) | ( (~ k2)  &  l2 ) | ( (~ k2)  &  (~ m2) ) | ( (~ l2)  &  (~ m2) ) ;
 assign z13 = ( (~ m2) ) | ( (~ l2) ) | ( k2 ) ;
 assign a14 = ( c1 ) | ( e1  &  n2 ) | ( n2  &  d1 ) | ( (~ k2)  &  n2  &  l2  &  m2 ) ;
 assign b14 = ( e1 ) | ( d1 ) | ( (~ k2)  &  l2  &  m2 ) ;
 assign c14 = ( c1 ) | ( (~ n2)  &  (~ o2) ) ;
 assign d14 = ( c1 ) | ( (~ n2)  &  (~ p2) ) | ( (~ o2)  &  (~ p2) ) ;
 assign e14 = ( q2  &  p2 ) ;
 assign f14 = ( c1 ) | ( (~ n2)  &  (~ q2) ) | ( (~ o2)  &  (~ q2) ) | ( (~ p2)  &  (~ q2) ) ;
 assign g14 = ( r2  &  q2  &  p2 ) ;
 assign h14 = ( (~ q2) ) | ( (~ p2) ) | ( (~ o2) ) | ( (~ n2) ) ;
 assign j14 = ( i0 ) | ( (~ b)  &  (~ u2) ) | ( (~ u2)  &  u0 ) ;
 assign k14 = ( (~ e1) ) | ( (~ n2) ) | ( (~ l14) ) ;
 assign l14 = ( i  &  (~ p2)  &  (~ o2)  &  r2 ) | ( q2  &  (~ p2)  &  (~ o2)  &  r2 ) ;


endmodule

