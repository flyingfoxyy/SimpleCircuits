module C5315 (
	P_4115_177_, P_4092_176_, P_4091_175_, P_4090_174_, P_4089_173_, P_4088_172_, P_4087_171_, P_3724_170_, 
	P_3717_169_, P_3552_168_, P_3550_167_, P_3548_166_, P_3546_165_, P_3173_164_, P_2824_163_, P_2358_162_, P_2174_161_, P_1694_160_, 
	P_1691_159_, P_1690_158_, P_1689_157_, P_1497_156_, P_562_155_, P_559_154_, P_556_153_, P_552_152_, P_549_151_, P_545_150_, 
	P_534_149_, P_523_148_, P_514_147_, P_503_146_, P_490_145_, P_479_144_, P_468_143_, P_457_142_, P_446_141_, P_435_140_, 
	P_422_139_, P_411_138_, P_400_137_, P_389_136_, P_386_135_, P_374_134_, P_373_133_, P_372_132_, P_369_131_, P_366_130_, 
	P_361_129_, P_358_128_, P_351_127_, P_348_126_, P_341_125_, P_338_124_, P_335_123_, P_332_122_, P_331_121_, P_324_120_, 
	P_323_119_, P_316_118_, P_315_117_, P_308_116_, P_307_115_, P_302_114_, P_299_113_, P_293_112_, P_292_111_, P_289_110_, 
	P_288_109_, P_281_108_, P_280_107_, P_273_106_, P_272_105_, P_265_104_, P_264_103_, P_257_102_, P_254_101_, P_251_100_, 
	P_248_99_, P_245_98_, P_242_97_, P_241_96_, P_234_95_, P_233_94_, P_226_93_, P_225_92_, P_218_91_, P_217_90_, 
	P_210_89_, P_209_88_, P_206_87_, P_203_86_, P_200_85_, P_197_84_, P_194_83_, P_191_82_, P_188_81_, P_185_80_, 
	P_182_79_, P_179_78_, P_176_77_, P_173_76_, P_170_75_, P_167_74_, P_164_73_, P_161_72_, P_158_71_, P_155_70_, 
	P_152_69_, P_149_68_, P_146_67_, P_145_66_, P_141_65_, P_140_64_, P_137_63_, P_136_62_, P_135_61_, P_132_60_, 
	P_131_59_, P_130_58_, P_129_57_, P_128_56_, P_127_55_, P_126_54_, P_123_53_, P_122_52_, P_121_51_, P_120_50_, 
	P_119_49_, P_118_48_, P_117_47_, P_116_46_, P_115_45_, P_114_44_, P_113_43_, P_112_42_, P_109_41_, P_106_40_, 
	P_103_39_, P_100_38_, P_97_37_, P_94_36_, P_91_35_, P_88_34_, P_87_33_, P_86_32_, P_83_31_, P_82_30_, 
	P_81_29_, P_80_28_, P_79_27_, P_76_26_, P_73_25_, P_70_24_, P_67_23_, P_64_22_, P_61_21_, P_54_20_, 
	P_53_19_, P_52_18_, P_49_17_, P_46_16_, P_43_15_, P_40_14_, P_37_13_, P_34_12_, P_31_11_, P_27_10_, 
	P_26_9_, P_25_8_, P_24_7_, P_23_6_, P_20_5_, P_17_4_, P_14_3_, P_11_2_, P_4_1_, P_1_0_, 
	P_1004_1977_, P_1002_1920_, P_1000_2168_, P_998_2163_, P_993_850_, P_978_851_, P_973_202_, P_949_852_, P_939_853_, P_926_624_, 
	P_923_619_, P_921_664_, P_892_408_, P_889_734_, P_887_528_, P_882_2456_, P_877_2126_, P_875_2125_, P_873_2124_, P_871_2127_, 
	P_869_2181_, P_867_2237_, P_865_2277_, P_863_2276_, P_861_2070_, P_859_2132_, P_854_2268_, P_851_218_, P_850_217_, P_849_219_, 
	P_848_330_, P_847_465_, P_845_845_, P_843_2455_, P_838_2064_, P_836_2128_, P_834_2123_, P_832_2133_, P_830_2182_, P_828_2233_, 
	P_826_2275_, P_824_2274_, P_822_1933_, P_820_1283_, P_818_2273_, P_815_627_, P_813_2260_, P_810_356_, P_809_655_, P_807_2480_, 
	P_802_2183_, P_797_2191_, P_792_2188_, P_787_2186_, P_782_2239_, P_777_2278_, P_772_2299_, P_767_2479_, P_762_2184_, P_757_2190_, 
	P_752_2189_, P_747_2187_, P_742_2238_, P_737_2279_, P_732_2300_, P_727_2298_, P_722_2131_, P_717_1282_, P_715_1278_, P_712_2297_, 
	P_707_1277_, P_704_1281_, P_702_2228_, P_699_2227_, P_696_2226_, P_693_2179_, P_690_2484_, P_688_2317_, P_685_2316_, P_682_2296_, 
	P_679_2272_, P_676_2229_, P_673_1276_, P_670_2225_, P_667_2224_, P_664_2223_, P_661_2178_, P_658_2483_, P_656_621_, P_654_2315_, 
	P_651_2314_, P_648_2295_, P_645_2271_, P_642_2222_, P_639_1275_, P_636_1280_, P_634_665_, P_632_1692_, P_629_1926_, P_626_1752_, 
	P_623_2152_, P_621_1893_, P_618_1925_, P_615_1750_, P_612_263_, P_611_275_, P_610_1519_, P_606_407_, P_604_223_, P_603_225_, 
	P_602_222_, P_601_220_, P_600_259_, P_599_269_, P_598_1623_, P_594_224_, P_593_733_, P_591_1894_, P_588_1696_, P_585_2236_, 
	P_575_2240_, P_298_299_, P_144_354_);

input P_4115_177_, P_4092_176_, P_4091_175_, P_4090_174_, P_4089_173_, P_4088_172_, P_4087_171_, P_3724_170_, P_3717_169_, P_3552_168_, P_3550_167_, P_3548_166_, P_3546_165_, P_3173_164_, P_2824_163_, P_2358_162_, P_2174_161_, P_1694_160_, P_1691_159_, P_1690_158_, P_1689_157_, P_1497_156_, P_562_155_, P_559_154_, P_556_153_, P_552_152_, P_549_151_, P_545_150_, P_534_149_, P_523_148_, P_514_147_, P_503_146_, P_490_145_, P_479_144_, P_468_143_, P_457_142_, P_446_141_, P_435_140_, P_422_139_, P_411_138_, P_400_137_, P_389_136_, P_386_135_, P_374_134_, P_373_133_, P_372_132_, P_369_131_, P_366_130_, P_361_129_, P_358_128_, P_351_127_, P_348_126_, P_341_125_, P_338_124_, P_335_123_, P_332_122_, P_331_121_, P_324_120_, P_323_119_, P_316_118_, P_315_117_, P_308_116_, P_307_115_, P_302_114_, P_299_113_, P_293_112_, P_292_111_, P_289_110_, P_288_109_, P_281_108_, P_280_107_, P_273_106_, P_272_105_, P_265_104_, P_264_103_, P_257_102_, P_254_101_, P_251_100_, P_248_99_, P_245_98_, P_242_97_, P_241_96_, P_234_95_, P_233_94_, P_226_93_, P_225_92_, P_218_91_, P_217_90_, P_210_89_, P_209_88_, P_206_87_, P_203_86_, P_200_85_, P_197_84_, P_194_83_, P_191_82_, P_188_81_, P_185_80_, P_182_79_, P_179_78_, P_176_77_, P_173_76_, P_170_75_, P_167_74_, P_164_73_, P_161_72_, P_158_71_, P_155_70_, P_152_69_, P_149_68_, P_146_67_, P_145_66_, P_141_65_, P_140_64_, P_137_63_, P_136_62_, P_135_61_, P_132_60_, P_131_59_, P_130_58_, P_129_57_, P_128_56_, P_127_55_, P_126_54_, P_123_53_, P_122_52_, P_121_51_, P_120_50_, P_119_49_, P_118_48_, P_117_47_, P_116_46_, P_115_45_, P_114_44_, P_113_43_, P_112_42_, P_109_41_, P_106_40_, P_103_39_, P_100_38_, P_97_37_, P_94_36_, P_91_35_, P_88_34_, P_87_33_, P_86_32_, P_83_31_, P_82_30_, P_81_29_, P_80_28_, P_79_27_, P_76_26_, P_73_25_, P_70_24_, P_67_23_, P_64_22_, P_61_21_, P_54_20_, P_53_19_, P_52_18_, P_49_17_, P_46_16_, P_43_15_, P_40_14_, P_37_13_, P_34_12_, P_31_11_, P_27_10_, P_26_9_, P_25_8_, P_24_7_, P_23_6_, P_20_5_, P_17_4_, P_14_3_, P_11_2_, P_4_1_, P_1_0_;

output P_1004_1977_, P_1002_1920_, P_1000_2168_, P_998_2163_, P_993_850_, P_978_851_, P_973_202_, P_949_852_, P_939_853_, P_926_624_, P_923_619_, P_921_664_, P_892_408_, P_889_734_, P_887_528_, P_882_2456_, P_877_2126_, P_875_2125_, P_873_2124_, P_871_2127_, P_869_2181_, P_867_2237_, P_865_2277_, P_863_2276_, P_861_2070_, P_859_2132_, P_854_2268_, P_851_218_, P_850_217_, P_849_219_, P_848_330_, P_847_465_, P_845_845_, P_843_2455_, P_838_2064_, P_836_2128_, P_834_2123_, P_832_2133_, P_830_2182_, P_828_2233_, P_826_2275_, P_824_2274_, P_822_1933_, P_820_1283_, P_818_2273_, P_815_627_, P_813_2260_, P_810_356_, P_809_655_, P_807_2480_, P_802_2183_, P_797_2191_, P_792_2188_, P_787_2186_, P_782_2239_, P_777_2278_, P_772_2299_, P_767_2479_, P_762_2184_, P_757_2190_, P_752_2189_, P_747_2187_, P_742_2238_, P_737_2279_, P_732_2300_, P_727_2298_, P_722_2131_, P_717_1282_, P_715_1278_, P_712_2297_, P_707_1277_, P_704_1281_, P_702_2228_, P_699_2227_, P_696_2226_, P_693_2179_, P_690_2484_, P_688_2317_, P_685_2316_, P_682_2296_, P_679_2272_, P_676_2229_, P_673_1276_, P_670_2225_, P_667_2224_, P_664_2223_, P_661_2178_, P_658_2483_, P_656_621_, P_654_2315_, P_651_2314_, P_648_2295_, P_645_2271_, P_642_2222_, P_639_1275_, P_636_1280_, P_634_665_, P_632_1692_, P_629_1926_, P_626_1752_, P_623_2152_, P_621_1893_, P_618_1925_, P_615_1750_, P_612_263_, P_611_275_, P_610_1519_, P_606_407_, P_604_223_, P_603_225_, P_602_222_, P_601_220_, P_600_259_, P_599_269_, P_598_1623_, P_594_224_, P_593_733_, P_591_1894_, P_588_1696_, P_585_2236_, P_575_2240_, P_298_299_, P_144_354_;

wire wire102, wire103, n193, n548, n287, n36, n40, n41, n39, n38, n44, n45, n43, n42, n48, n49, n47, n46, n52, n53, n51, n50, n56, n57, n55, n54, n60, n61, n59, n58, n64, n65, n63, n62, n68, n69, n67, n66, n72, n73, n71, n70, n76, n77, n75, n74, n80, n81, n79, n78, n84, n85, n83, n82, n88, n89, n87, n86, n92, n93, n91, n90, n96, n97, n95, n94, n100, n101, n99, n98, n104, n105, n103, n102, n108, n109, n107, n106, n112, n113, n111, n110, n116, n117, n115, n114, n120, n121, n119, n118, n124, n125, n123, n122, n128, n129, n127, n126, n132, n133, n131, n130, n140, n141, n139, n138, n147, n153, n156, n154, n158, n157, n160, n165, n166, n163, n164, n162, n167, n172, n171, n177, n178, n175, n176, n174, n180, n181, n179, n183, n184, n182, n186, n185, n188, n189, n187, n191, n190, n194, n197, n195, n199, n200, n198, n203, n204, n202, n207, n208, n209, n210, n206, n212, n213, n214, n215, n211, n217, n219, n221, n223, n225, n227, n229, n231, n233, n235, n237, n238, n239, n241, n243, n244, n245, n247, n249, n251, n253, n254, n258, n262, n263, n260, n259, n267, n268, n265, n266, n264, n271, n270, n269, n274, n275, n273, n272, n278, n279, n277, n276, n283, n280, n286, n284, n288, n289, n290, n291, n292, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n311, n312, n313, n314, n315, n316, n317, n319, n320, n321, n324, n325, n329, n333, n334, n332, n336, n337, n335, n339, n340, n338, n342, n343, n341, n345, n346, n344, n347, n348, n350, n351, n349, n353, n354, n352, n356, n357, n355, n358, n359, n360, n364, n365, n363, n367, n368, n366, n370, n371, n369, n373, n374, n372, n376, n377, n375, n379, n380, n378, n382, n383, n381, n385, n386, n384, n388, n392, n390, n391, n389, n394, n396, n397, n395, n399, n400, n398, n401, n402, n404, n405, n408, n409, n407, n411, n412, n410, n414, n415, n413, n416, n417, n419, n420, n418, n422, n423, n421, n424, n425, n427, n428, n426, n430, n431, n429, n433, n434, n432, n436, n437, n435, n439, n440, n438, n442, n443, n441, n445, n446, n444, n448, n449, n447, n451, n452, n450, n454, n455, n453, n457, n458, n456, n460, n459, n461, n462, n464, n463, n465, n466, n467, n468, n470, n469, n472, n473, n471, n474, n476, n477, n478, n480, n482, n483, n485, n484, n486, n487, n489, n488, n492, n491, n493, n494, n497, n501, n500, n504, n503, n505, n507, n511, n510, n512, n514, n515, n519, n518, n521, n520, n523, n522, n527, n526, n530, n529, n532, n535, n538, n537, n539, n541, n543, n542, n545, n544, n547, n549, n550, n552, n554, n556, n558, n560, n562, n566, n568, n569, n570, n572, n574, n575, n578, n580, n581, n582, n583, n586, n589, n597, n599, n608, n609, n611, n613, n623, n624, n626, n633, n634, n636, n638, n639, n640, n642, n644, n645, n646, n647, n648, n666, n668, n667, n669, n671, n673, n672, n675, n674, n678, n679, n677, n681, n682, n680, n684, n685, n683, n686, n688, n687, n690, n689, n692, n693, n691, n696, n697, n699, n701, n703, n704, n705, n706, n707, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n720, n721, n722, n723, n724, n726, n727, n725, n728, n730, n731, n732, n734, n735, n736, n737, n738, n739, n740, n741, n743, n744, n745, n748, n747, n750, n753, n754, n755, n758, n757, n760, n761, n762, n766, n768, n770, n771, n773, n778, n779, n781, n780, n783, n784, n786, n787, n789, n788, n790, n791, n793, n792, n794, n796, n799, n800, n801, n802, n805, n803, n806, n809, n810, n819, n820, n822, n824, n825, n826, n827, n829, n831, n833, n835, n837, n839, n840, n844, n846, n847, n848, n849, n850, n851, n852, n859, n860, n861, n862, n867, n868, n869, n871, n877;

assign P_1004_1977_ = ( (~ n482)  &  n483 ) | ( n482  &  (~ n483) ) ;
 assign P_1002_1920_ = ( (~ n476)  &  n477 ) | ( n476  &  (~ n477) ) ;
 assign P_1000_2168_ = ( (~ n493)  &  n494 ) | ( n493  &  (~ n494) ) ;
 assign P_998_2163_ = ( (~ n486)  &  n487 ) | ( n486  &  (~ n487) ) ;
 assign P_882_2456_ = ( (~ n302) ) ;
 assign P_877_2126_ = ( (~ P_126_54_)  &  n227 ) | ( n195  &  n227 ) ;
 assign P_875_2125_ = ( (~ P_127_55_)  &  n225 ) | ( n195  &  n225 ) ;
 assign P_873_2124_ = ( (~ P_128_56_)  &  n223 ) | ( n195  &  n223 ) ;
 assign P_871_2127_ = ( (~ P_122_52_)  &  n229 ) | ( n195  &  n229 ) ;
 assign P_869_2181_ = ( (~ P_113_43_)  &  n235 ) | ( n195  &  n235 ) ;
 assign P_867_2237_ = ( (~ P_53_19_)  &  n243 ) | ( n195  &  n243 ) ;
 assign P_865_2277_ = ( (~ P_114_44_)  &  n253 ) | ( n195  &  n253 ) ;
 assign P_863_2276_ = ( (~ P_115_45_)  &  n251 ) | ( n195  &  n251 ) ;
 assign P_861_2070_ = ( (~ P_117_47_)  &  n219 ) | ( n195  &  n219 ) ;
 assign P_859_2132_ = ( (~ n306) ) ;
 assign P_854_2268_ = ( (~ n254) ) ;
 assign P_851_218_ = ( (~ P_559_154_) ) ;
 assign P_850_217_ = ( (~ P_562_155_) ) ;
 assign P_849_219_ = ( (~ P_552_152_) ) ;
 assign P_848_330_ = ( (~ P_245_98_) ) ;
 assign P_847_465_ = ( (~ n316) ) ;
 assign P_845_845_ = ( P_2824_163_ ) | ( (~ P_27_10_) ) ;
 assign P_843_2455_ = ( (~ n303) ) ;
 assign P_838_2064_ = ( (~ P_129_57_)  &  n217 ) | ( n195  &  n217 ) ;
 assign P_836_2128_ = ( (~ P_119_49_)  &  n231 ) | ( n195  &  n231 ) ;
 assign P_834_2123_ = ( (~ P_130_58_)  &  n221 ) | ( n195  &  n221 ) ;
 assign P_832_2133_ = ( (~ P_52_18_)  &  n233 ) | ( n195  &  n233 ) ;
 assign P_830_2182_ = ( (~ P_112_42_)  &  n237 ) | ( n195  &  n237 ) ;
 assign P_828_2233_ = ( (~ P_116_46_)  &  n241 ) | ( n195  &  n241 ) ;
 assign P_826_2275_ = ( (~ P_121_51_)  &  n249 ) | ( n195  &  n249 ) ;
 assign P_824_2274_ = ( (~ P_123_53_)  &  n247 ) | ( n195  &  n247 ) ;
 assign P_822_1933_ = ( (~ P_131_59_)  &  n197 ) | ( n197  &  n195 ) ;
 assign P_820_1283_ = ( (~ n321) ) ;
 assign P_818_2273_ = ( (~ P_4115_177_)  &  n258 ) | ( (~ P_135_61_)  &  n258 ) ;
 assign P_815_627_ = ( (~ P_3173_164_)  &  P_136_62_ ) ;
 assign P_813_2260_ = ( P_623_2152_  &  n666 ) | ( (~ P_623_2152_)  &  (~ n666) ) ;
 assign P_810_356_ = ( P_141_65_  &  P_145_66_ ) ;
 assign P_809_655_ = ( (~ n36) ) ;
 assign P_807_2480_ = ( (~ n300) ) ;
 assign P_802_2183_ = ( (~ n305) ) ;
 assign P_797_2191_ = ( (~ n355) ) ;
 assign P_792_2188_ = ( (~ n352) ) ;
 assign P_787_2186_ = ( (~ n349) ) ;
 assign P_782_2239_ = ( (~ n384) ) ;
 assign P_777_2278_ = ( (~ n381) ) ;
 assign P_772_2299_ = ( (~ n378) ) ;
 assign P_767_2479_ = ( (~ n301) ) ;
 assign P_762_2184_ = ( (~ n304) ) ;
 assign P_757_2190_ = ( (~ n344) ) ;
 assign P_752_2189_ = ( (~ n341) ) ;
 assign P_747_2187_ = ( (~ n338) ) ;
 assign P_742_2238_ = ( (~ n375) ) ;
 assign P_737_2279_ = ( (~ n372) ) ;
 assign P_732_2300_ = ( (~ n369) ) ;
 assign P_727_2298_ = ( (~ n366) ) ;
 assign P_722_2131_ = ( (~ n307) ) ;
 assign P_717_1282_ = ( (~ n308) ) ;
 assign P_715_1278_ = ( P_141_65_  &  (~ n36) ) | ( P_141_65_  &  (~ n714) ) ;
 assign P_712_2297_ = ( (~ n363) ) ;
 assign P_707_1277_ = ( P_141_65_  &  (~ n36) ) | ( P_141_65_  &  (~ n713) ) ;
 assign P_704_1281_ = ( (~ n308) ) ;
 assign P_702_2228_ = ( (~ n429) ) ;
 assign P_699_2227_ = ( (~ n426) ) ;
 assign P_696_2226_ = ( (~ n245) ) ;
 assign P_693_2179_ = ( (~ n239) ) ;
 assign P_690_2484_ = ( (~ n298) ) ;
 assign P_688_2317_ = ( (~ n456) ) ;
 assign P_685_2316_ = ( (~ n453) ) ;
 assign P_682_2296_ = ( (~ n444) ) ;
 assign P_679_2272_ = ( (~ n438) ) ;
 assign P_676_2229_ = ( (~ n432) ) ;
 assign P_673_1276_ = ( P_141_65_  &  (~ n36) ) | ( P_141_65_  &  (~ n712) ) ;
 assign P_670_2225_ = ( (~ n421) ) ;
 assign P_667_2224_ = ( (~ n418) ) ;
 assign P_664_2223_ = ( (~ n244) ) ;
 assign P_661_2178_ = ( (~ n238) ) ;
 assign P_658_2483_ = ( (~ n299) ) ;
 assign P_656_621_ = ( (~ n317) ) ;
 assign P_654_2315_ = ( (~ n450) ) ;
 assign P_651_2314_ = ( (~ n447) ) ;
 assign P_648_2295_ = ( (~ n441) ) ;
 assign P_645_2271_ = ( (~ n435) ) ;
 assign P_642_2222_ = ( (~ n413) ) ;
 assign P_639_1275_ = ( P_141_65_  &  (~ n36) ) | ( P_141_65_  &  (~ n711) ) ;
 assign P_636_1280_ = ( (~ n309) ) ;
 assign P_634_665_ = ( P_373_133_  &  P_1_0_ ) ;
 assign P_632_1692_ = ( (~ n852) ) ;
 assign P_623_2152_ = ( (~ n193)  &  n770 ) | ( n193  &  n771 ) | ( n770  &  n771 ) ;
 assign P_621_1893_ = ( (~ n311) ) ;
 assign wire102 = ( n312 ) | ( n313 ) | ( n314 ) | ( n315 ) ;
 assign wire103 = ( (~ n189)  &  (~ n315)  &  n634 ) ;
 assign P_612_263_ = ( (~ P_358_128_) ) ;
 assign P_611_275_ = ( (~ P_338_124_) ) ;
 assign P_610_1519_ = ( (~ n74)  &  (~ n82)  &  (~ n90)  &  (~ n98)  &  (~ n102)  &  n147 ) ;
 assign P_606_407_ = ( (~ P_549_151_) ) ;
 assign P_604_223_ = ( (~ P_545_150_) ) ;
 assign P_603_225_ = ( (~ P_545_150_) ) ;
 assign P_602_222_ = ( (~ P_549_151_) ) ;
 assign P_601_220_ = ( P_552_152_  &  P_562_155_ ) ;
 assign P_600_259_ = ( (~ P_366_130_) ) ;
 assign P_599_269_ = ( (~ P_348_126_) ) ;
 assign P_598_1623_ = ( (~ n42)  &  (~ n46)  &  (~ n54)  &  (~ n62)  &  (~ n66)  &  n153 ) ;
 assign P_594_224_ = ( (~ P_545_150_) ) ;
 assign P_593_733_ = ( (~ P_299_113_) ) ;
 assign P_591_1894_ = ( (~ n311) ) ;
 assign P_588_1696_ = ( (~ n852) ) ;
 assign P_585_2236_ = ( P_623_2152_  &  n287  &  n288  &  n289  &  n290  &  n291 ) ;
 assign P_575_2240_ = ( n292  &  n294  &  n295  &  n296  &  n297  &  (~ n329) ) ;
 assign n193 = ( n163  &  n162 ) | ( n162  &  (~ n597) ) ;
 assign n548 = ( (~ P_490_145_)  &  n527 ) | ( P_490_145_  &  (~ n527) ) ;
 assign n287 = ( (~ n193)  &  n548 ) | ( n193  &  (~ n548) ) ;
 assign n36 = ( P_31_11_  &  P_27_10_ ) ;
 assign n40 = ( (~ P_534_149_) ) | ( P_351_127_ ) | ( (~ P_251_100_) ) ;
 assign n41 = ( (~ P_248_99_) ) | ( n556 ) ;
 assign n39 = ( (~ P_351_127_)  &  P_254_101_ ) | ( P_351_127_  &  P_242_97_ ) | ( P_254_101_  &  P_242_97_ ) ;
 assign n38 = ( n40  &  n41  &  P_534_149_ ) | ( n40  &  n41  &  n39 ) ;
 assign n44 = ( P_3550_167_ ) | ( (~ P_534_149_) ) | ( P_351_127_ ) ;
 assign n45 = ( P_3552_168_ ) | ( n556 ) ;
 assign n43 = ( (~ P_3548_166_)  &  (~ P_3546_165_) ) | ( (~ P_3546_165_)  &  P_351_127_ ) | ( (~ P_3548_166_)  &  (~ P_351_127_) ) ;
 assign n42 = ( n44  &  n45  &  P_534_149_ ) | ( n44  &  n45  &  n43 ) ;
 assign n48 = ( P_3550_167_ ) | ( (~ P_523_148_) ) | ( P_341_125_ ) ;
 assign n49 = ( P_3552_168_ ) | ( n572 ) ;
 assign n47 = ( (~ P_3548_166_)  &  (~ P_3546_165_) ) | ( (~ P_3546_165_)  &  P_341_125_ ) | ( (~ P_3548_166_)  &  (~ P_341_125_) ) ;
 assign n46 = ( n48  &  n49  &  P_523_148_ ) | ( n48  &  n49  &  n47 ) ;
 assign n52 = ( (~ P_523_148_) ) | ( P_341_125_ ) | ( (~ P_251_100_) ) ;
 assign n53 = ( (~ P_248_99_) ) | ( n572 ) ;
 assign n51 = ( (~ P_341_125_)  &  P_254_101_ ) | ( P_341_125_  &  P_242_97_ ) | ( P_254_101_  &  P_242_97_ ) ;
 assign n50 = ( n52  &  n53  &  P_523_148_ ) | ( n52  &  n53  &  n51 ) ;
 assign n56 = ( P_3550_167_ ) | ( (~ P_503_146_) ) | ( P_324_120_ ) ;
 assign n57 = ( P_3552_168_ ) | ( n568 ) ;
 assign n55 = ( (~ P_3548_166_)  &  (~ P_3546_165_) ) | ( (~ P_3546_165_)  &  P_324_120_ ) | ( (~ P_3548_166_)  &  (~ P_324_120_) ) ;
 assign n54 = ( n56  &  n57  &  P_503_146_ ) | ( n56  &  n57  &  n55 ) ;
 assign n60 = ( (~ P_503_146_) ) | ( P_324_120_ ) | ( (~ P_251_100_) ) ;
 assign n61 = ( (~ P_248_99_) ) | ( n568 ) ;
 assign n59 = ( (~ P_324_120_)  &  P_254_101_ ) | ( P_324_120_  &  P_242_97_ ) | ( P_254_101_  &  P_242_97_ ) ;
 assign n58 = ( n60  &  n61  &  P_503_146_ ) | ( n60  &  n61  &  n59 ) ;
 assign n64 = ( (~ P_490_145_) ) | ( P_316_118_ ) | ( (~ P_251_100_) ) ;
 assign n65 = ( (~ P_490_145_) ) | ( (~ P_316_118_) ) | ( (~ P_248_99_) ) ;
 assign n63 = ( (~ P_316_118_)  &  P_254_101_ ) | ( P_316_118_  &  P_242_97_ ) | ( P_254_101_  &  P_242_97_ ) ;
 assign n62 = ( n64  &  n65  &  P_490_145_ ) | ( n64  &  n65  &  n63 ) ;
 assign n68 = ( (~ P_479_144_) ) | ( (~ P_308_116_) ) | ( (~ P_248_99_) ) ;
 assign n69 = ( (~ P_479_144_) ) | ( P_308_116_ ) | ( (~ P_251_100_) ) ;
 assign n67 = ( (~ P_308_116_)  &  P_254_101_ ) | ( P_308_116_  &  P_242_97_ ) | ( P_254_101_  &  P_242_97_ ) ;
 assign n66 = ( n68  &  n69  &  P_479_144_ ) | ( n68  &  n69  &  n67 ) ;
 assign n72 = ( (~ P_468_143_) ) | ( (~ P_251_100_) ) | ( P_218_91_ ) ;
 assign n73 = ( (~ P_248_99_) ) | ( n611 ) ;
 assign n71 = ( P_254_101_  &  P_242_97_ ) | ( P_242_97_  &  P_218_91_ ) | ( P_254_101_  &  (~ P_218_91_) ) ;
 assign n70 = ( n72  &  n73  &  P_468_143_ ) | ( n72  &  n73  &  n71 ) ;
 assign n76 = ( P_3550_167_ ) | ( (~ P_468_143_) ) | ( P_218_91_ ) ;
 assign n77 = ( P_3552_168_ ) | ( n611 ) ;
 assign n75 = ( (~ P_3548_166_)  &  (~ P_3546_165_) ) | ( (~ P_3546_165_)  &  P_218_91_ ) | ( (~ P_3548_166_)  &  (~ P_218_91_) ) ;
 assign n74 = ( n76  &  n77  &  P_468_143_ ) | ( n76  &  n77  &  n75 ) ;
 assign n80 = ( (~ P_457_142_) ) | ( (~ P_251_100_) ) | ( P_210_89_ ) ;
 assign n81 = ( (~ P_248_99_) ) | ( n608 ) ;
 assign n79 = ( P_254_101_  &  P_242_97_ ) | ( P_242_97_  &  P_210_89_ ) | ( P_254_101_  &  (~ P_210_89_) ) ;
 assign n78 = ( n80  &  n81  &  P_457_142_ ) | ( n80  &  n81  &  n79 ) ;
 assign n84 = ( P_3550_167_ ) | ( (~ P_457_142_) ) | ( P_210_89_ ) ;
 assign n85 = ( P_3552_168_ ) | ( n608 ) ;
 assign n83 = ( (~ P_3548_166_)  &  (~ P_3546_165_) ) | ( (~ P_3546_165_)  &  P_210_89_ ) | ( (~ P_3548_166_)  &  (~ P_210_89_) ) ;
 assign n82 = ( n84  &  n85  &  P_457_142_ ) | ( n84  &  n85  &  n83 ) ;
 assign n88 = ( (~ P_435_140_) ) | ( (~ P_251_100_) ) | ( P_234_95_ ) ;
 assign n89 = ( (~ P_248_99_) ) | ( n580 ) ;
 assign n87 = ( P_254_101_  &  P_242_97_ ) | ( P_242_97_  &  P_234_95_ ) | ( P_254_101_  &  (~ P_234_95_) ) ;
 assign n86 = ( n88  &  n89  &  P_435_140_ ) | ( n88  &  n89  &  n87 ) ;
 assign n92 = ( P_3550_167_ ) | ( (~ P_435_140_) ) | ( P_234_95_ ) ;
 assign n93 = ( P_3552_168_ ) | ( n580 ) ;
 assign n91 = ( (~ P_3548_166_)  &  (~ P_3546_165_) ) | ( (~ P_3546_165_)  &  P_234_95_ ) | ( (~ P_3548_166_)  &  (~ P_234_95_) ) ;
 assign n90 = ( n92  &  n93  &  P_435_140_ ) | ( n92  &  n93  &  n91 ) ;
 assign n96 = ( (~ P_422_139_) ) | ( (~ P_251_100_) ) | ( P_226_93_ ) ;
 assign n97 = ( (~ P_248_99_) ) | ( n613 ) ;
 assign n95 = ( P_254_101_  &  P_242_97_ ) | ( P_242_97_  &  P_226_93_ ) | ( P_254_101_  &  (~ P_226_93_) ) ;
 assign n94 = ( n96  &  n97  &  P_422_139_ ) | ( n96  &  n97  &  n95 ) ;
 assign n100 = ( P_3550_167_ ) | ( (~ P_422_139_) ) | ( P_226_93_ ) ;
 assign n101 = ( P_3552_168_ ) | ( n613 ) ;
 assign n99 = ( (~ P_3548_166_)  &  (~ P_3546_165_) ) | ( (~ P_3546_165_)  &  P_226_93_ ) | ( (~ P_3548_166_)  &  (~ P_226_93_) ) ;
 assign n98 = ( n100  &  n101  &  P_422_139_ ) | ( n100  &  n101  &  n99 ) ;
 assign n104 = ( P_3550_167_ ) | ( (~ P_411_138_) ) | ( P_273_106_ ) ;
 assign n105 = ( P_3552_168_ ) | ( n589 ) ;
 assign n103 = ( (~ P_3548_166_)  &  (~ P_3546_165_) ) | ( (~ P_3546_165_)  &  P_273_106_ ) | ( (~ P_3548_166_)  &  (~ P_273_106_) ) ;
 assign n102 = ( n104  &  n105  &  P_411_138_ ) | ( n104  &  n105  &  n103 ) ;
 assign n108 = ( (~ P_411_138_) ) | ( P_273_106_ ) | ( (~ P_251_100_) ) ;
 assign n109 = ( (~ P_248_99_) ) | ( n589 ) ;
 assign n107 = ( (~ P_273_106_)  &  P_254_101_ ) | ( P_273_106_  &  P_242_97_ ) | ( P_254_101_  &  P_242_97_ ) ;
 assign n106 = ( n108  &  n109  &  P_411_138_ ) | ( n108  &  n109  &  n107 ) ;
 assign n112 = ( (~ P_400_137_) ) | ( P_265_104_ ) | ( (~ P_251_100_) ) ;
 assign n113 = ( (~ P_248_99_) ) | ( n586 ) ;
 assign n111 = ( (~ P_265_104_)  &  P_254_101_ ) | ( P_265_104_  &  P_242_97_ ) | ( P_254_101_  &  P_242_97_ ) ;
 assign n110 = ( n112  &  n113  &  P_400_137_ ) | ( n112  &  n113  &  n111 ) ;
 assign n116 = ( P_3550_167_ ) | ( (~ P_400_137_) ) | ( P_265_104_ ) ;
 assign n117 = ( P_3552_168_ ) | ( n586 ) ;
 assign n115 = ( (~ P_3548_166_)  &  (~ P_3546_165_) ) | ( (~ P_3546_165_)  &  P_265_104_ ) | ( (~ P_3548_166_)  &  (~ P_265_104_) ) ;
 assign n114 = ( n116  &  n117  &  P_400_137_ ) | ( n116  &  n117  &  n115 ) ;
 assign n120 = ( P_3550_167_ ) | ( (~ P_389_136_) ) | ( P_257_102_ ) ;
 assign n121 = ( P_3552_168_ ) | ( n583 ) ;
 assign n119 = ( (~ P_3548_166_)  &  (~ P_3546_165_) ) | ( (~ P_3546_165_)  &  P_257_102_ ) | ( (~ P_3548_166_)  &  (~ P_257_102_) ) ;
 assign n118 = ( n120  &  n121  &  P_389_136_ ) | ( n120  &  n121  &  n119 ) ;
 assign n124 = ( (~ P_389_136_) ) | ( P_257_102_ ) | ( (~ P_251_100_) ) ;
 assign n125 = ( (~ P_248_99_) ) | ( n583 ) ;
 assign n123 = ( (~ P_257_102_)  &  P_254_101_ ) | ( P_257_102_  &  P_242_97_ ) | ( P_254_101_  &  P_242_97_ ) ;
 assign n122 = ( n124  &  n125  &  P_389_136_ ) | ( n124  &  n125  &  n123 ) ;
 assign n128 = ( (~ P_374_134_) ) | ( P_281_108_ ) | ( (~ P_251_100_) ) ;
 assign n129 = ( (~ P_248_99_) ) | ( n560 ) ;
 assign n127 = ( (~ P_281_108_)  &  P_254_101_ ) | ( P_281_108_  &  P_242_97_ ) | ( P_254_101_  &  P_242_97_ ) ;
 assign n126 = ( n128  &  n129  &  P_374_134_ ) | ( n128  &  n129  &  n127 ) ;
 assign n132 = ( P_3550_167_ ) | ( (~ P_374_134_) ) | ( P_281_108_ ) ;
 assign n133 = ( P_3552_168_ ) | ( n560 ) ;
 assign n131 = ( (~ P_3548_166_)  &  (~ P_3546_165_) ) | ( (~ P_3546_165_)  &  P_281_108_ ) | ( (~ P_3548_166_)  &  (~ P_281_108_) ) ;
 assign n130 = ( n132  &  n133  &  P_374_134_ ) | ( n132  &  n133  &  n131 ) ;
 assign n140 = ( (~ P_446_141_) ) | ( (~ P_251_100_) ) | ( P_206_87_ ) ;
 assign n141 = ( (~ P_446_141_) ) | ( (~ P_248_99_) ) | ( (~ P_206_87_) ) ;
 assign n139 = ( P_254_101_  &  P_242_97_ ) | ( P_242_97_  &  P_206_87_ ) | ( P_254_101_  &  (~ P_206_87_) ) ;
 assign n138 = ( n140  &  n141  &  P_446_141_ ) | ( n140  &  n141  &  n139 ) ;
 assign n147 = ( (~ n114)  &  (~ n118)  &  (~ n130)  &  (~ n138) ) ;
 assign n153 = ( n701  &  (~ n703)  &  n717  &  n722 ) ;
 assign n156 = ( (~ n545)  &  n569 ) ;
 assign n154 = ( n156 ) | ( (~ n570) ) ;
 assign n158 = ( n535  &  n547  &  n164  &  n539 ) ;
 assign n157 = ( n158  &  (~ n624) ) ;
 assign n160 = ( n158  &  (~ n597) ) ;
 assign n165 = ( n163 ) | ( n535  &  n539 ) ;
 assign n166 = ( (~ P_503_146_)  &  n163 ) | ( (~ P_503_146_)  &  n547 ) | ( n163  &  (~ n699) ) | ( n547  &  (~ n699) ) ;
 assign n163 = ( P_503_146_  &  n699 ) | ( (~ P_503_146_)  &  (~ n699) ) ;
 assign n164 = ( (~ P_514_147_) ) | ( n541 ) ;
 assign n162 = ( n165  &  n166  &  n163 ) | ( n165  &  n166  &  n164 ) ;
 assign n167 = ( (~ P_457_142_)  &  (~ n198) ) | ( (~ n198)  &  (~ n697) ) ;
 assign n172 = ( P_457_142_  &  n697 ) | ( (~ P_457_142_)  &  (~ n697) ) ;
 assign n171 = ( n167  &  n172 ) | ( n167  &  (~ n518) ) ;
 assign n177 = ( n175 ) | ( n503  &  n507 ) ;
 assign n178 = ( (~ P_435_140_)  &  n175 ) | ( n175  &  (~ n489) ) | ( (~ P_435_140_)  &  n515 ) | ( (~ n489)  &  n515 ) ;
 assign n175 = ( P_435_140_  &  n489 ) | ( (~ P_435_140_)  &  (~ n489) ) ;
 assign n176 = ( (~ P_389_136_) ) | ( (~ n758) ) ;
 assign n174 = ( n177  &  n178  &  n175 ) | ( n177  &  n178  &  n176 ) ;
 assign n180 = ( n505  &  n500  &  n514 ) ;
 assign n181 = ( n501 ) | ( n582 ) ;
 assign n179 = ( n180  &  n181 ) ;
 assign n183 = ( n507  &  n515  &  n176  &  n503 ) ;
 assign n184 = ( n504 ) | ( n181 ) ;
 assign n182 = ( n183  &  n184 ) ;
 assign n186 = ( n504 ) | ( n626 ) ;
 assign n185 = ( n183  &  n186 ) ;
 assign n188 = ( (~ n312)  &  (~ n550)  &  (~ n849) ) ;
 assign n189 = ( n312 ) | ( (~ n325) ) ;
 assign n187 = ( n188  &  n189 ) ;
 assign n191 = ( (~ n312)  &  n360 ) ;
 assign n190 = ( n191  &  (~ n325) ) ;
 assign n194 = ( n174  &  n175 ) | ( n174  &  n184 ) ;
 assign n197 = ( n701  &  n715 ) | ( n552  &  n715 ) | ( n701  &  n554 ) | ( n552  &  n554 ) ;
 assign n195 = ( (~ P_4092_176_) ) | ( P_4091_175_ ) ;
 assign n199 = ( n762  &  P_468_143_ ) ;
 assign n200 = ( n266  &  n522 ) ;
 assign n198 = ( (~ n172)  &  n199 ) | ( (~ n172)  &  n200 ) ;
 assign n203 = ( (~ P_54_20_)  &  (~ n543) ) ;
 assign n204 = ( (~ n530)  &  P_534_149_ ) | ( n530  &  (~ P_534_149_) ) ;
 assign n202 = ( P_54_20_  &  n203 ) | ( P_54_20_  &  n204 ) | ( n203  &  (~ n558) ) | ( n204  &  (~ n558) ) ;
 assign n207 = ( n484 ) | ( n835 ) | ( (~ n848) ) ;
 assign n208 = ( (~ n484) ) | ( (~ n835) ) | ( (~ n848) ) ;
 assign n209 = ( n484 ) | ( (~ n835) ) | ( n848 ) ;
 assign n210 = ( (~ n484) ) | ( n835 ) | ( n848 ) ;
 assign n206 = ( n207  &  n208  &  n209  &  n210 ) ;
 assign n212 = ( n488 ) | ( (~ n491) ) | ( n837 ) ;
 assign n213 = ( (~ n488) ) | ( (~ n491) ) | ( (~ n837) ) ;
 assign n214 = ( n488 ) | ( n491 ) | ( (~ n837) ) ;
 assign n215 = ( (~ n488) ) | ( n491 ) | ( n837 ) ;
 assign n211 = ( n212  &  n213  &  n214  &  n215 ) ;
 assign n217 = ( (~ n42)  &  n202 ) | ( n202  &  n552 ) | ( (~ n42)  &  n554 ) | ( n552  &  n554 ) ;
 assign n219 = ( (~ n130)  &  (~ n329) ) | ( (~ n329)  &  n552 ) | ( (~ n130)  &  n554 ) | ( n552  &  n554 ) ;
 assign n221 = ( n717  &  n459 ) | ( n552  &  n459 ) | ( n717  &  n554 ) | ( n552  &  n554 ) ;
 assign n223 = ( (~ n118)  &  n554 ) | ( n552  &  n554 ) | ( (~ n118)  &  (~ n844) ) | ( n552  &  (~ n844) ) ;
 assign n225 = ( (~ n114)  &  n554 ) | ( n552  &  n554 ) | ( (~ n114)  &  n720 ) | ( n552  &  n720 ) ;
 assign n227 = ( (~ n102)  &  n554 ) | ( n552  &  n554 ) | ( (~ n102)  &  n721 ) | ( n552  &  n721 ) ;
 assign n229 = ( (~ n90)  &  n554 ) | ( n552  &  n554 ) | ( (~ n90)  &  n718 ) | ( n552  &  n718 ) ;
 assign n231 = ( (~ n46)  &  n290 ) | ( n290  &  n552 ) | ( (~ n46)  &  n554 ) | ( n552  &  n554 ) ;
 assign n233 = ( (~ n54)  &  n554 ) | ( n552  &  n554 ) | ( (~ n54)  &  n716 ) | ( n552  &  n716 ) ;
 assign n235 = ( (~ n98)  &  n292 ) | ( n292  &  n552 ) | ( (~ n98)  &  n554 ) | ( n552  &  n554 ) ;
 assign n237 = ( n287  &  (~ n62) ) | ( n287  &  n552 ) | ( (~ n62)  &  n554 ) | ( n552  &  n554 ) ;
 assign n238 = ( n408  &  n409  &  P_861_2070_ ) | ( n408  &  n409  &  n407 ) ;
 assign n239 = ( n411  &  n412  &  P_861_2070_ ) | ( n411  &  n412  &  n410 ) ;
 assign n241 = ( (~ n66)  &  n288 ) | ( n288  &  n552 ) | ( (~ n66)  &  n554 ) | ( n552  &  n554 ) ;
 assign n243 = ( (~ n74)  &  n294 ) | ( n294  &  n552 ) | ( (~ n74)  &  n554 ) | ( n552  &  n554 ) ;
 assign n244 = ( n416  &  n417  &  P_877_2126_ ) | ( n416  &  n417  &  n407 ) ;
 assign n245 = ( n424  &  n425  &  P_877_2126_ ) | ( n424  &  n425  &  n410 ) ;
 assign n247 = ( P_623_2152_  &  n552 ) | ( n552  &  n554 ) | ( P_623_2152_  &  (~ n703) ) | ( n554  &  (~ n703) ) ;
 assign n249 = ( n722  &  n289 ) | ( n552  &  n289 ) | ( n722  &  n554 ) | ( n552  &  n554 ) ;
 assign n251 = ( (~ n138)  &  n296 ) | ( n296  &  n552 ) | ( (~ n138)  &  n554 ) | ( n552  &  n554 ) ;
 assign n253 = ( (~ n82)  &  n295 ) | ( n295  &  n552 ) | ( (~ n82)  &  n554 ) | ( n552  &  n554 ) ;
 assign n254 = ( (~ P_559_154_) ) | ( (~ P_245_98_) ) | ( P_1004_1977_ ) | ( P_1002_1920_ ) | ( P_1000_2168_ ) | ( P_998_2163_ ) | ( (~ P_601_220_) ) | ( (~ n316) ) ;
 assign n258 = ( (~ P_3717_169_)  &  n839 ) | ( P_3717_169_  &  n840 ) | ( n839  &  n840 ) ;
 assign n262 = ( n548 ) | ( (~ n463) ) | ( n727 ) ;
 assign n263 = ( (~ n325) ) | ( n463 ) ;
 assign n260 = ( (~ n548)  &  n463 ) | ( n548  &  (~ n463) ) ;
 assign n259 = ( n262  &  n263  &  n260 ) | ( n262  &  n263  &  (~ n727) ) ;
 assign n267 = ( (~ n266) ) | ( (~ n469) ) | ( n519 ) ;
 assign n268 = ( n469 ) | ( (~ n518) ) ;
 assign n265 = ( (~ n519)  &  n469 ) | ( n519  &  (~ n469) ) ;
 assign n266 = ( (~ n762)  &  P_468_143_ ) | ( n762  &  (~ P_468_143_) ) ;
 assign n264 = ( n267  &  n268  &  n265 ) | ( n267  &  n268  &  n266 ) ;
 assign n271 = ( (~ n542)  &  (~ n558) ) | ( (~ n542)  &  n790 ) | ( (~ n558)  &  (~ n790) ) ;
 assign n270 = ( n543  &  n790 ) | ( (~ n543)  &  (~ n790) ) ;
 assign n269 = ( n271  &  n204 ) | ( n271  &  n270 ) ;
 assign n274 = ( P_2174_161_ ) | ( (~ n162) ) | ( n788 ) ;
 assign n275 = ( n789  &  n788 ) | ( n789  &  n787 ) ;
 assign n273 = ( (~ n461)  &  n462 ) | ( n461  &  (~ n462) ) ;
 assign n272 = ( n274  &  n275  &  n162 ) | ( n274  &  n275  &  n273 ) ;
 assign n278 = ( P_1497_156_ ) | ( (~ n174) ) | ( n803 ) ;
 assign n279 = ( (~ n802)  &  n805 ) | ( n805  &  n803 ) ;
 assign n277 = ( (~ n467)  &  n468 ) | ( n467  &  (~ n468) ) ;
 assign n276 = ( n278  &  n279  &  n174 ) | ( n278  &  n279  &  n277 ) ;
 assign n283 = ( n552  &  n554 ) | ( n552  &  n689 ) | ( n554  &  (~ n691) ) | ( n689  &  (~ n691) ) ;
 assign n280 = ( (~ P_4092_176_)  &  n283 ) | ( (~ P_97_37_)  &  n283 ) ;
 assign n286 = ( (~ n471)  &  n554 ) | ( n552  &  n554 ) | ( (~ n471)  &  n687 ) | ( n552  &  n687 ) ;
 assign n284 = ( (~ P_4092_176_)  &  n286 ) | ( (~ P_94_36_)  &  n286 ) ;
 assign n288 = ( (~ n193)  &  n667 ) | ( n193  &  (~ n705) ) | ( n667  &  (~ n705) ) ;
 assign n289 = ( n193  &  (~ n704) ) | ( (~ n193)  &  n773 ) | ( (~ n704)  &  n773 ) ;
 assign n290 = ( (~ n545)  &  n766 ) | ( (~ n569)  &  (~ n574)  &  n766 ) ;
 assign n291 = ( n715  &  n202  &  n459  &  n716 ) ;
 assign n292 = ( (~ n194)  &  n519 ) | ( n194  &  (~ n519) ) ;
 assign n294 = ( (~ n194)  &  n674 ) | ( n194  &  (~ n707) ) | ( n674  &  (~ n707) ) ;
 assign n295 = ( (~ n194)  &  n672 ) | ( n194  &  (~ n706) ) | ( n672  &  (~ n706) ) ;
 assign n296 = ( n194  &  n669 ) | ( (~ n194)  &  n671 ) | ( n669  &  n671 ) ;
 assign n297 = ( n718  &  n720  &  n721  &  (~ n844) ) ;
 assign n298 = ( P_137_63_  &  n404 ) | ( P_137_63_  &  n405 ) | ( P_137_63_  &  (~ n710) ) ;
 assign n299 = ( P_137_63_  &  n401 ) | ( P_137_63_  &  n402 ) | ( P_137_63_  &  (~ n709) ) ;
 assign n300 = ( n399  &  n400  &  n284 ) | ( n399  &  n400  &  n398 ) ;
 assign n301 = ( n396  &  n397  &  n284 ) | ( n396  &  n397  &  n395 ) ;
 assign n302 = ( (~ P_4092_176_)  &  n394 ) | ( (~ P_118_48_)  &  n394 ) ;
 assign n303 = ( (~ P_4092_176_)  &  n388 ) | ( (~ P_120_50_)  &  n388 ) ;
 assign n304 = ( n347  &  n348  &  P_877_2126_ ) | ( n347  &  n348  &  n332 ) ;
 assign n305 = ( n358  &  n359  &  P_877_2126_ ) | ( n358  &  n359  &  n335 ) ;
 assign n306 = ( n336  &  n337  &  P_861_2070_ ) | ( n336  &  n337  &  n335 ) ;
 assign n307 = ( n333  &  n334  &  P_861_2070_ ) | ( n333  &  n334  &  n332 ) ;
 assign n308 = ( (~ P_2358_162_)  &  n36  &  n320 ) | ( P_34_12_  &  n36  &  n320 ) ;
 assign n309 = ( (~ P_2358_162_)  &  n36  &  n319 ) | ( P_87_33_  &  n36  &  n319 ) ;
 assign n311 = ( (~ P_446_141_)  &  n324 ) | ( n324  &  (~ n696) ) ;
 assign n312 = ( P_332_122_  &  P_307_115_ ) | ( (~ P_332_122_)  &  P_302_114_ ) | ( P_307_115_  &  P_302_114_ ) ;
 assign n313 = ( n549 ) | ( n550 ) ;
 assign n314 = ( (~ n162)  &  n325 ) ;
 assign n315 = ( P_332_122_  &  P_299_113_ ) | ( (~ P_332_122_)  &  P_293_112_ ) | ( P_299_113_  &  P_293_112_ ) ;
 assign n316 = ( P_386_135_  &  P_556_153_ ) ;
 assign n317 = ( P_140_64_  &  n36 ) ;
 assign n319 = ( P_86_32_ ) | ( P_2358_162_ ) ;
 assign n320 = ( P_88_34_ ) | ( P_2358_162_ ) ;
 assign n321 = ( P_83_31_  &  n36 ) ;
 assign n324 = ( n174  &  n167 ) | ( n520  &  n167 ) | ( n174  &  n521 ) | ( n520  &  n521 ) ;
 assign n325 = ( n548  &  (~ n727) ) ;
 assign n329 = ( P_4_1_  &  (~ n581) ) | ( (~ n391)  &  (~ n581) ) ;
 assign n333 = ( (~ P_61_21_) ) | ( n566 ) ;
 assign n334 = ( (~ P_11_2_)  &  P_822_1933_ ) | ( (~ P_11_2_)  &  n395 ) | ( P_822_1933_  &  n562 ) | ( n395  &  n562 ) ;
 assign n332 = ( (~ P_4088_172_) ) | ( P_4087_171_ ) ;
 assign n336 = ( (~ P_61_21_) ) | ( n578 ) ;
 assign n337 = ( (~ P_11_2_)  &  P_822_1933_ ) | ( (~ P_11_2_)  &  n398 ) | ( P_822_1933_  &  n575 ) | ( n398  &  n575 ) ;
 assign n335 = ( P_4090_174_ ) | ( (~ P_4089_173_) ) ;
 assign n339 = ( (~ P_37_13_)  &  P_871_2127_ ) | ( (~ P_37_13_)  &  n332 ) | ( P_871_2127_  &  n566 ) | ( n332  &  n566 ) ;
 assign n340 = ( (~ P_43_15_)  &  P_832_2133_ ) | ( (~ P_43_15_)  &  n395 ) | ( P_832_2133_  &  n562 ) | ( n395  &  n562 ) ;
 assign n338 = ( n339  &  n340 ) ;
 assign n342 = ( (~ P_20_5_)  &  P_873_2124_ ) | ( (~ P_20_5_)  &  n332 ) | ( P_873_2124_  &  n566 ) | ( n332  &  n566 ) ;
 assign n343 = ( (~ P_76_26_)  &  P_834_2123_ ) | ( (~ P_76_26_)  &  n395 ) | ( P_834_2123_  &  n562 ) | ( n395  &  n562 ) ;
 assign n341 = ( n342  &  n343 ) ;
 assign n345 = ( (~ P_17_4_)  &  P_875_2125_ ) | ( (~ P_17_4_)  &  n332 ) | ( P_875_2125_  &  n566 ) | ( n332  &  n566 ) ;
 assign n346 = ( (~ P_73_25_)  &  P_836_2128_ ) | ( (~ P_73_25_)  &  n395 ) | ( P_836_2128_  &  n562 ) | ( n395  &  n562 ) ;
 assign n344 = ( n345  &  n346 ) ;
 assign n347 = ( (~ P_70_24_) ) | ( n566 ) ;
 assign n348 = ( (~ P_67_23_)  &  P_838_2064_ ) | ( (~ P_67_23_)  &  n395 ) | ( P_838_2064_  &  n562 ) | ( n395  &  n562 ) ;
 assign n350 = ( (~ P_37_13_)  &  P_871_2127_ ) | ( (~ P_37_13_)  &  n335 ) | ( P_871_2127_  &  n578 ) | ( n335  &  n578 ) ;
 assign n351 = ( (~ P_43_15_)  &  P_832_2133_ ) | ( (~ P_43_15_)  &  n398 ) | ( P_832_2133_  &  n575 ) | ( n398  &  n575 ) ;
 assign n349 = ( n350  &  n351 ) ;
 assign n353 = ( (~ P_20_5_)  &  P_873_2124_ ) | ( (~ P_20_5_)  &  n335 ) | ( P_873_2124_  &  n578 ) | ( n335  &  n578 ) ;
 assign n354 = ( (~ P_76_26_)  &  P_834_2123_ ) | ( (~ P_76_26_)  &  n398 ) | ( P_834_2123_  &  n575 ) | ( n398  &  n575 ) ;
 assign n352 = ( n353  &  n354 ) ;
 assign n356 = ( (~ P_17_4_)  &  P_875_2125_ ) | ( (~ P_17_4_)  &  n335 ) | ( P_875_2125_  &  n578 ) | ( n335  &  n578 ) ;
 assign n357 = ( (~ P_73_25_)  &  P_836_2128_ ) | ( (~ P_73_25_)  &  n398 ) | ( P_836_2128_  &  n575 ) | ( n398  &  n575 ) ;
 assign n355 = ( n356  &  n357 ) ;
 assign n358 = ( (~ P_70_24_) ) | ( n578 ) ;
 assign n359 = ( (~ P_67_23_)  &  P_838_2064_ ) | ( (~ P_67_23_)  &  n398 ) | ( P_838_2064_  &  n575 ) | ( n398  &  n575 ) ;
 assign n360 = ( n312  &  (~ n849) ) | ( (~ n550)  &  (~ n849) ) ;
 assign n364 = ( (~ P_106_40_)  &  P_863_2276_ ) | ( (~ P_106_40_)  &  n335 ) | ( P_863_2276_  &  n578 ) | ( n335  &  n578 ) ;
 assign n365 = ( (~ P_109_41_)  &  P_824_2274_ ) | ( (~ P_109_41_)  &  n398 ) | ( P_824_2274_  &  n575 ) | ( n398  &  n575 ) ;
 assign n363 = ( n364  &  n365 ) ;
 assign n367 = ( (~ P_106_40_)  &  P_863_2276_ ) | ( (~ P_106_40_)  &  n332 ) | ( P_863_2276_  &  n566 ) | ( n332  &  n566 ) ;
 assign n368 = ( (~ P_109_41_)  &  P_824_2274_ ) | ( (~ P_109_41_)  &  n395 ) | ( P_824_2274_  &  n562 ) | ( n395  &  n562 ) ;
 assign n366 = ( n367  &  n368 ) ;
 assign n370 = ( (~ P_49_17_)  &  P_865_2277_ ) | ( (~ P_49_17_)  &  n332 ) | ( P_865_2277_  &  n566 ) | ( n332  &  n566 ) ;
 assign n371 = ( (~ P_46_16_)  &  P_826_2275_ ) | ( (~ P_46_16_)  &  n395 ) | ( P_826_2275_  &  n562 ) | ( n395  &  n562 ) ;
 assign n369 = ( n370  &  n371 ) ;
 assign n373 = ( (~ P_103_39_)  &  P_867_2237_ ) | ( (~ P_103_39_)  &  n332 ) | ( P_867_2237_  &  n566 ) | ( n332  &  n566 ) ;
 assign n374 = ( (~ P_100_38_)  &  P_828_2233_ ) | ( (~ P_100_38_)  &  n395 ) | ( P_828_2233_  &  n562 ) | ( n395  &  n562 ) ;
 assign n372 = ( n373  &  n374 ) ;
 assign n376 = ( (~ P_40_14_)  &  P_869_2181_ ) | ( (~ P_40_14_)  &  n332 ) | ( P_869_2181_  &  n566 ) | ( n332  &  n566 ) ;
 assign n377 = ( (~ P_91_35_)  &  P_830_2182_ ) | ( (~ P_91_35_)  &  n395 ) | ( P_830_2182_  &  n562 ) | ( n395  &  n562 ) ;
 assign n375 = ( n376  &  n377 ) ;
 assign n379 = ( (~ P_49_17_)  &  P_865_2277_ ) | ( (~ P_49_17_)  &  n335 ) | ( P_865_2277_  &  n578 ) | ( n335  &  n578 ) ;
 assign n380 = ( (~ P_46_16_)  &  P_826_2275_ ) | ( (~ P_46_16_)  &  n398 ) | ( P_826_2275_  &  n575 ) | ( n398  &  n575 ) ;
 assign n378 = ( n379  &  n380 ) ;
 assign n382 = ( (~ P_103_39_)  &  P_867_2237_ ) | ( (~ P_103_39_)  &  n335 ) | ( P_867_2237_  &  n578 ) | ( n335  &  n578 ) ;
 assign n383 = ( (~ P_100_38_)  &  P_828_2233_ ) | ( (~ P_100_38_)  &  n398 ) | ( P_828_2233_  &  n575 ) | ( n398  &  n575 ) ;
 assign n381 = ( n382  &  n383 ) ;
 assign n385 = ( (~ P_40_14_)  &  P_869_2181_ ) | ( (~ P_40_14_)  &  n335 ) | ( P_869_2181_  &  n578 ) | ( n335  &  n578 ) ;
 assign n386 = ( (~ P_91_35_)  &  P_830_2182_ ) | ( (~ P_91_35_)  &  n398 ) | ( P_830_2182_  &  n575 ) | ( n398  &  n575 ) ;
 assign n384 = ( n385  &  n386 ) ;
 assign n388 = ( (~ P_4091_175_)  &  n734 ) | ( (~ P_4092_176_)  &  (~ n687)  &  n734 ) ;
 assign n392 = ( n497  &  n512 ) ;
 assign n390 = ( P_411_138_  &  n761 ) | ( (~ P_411_138_)  &  (~ n761) ) ;
 assign n391 = ( P_374_134_  &  n511 ) | ( (~ P_374_134_)  &  (~ n511) ) ;
 assign n389 = ( n392  &  n390 ) | ( n392  &  n391 ) ;
 assign n394 = ( (~ P_4091_175_)  &  n750 ) | ( (~ P_4092_176_)  &  (~ n689)  &  n750 ) ;
 assign n396 = ( (~ P_14_3_) ) | ( n562 ) ;
 assign n397 = ( (~ P_64_22_)  &  n280 ) | ( (~ P_64_22_)  &  n332 ) | ( n280  &  n566 ) | ( n332  &  n566 ) ;
 assign n395 = ( P_4088_172_ ) | ( P_4087_171_ ) ;
 assign n399 = ( (~ P_14_3_) ) | ( n575 ) ;
 assign n400 = ( (~ P_64_22_)  &  n280 ) | ( (~ P_64_22_)  &  n335 ) | ( n280  &  n578 ) | ( n335  &  n578 ) ;
 assign n398 = ( P_4089_173_ ) | ( P_4090_174_ ) ;
 assign n401 = ( (~ P_1690_158_)  &  (~ P_1689_157_)  &  (~ n284) ) ;
 assign n402 = ( P_1690_158_  &  (~ P_1689_157_)  &  P_176_77_ ) ;
 assign n404 = ( (~ P_1694_160_)  &  (~ P_1691_159_)  &  (~ n284) ) ;
 assign n405 = ( P_1694_160_  &  (~ P_1691_159_)  &  P_176_77_ ) ;
 assign n408 = ( P_822_1933_ ) | ( n638 ) ;
 assign n409 = ( (~ P_185_80_)  &  (~ P_182_79_) ) | ( (~ P_185_80_)  &  n640 ) | ( (~ P_182_79_)  &  n642 ) | ( n640  &  n642 ) ;
 assign n407 = ( P_1690_158_ ) | ( n639 ) ;
 assign n411 = ( P_822_1933_ ) | ( n645 ) ;
 assign n412 = ( (~ P_185_80_)  &  (~ P_182_79_) ) | ( (~ P_185_80_)  &  n647 ) | ( (~ P_182_79_)  &  n648 ) | ( n647  &  n648 ) ;
 assign n410 = ( P_1694_160_ ) | ( n646 ) ;
 assign n414 = ( (~ P_200_85_)  &  (~ P_170_75_) ) | ( (~ P_170_75_)  &  n640 ) | ( (~ P_200_85_)  &  n642 ) | ( n640  &  n642 ) ;
 assign n415 = ( P_832_2133_  &  P_871_2127_ ) | ( n638  &  P_871_2127_ ) | ( P_832_2133_  &  n407 ) | ( n638  &  n407 ) ;
 assign n413 = ( n414  &  n415 ) ;
 assign n416 = ( P_838_2064_ ) | ( n638 ) ;
 assign n417 = ( (~ P_188_81_)  &  (~ P_158_71_) ) | ( (~ P_158_71_)  &  n640 ) | ( (~ P_188_81_)  &  n642 ) | ( n640  &  n642 ) ;
 assign n419 = ( (~ P_155_70_)  &  (~ P_152_69_) ) | ( (~ P_152_69_)  &  n640 ) | ( (~ P_155_70_)  &  n642 ) | ( n640  &  n642 ) ;
 assign n420 = ( P_836_2128_  &  P_875_2125_ ) | ( n638  &  P_875_2125_ ) | ( P_836_2128_  &  n407 ) | ( n638  &  n407 ) ;
 assign n418 = ( n419  &  n420 ) ;
 assign n422 = ( (~ P_149_68_)  &  (~ P_146_67_) ) | ( (~ P_146_67_)  &  n640 ) | ( (~ P_149_68_)  &  n642 ) | ( n640  &  n642 ) ;
 assign n423 = ( P_834_2123_  &  P_873_2124_ ) | ( n638  &  P_873_2124_ ) | ( P_834_2123_  &  n407 ) | ( n638  &  n407 ) ;
 assign n421 = ( n422  &  n423 ) ;
 assign n424 = ( P_838_2064_ ) | ( n645 ) ;
 assign n425 = ( (~ P_188_81_)  &  (~ P_158_71_) ) | ( (~ P_158_71_)  &  n647 ) | ( (~ P_188_81_)  &  n648 ) | ( n647  &  n648 ) ;
 assign n427 = ( (~ P_155_70_)  &  (~ P_152_69_) ) | ( (~ P_152_69_)  &  n647 ) | ( (~ P_155_70_)  &  n648 ) | ( n647  &  n648 ) ;
 assign n428 = ( P_836_2128_  &  P_875_2125_ ) | ( n645  &  P_875_2125_ ) | ( P_836_2128_  &  n410 ) | ( n645  &  n410 ) ;
 assign n426 = ( n427  &  n428 ) ;
 assign n430 = ( (~ P_149_68_)  &  (~ P_146_67_) ) | ( (~ P_146_67_)  &  n647 ) | ( (~ P_149_68_)  &  n648 ) | ( n647  &  n648 ) ;
 assign n431 = ( P_834_2123_  &  P_873_2124_ ) | ( n645  &  P_873_2124_ ) | ( P_834_2123_  &  n410 ) | ( n645  &  n410 ) ;
 assign n429 = ( n430  &  n431 ) ;
 assign n433 = ( (~ P_200_85_)  &  (~ P_170_75_) ) | ( (~ P_170_75_)  &  n647 ) | ( (~ P_200_85_)  &  n648 ) | ( n647  &  n648 ) ;
 assign n434 = ( P_832_2133_  &  P_871_2127_ ) | ( n645  &  P_871_2127_ ) | ( P_832_2133_  &  n410 ) | ( n645  &  n410 ) ;
 assign n432 = ( n433  &  n434 ) ;
 assign n436 = ( (~ P_203_86_)  &  (~ P_173_76_) ) | ( (~ P_173_76_)  &  n640 ) | ( (~ P_203_86_)  &  n642 ) | ( n640  &  n642 ) ;
 assign n437 = ( P_830_2182_  &  P_869_2181_ ) | ( n638  &  P_869_2181_ ) | ( P_830_2182_  &  n407 ) | ( n638  &  n407 ) ;
 assign n435 = ( n436  &  n437 ) ;
 assign n439 = ( (~ P_203_86_)  &  (~ P_173_76_) ) | ( (~ P_173_76_)  &  n647 ) | ( (~ P_203_86_)  &  n648 ) | ( n647  &  n648 ) ;
 assign n440 = ( P_830_2182_  &  P_869_2181_ ) | ( n645  &  P_869_2181_ ) | ( P_830_2182_  &  n410 ) | ( n645  &  n410 ) ;
 assign n438 = ( n439  &  n440 ) ;
 assign n442 = ( (~ P_197_84_)  &  (~ P_167_74_) ) | ( (~ P_167_74_)  &  n640 ) | ( (~ P_197_84_)  &  n642 ) | ( n640  &  n642 ) ;
 assign n443 = ( P_828_2233_  &  P_867_2237_ ) | ( n638  &  P_867_2237_ ) | ( P_828_2233_  &  n407 ) | ( n638  &  n407 ) ;
 assign n441 = ( n442  &  n443 ) ;
 assign n445 = ( (~ P_197_84_)  &  (~ P_167_74_) ) | ( (~ P_167_74_)  &  n647 ) | ( (~ P_197_84_)  &  n648 ) | ( n647  &  n648 ) ;
 assign n446 = ( P_828_2233_  &  P_867_2237_ ) | ( n645  &  P_867_2237_ ) | ( P_828_2233_  &  n410 ) | ( n645  &  n410 ) ;
 assign n444 = ( n445  &  n446 ) ;
 assign n448 = ( (~ P_194_83_)  &  (~ P_164_73_) ) | ( (~ P_164_73_)  &  n640 ) | ( (~ P_194_83_)  &  n642 ) | ( n640  &  n642 ) ;
 assign n449 = ( P_826_2275_  &  P_865_2277_ ) | ( n638  &  P_865_2277_ ) | ( P_826_2275_  &  n407 ) | ( n638  &  n407 ) ;
 assign n447 = ( n448  &  n449 ) ;
 assign n451 = ( (~ P_191_82_)  &  (~ P_161_72_) ) | ( (~ P_161_72_)  &  n640 ) | ( (~ P_191_82_)  &  n642 ) | ( n640  &  n642 ) ;
 assign n452 = ( P_824_2274_  &  P_863_2276_ ) | ( n638  &  P_863_2276_ ) | ( P_824_2274_  &  n407 ) | ( n638  &  n407 ) ;
 assign n450 = ( n451  &  n452 ) ;
 assign n454 = ( (~ P_194_83_)  &  (~ P_164_73_) ) | ( (~ P_164_73_)  &  n647 ) | ( (~ P_194_83_)  &  n648 ) | ( n647  &  n648 ) ;
 assign n455 = ( P_826_2275_  &  P_865_2277_ ) | ( n645  &  P_865_2277_ ) | ( P_826_2275_  &  n410 ) | ( n645  &  n410 ) ;
 assign n453 = ( n454  &  n455 ) ;
 assign n457 = ( (~ P_191_82_)  &  (~ P_161_72_) ) | ( (~ P_161_72_)  &  n647 ) | ( (~ P_191_82_)  &  n648 ) | ( n647  &  n648 ) ;
 assign n458 = ( P_824_2274_  &  P_863_2276_ ) | ( n645  &  P_863_2276_ ) | ( P_824_2274_  &  n410 ) | ( n645  &  n410 ) ;
 assign n456 = ( n457  &  n458 ) ;
 assign n460 = ( (~ P_514_147_)  &  n541 ) | ( P_514_147_  &  (~ n541) ) ;
 assign n459 = ( (~ n154)  &  n460 ) | ( n154  &  (~ n460) ) ;
 assign n461 = ( (~ n724)  &  n725 ) | ( n724  &  (~ n725) ) ;
 assign n462 = ( (~ n312)  &  n867 ) | ( n312  &  (~ n867) ) ;
 assign n464 = ( (~ n526)  &  n313 ) | ( n526  &  (~ n313) ) ;
 assign n463 = ( (~ n191)  &  n464 ) | ( n191  &  (~ n464) ) ;
 assign n465 = ( (~ n86)  &  n122 ) | ( n86  &  (~ n122) ) ;
 assign n466 = ( (~ n106)  &  n110 ) | ( n106  &  (~ n110) ) ;
 assign n467 = ( (~ n736)  &  n737 ) | ( n736  &  (~ n737) ) ;
 assign n468 = ( (~ n519)  &  n869 ) | ( n519  &  (~ n869) ) ;
 assign n470 = ( (~ n522)  &  n609 ) | ( n522  &  (~ n609) ) ;
 assign n469 = ( (~ n167)  &  n470 ) | ( n167  &  (~ n470) ) ;
 assign n472 = ( n784 ) | ( n786 ) | ( n780 ) | ( n783 ) ;
 assign n473 = ( (~ n723)  &  n859 ) | ( n723  &  (~ n859) ) ;
 assign n471 = ( (~ n472)  &  n473 ) | ( n472  &  (~ n473) ) ;
 assign n474 = ( P_369_131_  &  P_361_129_ ) | ( (~ P_369_131_)  &  (~ P_361_129_) ) ;
 assign n476 = ( P_302_114_  &  n753 ) | ( (~ P_302_114_)  &  (~ n753) ) ;
 assign n477 = ( P_293_112_  &  n850 ) | ( (~ P_293_112_)  &  (~ n850) ) ;
 assign n478 = ( P_257_102_  &  P_234_95_ ) | ( (~ P_257_102_)  &  (~ P_234_95_) ) ;
 assign n480 = ( P_289_110_  &  P_281_108_ ) | ( (~ P_289_110_)  &  (~ P_281_108_) ) ;
 assign n482 = ( P_226_93_  &  n754 ) | ( (~ P_226_93_)  &  (~ n754) ) ;
 assign n483 = ( P_206_87_  &  n851 ) | ( (~ P_206_87_)  &  (~ n851) ) ;
 assign n485 = ( (~ P_372_132_)  &  (~ P_369_131_) ) | ( (~ P_372_132_)  &  P_332_122_ ) | ( (~ P_369_131_)  &  (~ P_332_122_) ) ;
 assign n484 = ( n485  &  n543 ) | ( (~ n485)  &  (~ n543) ) ;
 assign n486 = ( n527  &  n755 ) | ( (~ n527)  &  (~ n755) ) ;
 assign n487 = ( (~ n312)  &  n315 ) | ( n312  &  (~ n315) ) ;
 assign n489 = ( P_335_123_  &  P_241_96_ ) | ( (~ P_335_123_)  &  P_234_95_ ) | ( P_241_96_  &  P_234_95_ ) ;
 assign n488 = ( n489  &  n523 ) | ( (~ n489)  &  (~ n523) ) ;
 assign n492 = ( P_335_123_  &  (~ P_292_111_) ) | ( (~ P_335_123_)  &  (~ P_289_110_) ) | ( (~ P_292_111_)  &  (~ P_289_110_) ) ;
 assign n491 = ( n492  &  n696 ) | ( (~ n492)  &  (~ n696) ) ;
 assign n493 = ( n757  &  n760 ) | ( (~ n757)  &  (~ n760) ) ;
 assign n494 = ( (~ n511)  &  n761 ) | ( n511  &  (~ n761) ) ;
 assign n497 = ( (~ P_411_138_) ) | ( (~ n761) ) ;
 assign n501 = ( P_400_137_  &  n760 ) | ( (~ P_400_137_)  &  (~ n760) ) ;
 assign n500 = ( n501 ) | ( n497 ) ;
 assign n504 = ( P_389_136_  &  n758 ) | ( (~ P_389_136_)  &  (~ n758) ) ;
 assign n503 = ( n504 ) | ( n500 ) ;
 assign n505 = ( (~ P_400_137_) ) | ( (~ n760) ) ;
 assign n507 = ( n504 ) | ( n505 ) ;
 assign n511 = ( P_335_123_  &  P_288_109_ ) | ( (~ P_335_123_)  &  P_281_108_ ) | ( P_288_109_  &  P_281_108_ ) ;
 assign n510 = ( n511  &  P_374_134_ ) ;
 assign n512 = ( n390 ) | ( (~ n510) ) ;
 assign n514 = ( n501 ) | ( n512 ) ;
 assign n515 = ( n504 ) | ( n514 ) ;
 assign n519 = ( (~ n523)  &  P_422_139_ ) | ( n523  &  (~ P_422_139_) ) ;
 assign n518 = ( n266  &  n519 ) ;
 assign n521 = ( P_446_141_  &  n696 ) | ( (~ P_446_141_)  &  (~ n696) ) ;
 assign n520 = ( n172 ) | ( (~ n518) ) | ( n521 ) ;
 assign n523 = ( P_335_123_  &  P_233_94_ ) | ( (~ P_335_123_)  &  P_226_93_ ) | ( P_233_94_  &  P_226_93_ ) ;
 assign n522 = ( n523  &  P_422_139_ ) ;
 assign n527 = ( P_332_122_  &  P_323_119_ ) | ( (~ P_332_122_)  &  P_316_118_ ) | ( P_323_119_  &  P_316_118_ ) ;
 assign n526 = ( n527  &  P_490_145_ ) ;
 assign n530 = ( P_358_128_  &  P_351_127_ ) | ( P_358_128_  &  P_332_122_ ) | ( P_351_127_  &  (~ P_332_122_) ) ;
 assign n529 = ( n530  &  P_534_149_ ) ;
 assign n532 = ( n529  &  (~ n545) ) ;
 assign n535 = ( n460 ) | ( (~ n532) ) ;
 assign n538 = ( P_348_126_  &  P_341_125_ ) | ( P_348_126_  &  P_332_122_ ) | ( P_341_125_  &  (~ P_332_122_) ) ;
 assign n537 = ( n538  &  P_523_148_ ) ;
 assign n539 = ( n460 ) | ( (~ n537) ) ;
 assign n541 = ( (~ P_338_124_)  &  P_332_122_ ) ;
 assign n543 = ( P_366_130_  &  P_361_129_ ) | ( P_366_130_  &  P_332_122_ ) | ( P_361_129_  &  (~ P_332_122_) ) ;
 assign n542 = ( n543  &  n204 ) ;
 assign n545 = ( P_523_148_  &  n538 ) | ( (~ P_523_148_)  &  (~ n538) ) ;
 assign n544 = ( (~ n542) ) | ( n545 ) ;
 assign n547 = ( n460 ) | ( n544 ) ;
 assign n549 = ( n599  &  P_479_144_ ) ;
 assign n550 = ( n526  &  (~ n727) ) ;
 assign n552 = ( P_4091_175_ ) | ( P_4092_176_ ) ;
 assign n554 = ( P_4092_176_ ) | ( (~ P_4091_175_) ) ;
 assign n556 = ( (~ P_534_149_) ) | ( (~ P_351_127_) ) ;
 assign n558 = ( n204  &  (~ n543) ) ;
 assign n560 = ( (~ P_374_134_) ) | ( (~ P_281_108_) ) ;
 assign n562 = ( P_4088_172_ ) | ( (~ P_4087_171_) ) ;
 assign n566 = ( (~ P_4088_172_) ) | ( (~ P_4087_171_) ) ;
 assign n568 = ( (~ P_503_146_) ) | ( (~ P_324_120_) ) ;
 assign n569 = ( P_54_20_  &  n558 ) ;
 assign n570 = ( (~ n532)  &  (~ n537)  &  n544 ) ;
 assign n572 = ( (~ P_523_148_) ) | ( (~ P_341_125_) ) ;
 assign n574 = ( n529 ) | ( n542 ) ;
 assign n575 = ( (~ P_4090_174_) ) | ( P_4089_173_ ) ;
 assign n578 = ( (~ P_4090_174_) ) | ( (~ P_4089_173_) ) ;
 assign n580 = ( (~ P_435_140_) ) | ( (~ P_234_95_) ) ;
 assign n581 = ( P_4_1_  &  (~ n391) ) ;
 assign n582 = ( n390 ) | ( (~ n581) ) ;
 assign n583 = ( (~ P_389_136_) ) | ( (~ P_257_102_) ) ;
 assign n586 = ( (~ P_400_137_) ) | ( (~ P_265_104_) ) ;
 assign n589 = ( (~ P_411_138_) ) | ( (~ P_273_106_) ) ;
 assign n597 = ( n156  &  (~ n460) ) ;
 assign n599 = ( P_332_122_  &  P_315_117_ ) | ( (~ P_332_122_)  &  P_308_116_ ) | ( P_315_117_  &  P_308_116_ ) ;
 assign n608 = ( (~ P_457_142_) ) | ( (~ P_210_89_) ) ;
 assign n609 = ( n200 ) | ( n199 ) ;
 assign n611 = ( (~ P_468_143_) ) | ( (~ P_218_91_) ) ;
 assign n613 = ( (~ P_422_139_) ) | ( (~ P_226_93_) ) ;
 assign n623 = ( (~ n545)  &  n558 ) ;
 assign n624 = ( (~ n460)  &  n623 ) ;
 assign n626 = ( n501 ) | ( n390 ) | ( n391 ) ;
 assign n633 = ( n175 ) | ( n186 ) ;
 assign n634 = ( (~ n163)  &  n624 ) ;
 assign n636 = ( P_1689_157_ ) | ( (~ P_137_63_) ) ;
 assign n638 = ( P_1690_158_ ) | ( n636 ) ;
 assign n639 = ( (~ P_1689_157_) ) | ( (~ P_137_63_) ) ;
 assign n640 = ( (~ P_1690_158_) ) | ( n636 ) ;
 assign n642 = ( (~ P_1690_158_) ) | ( n639 ) ;
 assign n644 = ( P_1691_159_ ) | ( (~ P_137_63_) ) ;
 assign n645 = ( P_1694_160_ ) | ( n644 ) ;
 assign n646 = ( (~ P_1691_159_) ) | ( (~ P_137_63_) ) ;
 assign n647 = ( (~ P_1694_160_) ) | ( n644 ) ;
 assign n648 = ( (~ P_1694_160_) ) | ( n646 ) ;
 assign n666 = ( P_132_60_  &  n315 ) | ( (~ P_132_60_)  &  (~ n315) ) ;
 assign n668 = ( (~ P_490_145_)  &  (~ n527) ) ;
 assign n667 = ( n668  &  n727 ) | ( (~ n668)  &  (~ n727) ) ;
 assign n669 = ( n167  &  n521 ) | ( (~ n167)  &  (~ n521) ) ;
 assign n671 = ( n171  &  n521 ) | ( (~ n171)  &  (~ n521) ) ;
 assign n673 = ( n518 ) | ( n609 ) ;
 assign n672 = ( (~ n673)  &  n172 ) | ( n673  &  (~ n172) ) ;
 assign n675 = ( (~ P_422_139_)  &  (~ n523) ) ;
 assign n674 = ( (~ n675)  &  n266 ) | ( n675  &  (~ n266) ) ;
 assign n678 = ( n163  &  n269 ) | ( (~ n163)  &  (~ n269) ) ;
 assign n679 = ( n460  &  n545 ) | ( (~ n460)  &  (~ n545) ) ;
 assign n677 = ( (~ n678)  &  n679 ) | ( n678  &  (~ n679) ) ;
 assign n681 = ( (~ n743)  &  n744 ) | ( n743  &  (~ n744) ) ;
 assign n682 = ( (~ n745)  &  n747 ) | ( n745  &  (~ n747) ) ;
 assign n680 = ( (~ n681)  &  n682 ) | ( n681  &  (~ n682) ) ;
 assign n684 = ( (~ n738)  &  n739 ) | ( n738  &  (~ n739) ) ;
 assign n685 = ( (~ n740)  &  n741 ) | ( n740  &  (~ n741) ) ;
 assign n683 = ( (~ n684)  &  n685 ) | ( n684  &  (~ n685) ) ;
 assign n686 = ( (~ n504)  &  n683 ) | ( n504  &  (~ n683) ) ;
 assign n688 = ( (~ P_2174_161_)  &  n677 ) | ( P_2174_161_  &  n794 ) | ( n677  &  n794 ) ;
 assign n687 = ( (~ n272)  &  n688 ) | ( n272  &  (~ n688) ) ;
 assign n690 = ( P_1497_156_  &  n680 ) | ( (~ P_1497_156_)  &  n686 ) | ( n680  &  n686 ) ;
 assign n689 = ( (~ n276)  &  n690 ) | ( n276  &  (~ n690) ) ;
 assign n692 = ( n800 ) | ( n801 ) | ( n796 ) | ( n799 ) ;
 assign n693 = ( (~ n735)  &  n861 ) | ( n735  &  (~ n861) ) ;
 assign n691 = ( (~ n692)  &  n693 ) | ( n692  &  (~ n693) ) ;
 assign n696 = ( P_335_123_  &  P_209_88_ ) | ( (~ P_335_123_)  &  P_206_87_ ) | ( P_209_88_  &  P_206_87_ ) ;
 assign n697 = ( P_335_123_  &  P_217_90_ ) | ( (~ P_335_123_)  &  P_210_89_ ) | ( P_217_90_  &  P_210_89_ ) ;
 assign n699 = ( P_332_122_  &  P_331_121_ ) | ( (~ P_332_122_)  &  P_324_120_ ) | ( P_331_121_  &  P_324_120_ ) ;
 assign n701 = ( (~ P_361_129_)  &  P_251_100_ ) | ( P_361_129_  &  P_248_99_ ) | ( P_251_100_  &  P_248_99_ ) ;
 assign n703 = ( (~ P_293_112_)  &  P_254_101_ ) | ( P_293_112_  &  P_242_97_ ) | ( P_254_101_  &  P_242_97_ ) ;
 assign n704 = ( (~ n312)  &  n360 ) | ( n313  &  n360 ) ;
 assign n705 = ( n526  &  (~ n550) ) | ( (~ n550)  &  (~ n727) ) ;
 assign n706 = ( (~ n172)  &  (~ n198) ) | ( (~ n198)  &  n609 ) ;
 assign n707 = ( (~ n200)  &  n266 ) | ( (~ n200)  &  n522 ) ;
 assign n709 = ( P_1690_158_  &  n809 ) | ( (~ P_1689_157_)  &  n809 ) | ( n280  &  n809 ) ;
 assign n710 = ( P_1694_160_  &  n810 ) | ( (~ P_1691_159_)  &  n810 ) | ( n280  &  n810 ) ;
 assign n711 = ( P_2358_162_  &  (~ P_25_8_) ) | ( (~ P_2358_162_)  &  (~ P_24_7_) ) | ( (~ P_25_8_)  &  (~ P_24_7_) ) ;
 assign n712 = ( P_2358_162_  &  (~ P_81_29_) ) | ( (~ P_2358_162_)  &  (~ P_26_9_) ) | ( (~ P_81_29_)  &  (~ P_26_9_) ) ;
 assign n713 = ( (~ P_2358_162_)  &  (~ P_79_27_) ) | ( P_2358_162_  &  (~ P_23_6_) ) | ( (~ P_79_27_)  &  (~ P_23_6_) ) ;
 assign n714 = ( (~ P_2358_162_)  &  (~ P_82_30_) ) | ( P_2358_162_  &  (~ P_80_28_) ) | ( (~ P_82_30_)  &  (~ P_80_28_) ) ;
 assign n715 = ( (~ P_54_20_)  &  n543 ) | ( P_54_20_  &  (~ n543) ) ;
 assign n716 = ( n160  &  n163 ) | ( (~ n160)  &  (~ n163) ) ;
 assign n717 = ( (~ P_3552_168_)  &  P_3546_165_ ) | ( (~ P_3552_168_)  &  P_514_147_ ) | ( P_3546_165_  &  (~ P_514_147_) ) ;
 assign n718 = ( n175  &  n182 ) | ( (~ n175)  &  (~ n182) ) ;
 assign n720 = ( (~ n501)  &  (~ n871) ) | ( n392  &  n582  &  (~ n871) ) ;
 assign n721 = ( (~ n390)  &  n768 ) | ( (~ n510)  &  (~ n581)  &  n768 ) ;
 assign n722 = ( (~ P_302_114_)  &  P_251_100_ ) | ( P_302_114_  &  P_248_99_ ) | ( P_251_100_  &  P_248_99_ ) ;
 assign n723 = ( n62  &  n66 ) | ( (~ n62)  &  (~ n66) ) ;
 assign n724 = ( (~ n668)  &  n190 ) | ( n668  &  (~ n190) ) ;
 assign n726 = ( n325 ) | ( n313 ) ;
 assign n727 = ( P_479_144_  &  n599 ) | ( (~ P_479_144_)  &  (~ n599) ) ;
 assign n725 = ( (~ n726)  &  n727 ) | ( n726  &  (~ n727) ) ;
 assign n728 = ( n158  &  n574 ) | ( (~ n158)  &  (~ n574) ) ;
 assign n730 = ( n157  &  n163 ) | ( (~ n157)  &  (~ n163) ) ;
 assign n731 = ( n460  &  n545 ) | ( (~ n460)  &  (~ n545) ) ;
 assign n732 = ( (~ n730)  &  n731 ) | ( n730  &  (~ n731) ) ;
 assign n734 = ( n552 ) | ( n471 ) ;
 assign n735 = ( (~ n70)  &  n78 ) | ( n70  &  (~ n78) ) ;
 assign n736 = ( (~ n675)  &  n171 ) | ( n675  &  (~ n171) ) ;
 assign n737 = ( (~ n673)  &  n521 ) | ( n673  &  (~ n521) ) ;
 assign n738 = ( n392  &  n510 ) | ( (~ n392)  &  (~ n510) ) ;
 assign n739 = ( (~ n183)  &  n180 ) | ( n183  &  (~ n180) ) ;
 assign n740 = ( (~ n175)  &  n501 ) | ( n175  &  (~ n501) ) ;
 assign n741 = ( (~ n390)  &  n391 ) | ( n390  &  (~ n391) ) ;
 assign n743 = ( (~ n185)  &  n389 ) | ( n185  &  (~ n389) ) ;
 assign n744 = ( (~ n175)  &  n504 ) | ( n175  &  (~ n504) ) ;
 assign n745 = ( (~ n390)  &  n501 ) | ( n390  &  (~ n501) ) ;
 assign n748 = ( n806  &  (~ n877) ) | ( (~ P_374_134_)  &  (~ n511)  &  (~ n877) ) ;
 assign n747 = ( n391  &  n748 ) | ( (~ n391)  &  (~ n748) ) ;
 assign n750 = ( n691 ) | ( n552 ) ;
 assign n753 = ( (~ P_316_118_)  &  P_308_116_ ) | ( P_316_118_  &  (~ P_308_116_) ) ;
 assign n754 = ( (~ P_210_89_)  &  P_218_91_ ) | ( P_210_89_  &  (~ P_218_91_) ) ;
 assign n755 = ( (~ n206)  &  n599 ) | ( n206  &  (~ n599) ) ;
 assign n758 = ( P_335_123_  &  P_264_103_ ) | ( (~ P_335_123_)  &  P_257_102_ ) | ( P_264_103_  &  P_257_102_ ) ;
 assign n757 = ( (~ n211)  &  n758 ) | ( n211  &  (~ n758) ) ;
 assign n760 = ( P_335_123_  &  P_272_105_ ) | ( (~ P_335_123_)  &  P_265_104_ ) | ( P_272_105_  &  P_265_104_ ) ;
 assign n761 = ( P_335_123_  &  P_280_107_ ) | ( (~ P_335_123_)  &  P_273_106_ ) | ( P_280_107_  &  P_273_106_ ) ;
 assign n762 = ( P_335_123_  &  P_225_92_ ) | ( (~ P_335_123_)  &  P_218_91_ ) | ( P_225_92_  &  P_218_91_ ) ;
 assign n766 = ( n569 ) | ( n574 ) | ( n545 ) ;
 assign n768 = ( n510 ) | ( n581 ) | ( n390 ) ;
 assign n770 = ( n187  &  n315 ) | ( (~ n187)  &  (~ n315) ) ;
 assign n771 = ( n188  &  n315 ) | ( (~ n188)  &  (~ n315) ) ;
 assign n773 = ( (~ n726)  &  n312 ) | ( n726  &  (~ n312) ) ;
 assign n778 = ( P_514_147_  &  P_248_99_ ) | ( (~ P_514_147_)  &  (~ P_242_97_) ) | ( P_248_99_  &  (~ P_242_97_) ) ;
 assign n779 = ( (~ n38)  &  n50 ) | ( n38  &  (~ n50) ) ;
 assign n781 = ( (~ n58)  &  n778 ) | ( n58  &  (~ n778) ) ;
 assign n780 = ( n701  &  (~ n779)  &  n781 ) ;
 assign n783 = ( (~ n701)  &  n779  &  n781 ) ;
 assign n784 = ( n701  &  n779  &  (~ n781) ) ;
 assign n786 = ( (~ n701)  &  (~ n779)  &  (~ n781) ) ;
 assign n787 = ( (~ n162) ) | ( n634 ) ;
 assign n789 = ( (~ P_2174_161_) ) | ( n273 ) | ( (~ n787) ) ;
 assign n788 = ( n312  &  n860 ) | ( (~ n312)  &  (~ n860) ) ;
 assign n790 = ( (~ n728)  &  n846 ) | ( n728  &  (~ n846) ) ;
 assign n791 = ( (~ n570) ) | ( n623 ) ;
 assign n793 = ( n558 ) | ( n574 ) | ( (~ n791) ) ;
 assign n792 = ( n791  &  n793 ) | ( (~ n558)  &  (~ n574)  &  n793 ) ;
 assign n794 = ( (~ n732)  &  n847 ) | ( n732  &  (~ n847) ) ;
 assign n796 = ( (~ n126)  &  (~ n465)  &  (~ n466) ) ;
 assign n799 = ( n126  &  (~ n465)  &  n466 ) ;
 assign n800 = ( (~ n126)  &  n465  &  n466 ) ;
 assign n801 = ( n126  &  n465  &  (~ n466) ) ;
 assign n802 = ( n633  &  n174 ) ;
 assign n805 = ( (~ P_1497_156_) ) | ( n277 ) | ( n802 ) ;
 assign n803 = ( (~ n172)  &  n862 ) | ( n172  &  (~ n862) ) ;
 assign n806 = ( n626  &  n180 ) ;
 assign n809 = ( (~ P_1690_158_) ) | ( (~ P_1689_157_) ) | ( (~ P_179_78_) ) ;
 assign n810 = ( (~ P_1694_160_) ) | ( (~ P_1691_159_) ) | ( (~ P_179_78_) ) ;
 assign n819 = ( P_351_127_  &  P_341_125_ ) | ( (~ P_351_127_)  &  (~ P_341_125_) ) ;
 assign n820 = ( P_324_120_  &  n474  &  (~ n819) ) ;
 assign n822 = ( P_324_120_  &  (~ n474)  &  n819 ) ;
 assign n824 = ( (~ P_324_120_)  &  n474  &  n819 ) ;
 assign n825 = ( (~ P_324_120_)  &  (~ n474)  &  (~ n819) ) ;
 assign n826 = ( P_273_106_  &  P_265_104_ ) | ( (~ P_273_106_)  &  (~ P_265_104_) ) ;
 assign n827 = ( n478  &  n480  &  (~ n826) ) ;
 assign n829 = ( n478  &  (~ n480)  &  n826 ) ;
 assign n831 = ( (~ n478)  &  n480  &  n826 ) ;
 assign n833 = ( (~ n478)  &  (~ n480)  &  (~ n826) ) ;
 assign n835 = ( (~ n530)  &  n538 ) | ( n530  &  (~ n538) ) ;
 assign n837 = ( n697  &  n762 ) | ( (~ n697)  &  (~ n762) ) ;
 assign n839 = ( P_3724_170_  &  n666 ) | ( (~ P_3724_170_)  &  n703 ) | ( n666  &  n703 ) ;
 assign n840 = ( (~ P_3724_170_)  &  P_123_53_ ) | ( P_3724_170_  &  (~ P_623_2152_) ) | ( P_123_53_  &  (~ P_623_2152_) ) ;
 assign n844 = ( (~ n179)  &  n504 ) | ( n179  &  (~ n504) ) ;
 assign n846 = ( n543  &  n570 ) | ( (~ n543)  &  (~ n570) ) ;
 assign n847 = ( (~ n792)  &  n868 ) | ( n792  &  (~ n868) ) ;
 assign n848 = ( n541  &  n699 ) | ( (~ n541)  &  (~ n699) ) ;
 assign n849 = ( (~ n312)  &  n549 ) ;
 assign n850 = ( n824 ) | ( n825 ) | ( n820 ) | ( n822 ) ;
 assign n851 = ( n831 ) | ( n833 ) | ( n827 ) | ( n829 ) ;
 assign n852 = ( n520 ) | ( n633 ) ;
 assign n859 = ( (~ n703)  &  n722 ) | ( n703  &  (~ n722) ) ;
 assign n860 = ( n259  &  n315 ) | ( (~ n259)  &  (~ n315) ) ;
 assign n861 = ( (~ n94)  &  n138 ) | ( n94  &  (~ n138) ) ;
 assign n862 = ( (~ n264)  &  n521 ) | ( n264  &  (~ n521) ) ;
 assign n867 = ( n548  &  n315 ) | ( (~ n548)  &  (~ n315) ) ;
 assign n868 = ( n204  &  n543 ) | ( (~ n204)  &  (~ n543) ) ;
 assign n869 = ( (~ n172)  &  n266 ) | ( n172  &  (~ n266) ) ;
 assign n871 = ( n392  &  (~ n501)  &  n582 ) ;
 assign n877 = ( (~ P_374_134_)  &  (~ n511)  &  n806 ) ;
 assign P_993_850_ = ( P_1_0_ ) ;
 assign P_978_851_ = ( P_1_0_ ) ;
 assign P_973_202_ = ( P_3173_164_ ) ;
 assign P_949_852_ = ( P_1_0_ ) ;
 assign P_939_853_ = ( P_1_0_ ) ;
 assign P_926_624_ = ( P_137_63_ ) ;
 assign P_923_619_ = ( P_141_65_ ) ;
 assign P_921_664_ = ( P_1_0_ ) ;
 assign P_892_408_ = ( P_549_151_ ) ;
 assign P_889_734_ = ( P_299_113_ ) ;
 assign P_887_528_ = ( P_299_113_ ) ;
 assign P_629_1926_ = ( wire102 ) ;
 assign P_626_1752_ = ( wire103 ) ;
 assign P_618_1925_ = ( wire102 ) ;
 assign P_615_1750_ = ( wire103 ) ;
 assign P_298_299_ = ( P_293_112_ ) ;
 assign P_144_354_ = ( P_141_65_ ) ;


endmodule

