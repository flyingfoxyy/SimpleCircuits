module pair (
	Pz4, Pz3, Pz2, Pz1, Pz0, Pz, Py4, Py3, 
	Py2, Py1, Py0, Py, Px4, Px3, Px2, Px1, Px0, Pw4, 
	Pw3, Pw2, Pw1, Pw0, Pw, Pv4, Pv3, Pv2, Pv1, Pv0, 
	Pv, Pu4, Pu3, Pu2, Pu1, Pu0, Pu, Pt4, Pt3, Pt2, 
	Pt1, Pt0, Pt, Ps4, Ps3, Ps2, Ps1, Ps0, Ps, Pr5, 
	Pr4, Pr3, Pr2, Pr1, Pr0, Pr, Pq5, Pq4, Pq3, Pq2, 
	Pq1, Pq0, Pq, Pp5, Pp4, Pp3, Pp2, Pp1, Pp0, Pp, 
	Po5, Po4, Po3, Po2, Po1, Po0, Po, Pn5, Pn4, Pn3, 
	Pn2, Pn1, Pn0, Pn, Pm5, Pm4, Pm3, Pm2, Pm1, Pm0, 
	Pm, Pl5, Pl4, Pl3, Pl2, Pl1, Pl0, Pl, Pk5, Pk4, 
	Pk3, Pk2, Pk1, Pk0, Pk, Pj5, Pj4, Pj3, Pj2, Pj1, 
	Pj0, Pj, Pi5, Pi4, Pi3, Pi2, Pi1, Pi0, Pi, Ph5, 
	Ph4, Ph3, Ph2, Ph1, Ph0, Ph, Pg5, Pg4, Pg3, Pg2, 
	Pg1, Pg0, Pg, Pf5, Pf4, Pf3, Pf2, Pf1, Pf0, Pf, 
	Pe5, Pe4, Pe3, Pe2, Pe1, Pe0, Pe, Pd5, Pd4, Pd3, 
	Pd2, Pd1, Pd0, Pd, Pc5, Pc4, Pc3, Pc2, Pc1, Pc0, 
	Pc, Pb5, Pb4, Pb3, Pb2, Pb1, Pb0, Pb, Pa5, Pa4, 
	Pa3, Pa2, Pa1, Pa0, Pa, Pz9, Pz8, Pz7, Pz6, Pz5, 
	Py10, Py9, Py8, Py7, Py6, Py5, Px10, Px9, Px8, Px7, 
	Px6, Px5, Pw10, Pw9, Pw8, Pw7, Pw6, Pw5, Pv10, Pv9, 
	Pv8, Pv7, Pv6, Pv5, Pu10, Pu9, Pu8, Pu7, Pu6, Pu5, 
	Pt10, Pt9, Pt8, Pt7, Pt6, Pt5, Ps10, Ps9, Ps8, Ps7, 
	Ps6, Ps5, Pr10, Pr9, Pr8, Pr7, Pr6, Pq10, Pq9, Pq8, 
	Pq7, Pq6, Pp10, Pp9, Pp8, Pp7, Pp6, Po10, Po9, Po8, 
	Po7, Po6, Pn10, Pn9, Pn8, Pn7, Pn6, Pm10, Pm9, Pm8, 
	Pm7, Pm6, Pl10, Pl9, Pl8, Pl7, Pl6, Pk10, Pk9, Pk8, 
	Pk7, Pk6, Pj10, Pj9, Pj8, Pj7, Pj6, Pi10, Pi9, Pi8, 
	Pi7, Pi6, Ph10, Ph9, Ph8, Ph7, Ph6, Pg10, Pg9, Pg8, 
	Pg7, Pg6, Pf10, Pf9, Pf8, Pf7, Pf6, Pe10, Pe9, Pe8, 
	Pe7, Pe6, Pd10, Pd9, Pd8, Pd7, Pd6, Pc10, Pc9, Pc8, 
	Pc7, Pc6, Pb10, Pb9, Pb8, Pb7, Pb6, Pa10, Pa9, Pa8, 
	Pa7, Pa6);

input Pz4, Pz3, Pz2, Pz1, Pz0, Pz, Py4, Py3, Py2, Py1, Py0, Py, Px4, Px3, Px2, Px1, Px0, Pw4, Pw3, Pw2, Pw1, Pw0, Pw, Pv4, Pv3, Pv2, Pv1, Pv0, Pv, Pu4, Pu3, Pu2, Pu1, Pu0, Pu, Pt4, Pt3, Pt2, Pt1, Pt0, Pt, Ps4, Ps3, Ps2, Ps1, Ps0, Ps, Pr5, Pr4, Pr3, Pr2, Pr1, Pr0, Pr, Pq5, Pq4, Pq3, Pq2, Pq1, Pq0, Pq, Pp5, Pp4, Pp3, Pp2, Pp1, Pp0, Pp, Po5, Po4, Po3, Po2, Po1, Po0, Po, Pn5, Pn4, Pn3, Pn2, Pn1, Pn0, Pn, Pm5, Pm4, Pm3, Pm2, Pm1, Pm0, Pm, Pl5, Pl4, Pl3, Pl2, Pl1, Pl0, Pl, Pk5, Pk4, Pk3, Pk2, Pk1, Pk0, Pk, Pj5, Pj4, Pj3, Pj2, Pj1, Pj0, Pj, Pi5, Pi4, Pi3, Pi2, Pi1, Pi0, Pi, Ph5, Ph4, Ph3, Ph2, Ph1, Ph0, Ph, Pg5, Pg4, Pg3, Pg2, Pg1, Pg0, Pg, Pf5, Pf4, Pf3, Pf2, Pf1, Pf0, Pf, Pe5, Pe4, Pe3, Pe2, Pe1, Pe0, Pe, Pd5, Pd4, Pd3, Pd2, Pd1, Pd0, Pd, Pc5, Pc4, Pc3, Pc2, Pc1, Pc0, Pc, Pb5, Pb4, Pb3, Pb2, Pb1, Pb0, Pb, Pa5, Pa4, Pa3, Pa2, Pa1, Pa0, Pa;

output Pz9, Pz8, Pz7, Pz6, Pz5, Py10, Py9, Py8, Py7, Py6, Py5, Px10, Px9, Px8, Px7, Px6, Px5, Pw10, Pw9, Pw8, Pw7, Pw6, Pw5, Pv10, Pv9, Pv8, Pv7, Pv6, Pv5, Pu10, Pu9, Pu8, Pu7, Pu6, Pu5, Pt10, Pt9, Pt8, Pt7, Pt6, Pt5, Ps10, Ps9, Ps8, Ps7, Ps6, Ps5, Pr10, Pr9, Pr8, Pr7, Pr6, Pq10, Pq9, Pq8, Pq7, Pq6, Pp10, Pp9, Pp8, Pp7, Pp6, Po10, Po9, Po8, Po7, Po6, Pn10, Pn9, Pn8, Pn7, Pn6, Pm10, Pm9, Pm8, Pm7, Pm6, Pl10, Pl9, Pl8, Pl7, Pl6, Pk10, Pk9, Pk8, Pk7, Pk6, Pj10, Pj9, Pj8, Pj7, Pj6, Pi10, Pi9, Pi8, Pi7, Pi6, Ph10, Ph9, Ph8, Ph7, Ph6, Pg10, Pg9, Pg8, Pg7, Pg6, Pf10, Pf9, Pf8, Pf7, Pf6, Pe10, Pe9, Pe8, Pe7, Pe6, Pd10, Pd9, Pd8, Pd7, Pd6, Pc10, Pc9, Pc8, Pc7, Pc6, Pb10, Pb9, Pb8, Pb7, Pb6, Pa10, Pa9, Pa8, Pa7, Pa6;

wire n13, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n31, n32, n33, n34, n30, n35, n38, n36, n39, n43, n42, n45, n44, n47, n46, n48, n49, n50, n52, n51, n53, n54, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n76, n74, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n94, n92, n96, n97, n98, n99, n100, n101, n102, n103, n104, n107, n106, n110, n109, n112, n111, n113, n114, n115, n117, n116, n118, n119, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n136, n137, n138, n139, n140, n141, n142, n143, n144, n147, n145, n146, n150, n151, n152, n153, n154, n155, n156, n159, n160, n161, n158, n163, n166, n164, n167, n172, n169, n173, n176, n182, n179, n184, n183, n186, n185, n187, n191, n190, n195, n192, n198, n197, n201, n206, n207, n205, n203, n208, n211, n214, n213, n219, n217, n221, n220, n222, n227, n225, n229, n230, n228, n233, n231, n235, n236, n237, n234, n239, n240, n238, n241, n246, n247, n248, n245, n249, n253, n252, n254, n260, n257, n263, n262, n265, n266, n264, n267, n269, n270, n271, n268, n273, n274, n272, n275, n277, n276, n278, n282, n284, n285, n286, n287, n288, n289, n283, n291, n290, n293, n292, n294, n298, n295, n301, n299, n300, n303, n304, n305, n302, n307, n306, n308, n310, n311, n313, n314, n315, n312, n318, n320, n319, n322, n321, n324, n323, n326, n325, n329, n332, n333, n334, n331, n336, n335, n339, n341, n340, n343, n342, n344, n345, n348, n349, n350, n347, n351, n352, n355, n354, n357, n356, n359, n361, n360, n363, n362, n365, n364, n369, n367, n368, n366, n370, n372, n371, n374, n373, n375, n377, n376, n378, n380, n379, n381, n383, n382, n387, n384, n390, n389, n393, n396, n395, n401, n399, n403, n402, n404, n405, n406, n407, n410, n408, n411, n414, n413, n415, n422, n419, n424, n423, n426, n427, n425, n429, n428, n430, n431, n433, n434, n432, n436, n437, n435, n438, n439, n442, n441, n443, n450, n447, n452, n451, n454, n453, n455, n457, n456, n459, n460, n458, n462, n461, n464, n465, n463, n466, n468, n467, n470, n471, n469, n473, n472, n474, n476, n477, n475, n479, n478, n480, n482, n481, n484, n485, n486, n487, n488, n489, n483, n490, n492, n493, n491, n495, n497, n498, n499, n496, n500, n501, n503, n506, n508, n510, n514, n515, n517, n531, n532, n538, n541, n543, n544, n566, n568, n573, n575, n578, n581, n588, n609, n611, n617, n624, n625, n626, n627, n628, n629, n631, n632, n633, n636, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n681, n682, n683, n684, n685, n686, n687, n689, n690, n691, n692, n693, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n720, n722, n723, n724, n725, n726, n727, n728, n729, n733, n734, n735, n738, n741, n742, n743, n744, n745, n746, n747, n749, n748, n750, n751, n753, n752, n754, n755, n759, n760, n763, n764;

assign Pz9 = ( n136  &  (~ n515) ) ;
 assign Pz8 = ( (~ n103) ) ;
 assign Pz7 = ( n72  &  n70 ) ;
 assign Pz6 = ( (~ Pb)  &  n43  &  n42 ) | ( (~ Pb)  &  n43  &  (~ n169) ) ;
 assign Pz5 = ( (~ n234) ) ;
 assign Py10 = ( n166  &  (~ n679) ) | ( Pp5  &  n166  &  n164 ) ;
 assign Py9 = ( n134  &  (~ n515) ) ;
 assign Py8 = ( n102  &  n88 ) ;
 assign Py7 = ( n70  &  n71 ) ;
 assign Py6 = ( n38  &  (~ n674) ) | ( Pp1  &  n38  &  n36 ) ;
 assign Py5 = ( (~ n245) ) ;
 assign Px10 = ( n166  &  (~ n686) ) | ( Pr5  &  n166  &  n164 ) ;
 assign Px9 = ( (~ n133) ) ;
 assign Px8 = ( (~ n101) ) ;
 assign Px7 = ( n69  &  n70 ) ;
 assign Px6 = ( n38  &  (~ n681) ) | ( Pr1  &  n38  &  n36 ) ;
 assign Px5 = ( (~ n268) ) ;
 assign Pw10 = ( (~ n163) ) ;
 assign Pw9 = ( Pq4  &  Pm4  &  Pl4  &  Ph4  &  Po4  &  Pk4  &  n132  &  Pn4 ) ;
 assign Pw8 = ( (~ n100) ) ;
 assign Pw7 = ( (~ n658) ) ;
 assign Pw6 = ( (~ n35) ) ;
 assign Pw5 = ( (~ n283) ) ;
 assign Pv10 = ( (~ n94) ) ;
 assign Pv9 = ( (~ n131) ) ;
 assign Pv8 = ( (~ n99) ) ;
 assign Pv7 = ( (~ n68) ) ;
 assign Pv6 = ( (~ n76) ) ;
 assign Pv5 = ( (~ n302) ) ;
 assign Pu10 = ( (~ n158) ) ;
 assign Pu9 = ( (~ n130) ) ;
 assign Pu8 = ( n88  &  n98 ) ;
 assign Pu7 = ( Po2  &  Pm2  &  Pl2  &  Pk2  &  Pi2  &  Pj2  &  n67  &  Pf2 ) ;
 assign Pu6 = ( (~ n30) ) ;
 assign Pu5 = ( (~ n312) ) ;
 assign Pt10 = ( (~ Pz)  &  n155 ) | ( (~ Pz)  &  n156 ) | ( (~ Pz)  &  (~ n704) ) ;
 assign Pt9 = ( (~ n129) ) ;
 assign Pt8 = ( n97  &  n88 ) ;
 assign Pt7 = ( (~ n66) ) ;
 assign Pt6 = ( (~ Pb)  &  n26 ) | ( (~ Pb)  &  n27 ) | ( (~ Pb)  &  (~ n699) ) ;
 assign Pt5 = ( (~ n331) ) ;
 assign Ps10 = ( (~ n154) ) ;
 assign Ps9 = ( (~ n128) ) ;
 assign Ps8 = ( n96  &  n88 ) ;
 assign Ps7 = ( (~ n65) ) ;
 assign Ps6 = ( (~ n25) ) ;
 assign Ps5 = ( (~ n347) ) ;
 assign Pr10 = ( n151  &  n153 ) ;
 assign Pr9 = ( (~ n127) ) ;
 assign Pr8 = ( Pn3  &  n88  &  Po3  &  Pm3  &  Pl3 ) ;
 assign Pr7 = ( (~ n64) ) ;
 assign Pq10 = ( n151  &  n152 ) ;
 assign Pq9 = ( (~ n126) ) ;
 assign Pq8 = ( (~ n659) ) ;
 assign Pq7 = ( (~ n63) ) ;
 assign Pq6 = ( (~ n24) ) ;
 assign Pp9 = ( Pz ) | ( n125 ) ;
 assign Pp8 = ( (~ n91) ) ;
 assign Pp7 = ( (~ n62) ) ;
 assign Pp6 = ( (~ n660) ) ;
 assign Po10 = ( (~ n150) ) ;
 assign Po9 = ( (~ n124) ) ;
 assign Po8 = ( n90  &  n88 ) ;
 assign Po7 = ( (~ n61) ) ;
 assign Po6 = ( (~ n661) ) ;
 assign Pn10 = ( (~ Pz)  &  (~ n147) ) | ( (~ Pz)  &  (~ n662) ) ;
 assign Pn9 = ( (~ n123) ) ;
 assign Pn8 = ( n88  &  n89 ) ;
 assign Pn7 = ( Pb ) | ( n60 ) ;
 assign Pn6 = ( n23 ) | ( Pi1 ) ;
 assign Pm10 = ( n147  &  n145 ) | ( n147  &  n146 ) | ( n147  &  Pz ) ;
 assign Pm9 = ( Pz ) | ( n122 ) ;
 assign Pm8 = ( n87  &  n88 ) ;
 assign Pm7 = ( (~ n59) ) ;
 assign Pl10 = ( (~ n663) ) ;
 assign Pl9 = ( Pz ) | ( n121 ) ;
 assign Pl8 = ( (~ n86) ) ;
 assign Pl7 = ( (~ n58) ) ;
 assign Pk10 = ( (~ n664) ) ;
 assign Pk9 = ( Pz ) | ( (~ Pd4) ) ;
 assign Pk8 = ( (~ n85) ) ;
 assign Pk7 = ( Pb ) | ( n57 ) ;
 assign Pk6 = ( n22  &  (~ n633) ) ;
 assign Pj10 = ( n144 ) | ( Pe5 ) ;
 assign Pj9 = ( (~ n119) ) ;
 assign Pj8 = ( n84  &  n70 ) ;
 assign Pj7 = ( Pb ) | ( n56 ) ;
 assign Pj6 = ( n21  &  (~ n633) ) ;
 assign Pi9 = ( (~ n118) ) ;
 assign Pi8 = ( (~ n83) ) ;
 assign Pi7 = ( (~ Pb2) ) | ( Pb ) ;
 assign Pi6 = ( n20  &  (~ n633) ) ;
 assign Ph9 = ( (~ Pz)  &  n117  &  n116 ) | ( (~ Pz)  &  n117  &  (~ n179) ) ;
 assign Ph8 = ( (~ n82) ) ;
 assign Ph7 = ( (~ n54) ) ;
 assign Ph6 = ( n19  &  (~ n633) ) ;
 assign Pg10 = ( n143  &  (~ n515) ) ;
 assign Pg9 = ( (~ n115) ) ;
 assign Pg8 = ( (~ n81) ) ;
 assign Pg7 = ( (~ n53) ) ;
 assign Pg6 = ( n18  &  (~ n633) ) ;
 assign Pf10 = ( n142  &  (~ n515) ) ;
 assign Pf9 = ( (~ n114) ) ;
 assign Pf8 = ( n70  &  n80 ) ;
 assign Pf7 = ( (~ Pb)  &  n52  &  n51 ) | ( (~ Pb)  &  n52  &  (~ n169) ) ;
 assign Pf6 = ( n17  &  (~ n633) ) ;
 assign Pe10 = ( n141  &  (~ n515) ) ;
 assign Pe9 = ( (~ n113) ) ;
 assign Pe8 = ( n79  &  n70 ) ;
 assign Pe7 = ( (~ n50) ) ;
 assign Pe6 = ( n16  &  (~ n633) ) ;
 assign Pd10 = ( n140  &  (~ n515) ) ;
 assign Pd9 = ( (~ Pz)  &  n112  &  n111 ) | ( (~ Pz)  &  n112  &  (~ n179) ) ;
 assign Pd8 = ( n78  &  n70 ) ;
 assign Pd7 = ( (~ n49) ) ;
 assign Pd6 = ( n15  &  (~ n633) ) ;
 assign Pc10 = ( n139  &  (~ n515) ) ;
 assign Pc9 = ( (~ Pz)  &  n110  &  n109 ) | ( (~ Pz)  &  n110  &  (~ n179) ) ;
 assign Pc8 = ( Pw2  &  n70  &  Py2  &  Pz2  &  Px2 ) ;
 assign Pc7 = ( (~ n48) ) ;
 assign Pc6 = ( n13  &  (~ n633) ) ;
 assign Pb10 = ( n138  &  (~ n515) ) ;
 assign Pb9 = ( (~ Pz)  &  n107  &  n106 ) | ( (~ Pz)  &  n107  &  (~ n179) ) ;
 assign Pb8 = ( (~ n665) ) ;
 assign Pb7 = ( (~ Pb)  &  n47  &  n46 ) | ( (~ Pb)  &  n47  &  (~ n169) ) ;
 assign Pb6 = ( (~ n483) ) ;
 assign Pa10 = ( n137  &  (~ n515) ) ;
 assign Pa9 = ( (~ n104) ) ;
 assign Pa8 = ( (~ n73) ) ;
 assign Pa7 = ( (~ Pb)  &  n45  &  n44 ) | ( (~ Pb)  &  n45  &  (~ n169) ) ;
 assign Pa6 = ( (~ n496) ) ;
 assign n13 = ( Pv0  &  n323 ) | ( (~ Pv0)  &  (~ n323) ) ;
 assign n15 = ( Pw0  &  n639 ) | ( (~ Pw0)  &  (~ n639) ) ;
 assign n16 = ( Px0  &  n640 ) | ( (~ Px0)  &  (~ n640) ) ;
 assign n17 = ( Py0  &  n653 ) | ( (~ Py0)  &  (~ n653) ) ;
 assign n18 = ( Pz0  &  n624 ) | ( (~ Pz0)  &  (~ n624) ) ;
 assign n19 = ( Pa1  &  n625 ) | ( (~ Pa1)  &  (~ n625) ) ;
 assign n20 = ( Pb1  &  n648 ) | ( (~ Pb1)  &  (~ n648) ) ;
 assign n21 = ( Pc1  &  n626 ) | ( (~ Pc1)  &  (~ n626) ) ;
 assign n22 = ( Pd1  &  n326 ) | ( (~ Pd1)  &  (~ n326) ) ;
 assign n23 = ( (~ Ph1)  &  (~ n310)  &  n538 ) ;
 assign n24 = ( n365  &  n172  &  Pb ) | ( n365  &  n172  &  n364 ) ;
 assign n25 = ( n32  &  n310  &  (~ n344) ) | ( n32  &  (~ n344)  &  n345 ) ;
 assign n26 = ( (~ n308)  &  n310 ) | ( (~ n308)  &  n329 ) ;
 assign n27 = ( Pn1  &  Pm1 ) ;
 assign n31 = ( n308 ) | ( n310 ) | ( n311 ) ;
 assign n32 = ( n172  &  n308 ) | ( n172  &  (~ n329) ) ;
 assign n33 = ( (~ Pn1) ) | ( (~ Pm1) ) | ( n531 ) ;
 assign n34 = ( (~ Pn1) ) | ( Pm1 ) | ( Pl1 ) | ( Pb ) ;
 assign n30 = ( n31  &  n32  &  n33  &  n34 ) ;
 assign n35 = ( (~ Pr1)  &  n38  &  n282 ) | ( n38  &  n282  &  (~ n566) ) ;
 assign n38 = ( n39  &  Pr1 ) | ( n39  &  Pp1 ) | ( n39  &  Pq1 ) ;
 assign n36 = ( Pd ) | ( (~ n34) ) ;
 assign n39 = ( (~ Pb)  &  n241 ) | ( (~ Pq1)  &  (~ Pp1)  &  (~ Pb) ) ;
 assign n43 = ( n169 ) | ( Pw2 ) ;
 assign n42 = ( Ps1  &  n173 ) | ( (~ Ps1)  &  (~ n173) ) ;
 assign n45 = ( n169 ) | ( Px2 ) ;
 assign n44 = ( Pt1  &  n755 ) | ( (~ Pt1)  &  (~ n755) ) ;
 assign n47 = ( n169 ) | ( Py2 ) ;
 assign n46 = ( Pu1  &  n752 ) | ( (~ Pu1)  &  (~ n752) ) ;
 assign n48 = ( (~ Pb)  &  (~ n169)  &  n482 ) | ( (~ Pb)  &  n482  &  n481 ) ;
 assign n49 = ( (~ Pb)  &  (~ n169)  &  n479 ) | ( (~ Pb)  &  n479  &  n478 ) ;
 assign n50 = ( (~ Pb)  &  (~ n169)  &  n473 ) | ( (~ Pb)  &  n473  &  n472 ) ;
 assign n52 = ( n169 ) | ( Pc3 ) ;
 assign n51 = ( Py1  &  n463 ) | ( (~ Py1)  &  (~ n463) ) ;
 assign n53 = ( (~ Pb)  &  (~ n169)  &  n457 ) | ( (~ Pb)  &  n457  &  n456 ) ;
 assign n54 = ( (~ Pb)  &  (~ n169)  &  n452 ) | ( (~ Pb)  &  n452  &  n451 ) ;
 assign n56 = ( (~ Pc2)  &  Pb2 ) | ( Pc2  &  (~ Pb2) ) ;
 assign n57 = ( (~ Pd2)  &  n405 ) | ( Pd2  &  (~ n405) ) ;
 assign n58 = ( (~ Pb)  &  n299  &  n403 ) | ( (~ Pb)  &  n403  &  n402 ) ;
 assign n59 = ( (~ Pb)  &  n299  &  n383 ) | ( (~ Pb)  &  n383  &  n382 ) ;
 assign n60 = ( Pg2  &  n276 ) | ( (~ Pg2)  &  (~ n276) ) ;
 assign n61 = ( (~ Pb)  &  n299  &  n377 ) | ( (~ Pb)  &  n377  &  n376 ) ;
 assign n62 = ( (~ Pb)  &  n299  &  n372 ) | ( (~ Pb)  &  n372  &  n371 ) ;
 assign n63 = ( (~ Pb)  &  n299  &  n363 ) | ( (~ Pb)  &  n363  &  n362 ) ;
 assign n64 = ( (~ Pb)  &  n299  &  n357 ) | ( (~ Pb)  &  n357  &  n356 ) ;
 assign n65 = ( (~ Pb)  &  n299  &  n343 ) | ( (~ Pb)  &  n343  &  n342 ) ;
 assign n66 = ( (~ Pb)  &  n299  &  n322 ) | ( (~ Pb)  &  n322  &  n321 ) ;
 assign n67 = ( Ph2  &  Pb ) | ( Ph2  &  (~ n299) ) ;
 assign n68 = ( (~ Pb)  &  n301  &  n299 ) | ( (~ Pb)  &  n301  &  n300 ) ;
 assign n69 = ( Pq2  &  n225 ) | ( (~ Pq2)  &  (~ n225) ) ;
 assign n70 = ( (~ Pb)  &  n345 ) ;
 assign n71 = ( Pr2  &  n715 ) | ( (~ Pr2)  &  (~ n715) ) ;
 assign n72 = ( Ps2  &  n228 ) | ( (~ Ps2)  &  (~ n228) ) ;
 assign n73 = ( (~ n70)  &  n401 ) | ( n401  &  n495 ) ;
 assign n76 = ( Pn1  &  (~ Pb) ) | ( Pm1  &  (~ Pb) ) | ( Pl1  &  (~ Pb) ) ;
 assign n74 = ( (~ Pg)  &  n76 ) | ( (~ Pg)  &  (~ n543) ) ;
 assign n78 = ( Pw2  &  n474 ) | ( (~ Pw2)  &  (~ n474) ) ;
 assign n79 = ( Px2  &  n469 ) | ( (~ Px2)  &  (~ n469) ) ;
 assign n80 = ( Py2  &  n746 ) | ( (~ Py2)  &  (~ n746) ) ;
 assign n81 = ( (~ n70)  &  n401 ) | ( n401  &  n455 ) ;
 assign n82 = ( (~ n70)  &  n401 ) | ( n401  &  n438 ) ;
 assign n83 = ( (~ n70)  &  n401 ) | ( n401  &  n431 ) ;
 assign n84 = ( Pc3  &  n425 ) | ( (~ Pc3)  &  (~ n425) ) ;
 assign n85 = ( (~ n70)  &  n401 ) | ( n401  &  n404 ) ;
 assign n86 = ( (~ n70)  &  n401 ) | ( n401  &  n399 ) ;
 assign n87 = ( (~ Pf3)  &  n369 ) | ( Pf3  &  (~ n369) ) ;
 assign n88 = ( (~ Pz)  &  n352 ) ;
 assign n89 = ( Pg3  &  n735 ) | ( (~ Pg3)  &  (~ n735) ) ;
 assign n90 = ( Ph3  &  n375 ) | ( (~ Ph3)  &  (~ n375) ) ;
 assign n91 = ( (~ n88)  &  n219 ) | ( n219  &  n370 ) ;
 assign n94 = ( (~ Pz)  &  Pn5 ) | ( (~ Pz)  &  Pm5 ) | ( (~ Pz)  &  Pl5 ) ;
 assign n92 = ( (~ Pe0)  &  n94 ) | ( (~ Pe0)  &  (~ n205) ) ;
 assign n96 = ( Pl3  &  n760 ) | ( (~ Pl3)  &  (~ n760) ) ;
 assign n97 = ( Pm3  &  n759 ) | ( (~ Pm3)  &  (~ n759) ) ;
 assign n98 = ( Pn3  &  n724 ) | ( (~ Pn3)  &  (~ n724) ) ;
 assign n99 = ( (~ n88)  &  n219 ) | ( n219  &  n294 ) ;
 assign n100 = ( (~ n88)  &  n219 ) | ( n219  &  n275 ) ;
 assign n101 = ( (~ n88)  &  n219 ) | ( n219  &  n267 ) ;
 assign n102 = ( Pr3  &  n238 ) | ( (~ Pr3)  &  (~ n238) ) ;
 assign n103 = ( (~ n88)  &  n219 ) | ( n219  &  n217 ) ;
 assign n104 = ( (~ n88)  &  n219 ) | ( n219  &  n490 ) ;
 assign n107 = ( Pl3 ) | ( n179 ) ;
 assign n106 = ( Pu3  &  n176 ) | ( (~ Pu3)  &  (~ n176) ) ;
 assign n110 = ( Pm3 ) | ( n179 ) ;
 assign n109 = ( Pv3  &  n750 ) | ( (~ Pv3)  &  (~ n750) ) ;
 assign n112 = ( Pn3 ) | ( n179 ) ;
 assign n111 = ( Pw3  &  n748 ) | ( (~ Pw3)  &  (~ n748) ) ;
 assign n113 = ( (~ Pz)  &  (~ n179)  &  n468 ) | ( (~ Pz)  &  n468  &  n467 ) ;
 assign n114 = ( (~ Pz)  &  (~ n179)  &  n462 ) | ( (~ Pz)  &  n462  &  n461 ) ;
 assign n115 = ( (~ Pz)  &  (~ n179)  &  n454 ) | ( (~ Pz)  &  n454  &  n453 ) ;
 assign n117 = ( Pr3 ) | ( n179 ) ;
 assign n116 = ( Pa4  &  n432 ) | ( (~ Pa4)  &  (~ n432) ) ;
 assign n118 = ( (~ Pz)  &  (~ n179)  &  n429 ) | ( (~ Pz)  &  n429  &  n428 ) ;
 assign n119 = ( (~ Pz)  &  (~ n179)  &  n424 ) | ( (~ Pz)  &  n424  &  n423 ) ;
 assign n121 = ( (~ Pe4)  &  Pd4 ) | ( Pe4  &  (~ Pd4) ) ;
 assign n122 = ( (~ Pf4)  &  n381 ) | ( Pf4  &  (~ n381) ) ;
 assign n123 = ( (~ Pz)  &  n380  &  n379 ) | ( (~ Pz)  &  n380  &  (~ n687) ) ;
 assign n124 = ( (~ Pz)  &  n374  &  n373 ) | ( (~ Pz)  &  n374  &  (~ n687) ) ;
 assign n125 = ( Pi4  &  n252 ) | ( (~ Pi4)  &  (~ n252) ) ;
 assign n126 = ( (~ Pz)  &  n361  &  n360 ) | ( (~ Pz)  &  n361  &  (~ n687) ) ;
 assign n127 = ( (~ Pz)  &  n355  &  n354 ) | ( (~ Pz)  &  n355  &  (~ n687) ) ;
 assign n128 = ( (~ Pz)  &  n341  &  n340 ) | ( (~ Pz)  &  n341  &  (~ n687) ) ;
 assign n129 = ( (~ Pz)  &  n320  &  n319 ) | ( (~ Pz)  &  n320  &  (~ n687) ) ;
 assign n130 = ( (~ Pz)  &  n307  &  n306 ) | ( (~ Pz)  &  n307  &  (~ n687) ) ;
 assign n131 = ( (~ Pz)  &  n293  &  n292 ) | ( (~ Pz)  &  n293  &  (~ n687) ) ;
 assign n132 = ( Pj4  &  Pz ) | ( Pj4  &  n687 ) ;
 assign n133 = ( (~ Pz)  &  n263  &  n262 ) | ( (~ Pz)  &  n263  &  (~ n687) ) ;
 assign n134 = ( Pr4  &  n187 ) | ( (~ Pr4)  &  (~ n187) ) ;
 assign n136 = ( Ps4  &  n514 ) | ( (~ Ps4)  &  (~ n514) ) ;
 assign n137 = ( Pt4  &  n641 ) | ( (~ Pt4)  &  (~ n641) ) ;
 assign n138 = ( Pu4  &  n656 ) | ( (~ Pu4)  &  (~ n656) ) ;
 assign n139 = ( Pv4  &  n627 ) | ( (~ Pv4)  &  (~ n627) ) ;
 assign n140 = ( Pw4  &  n628 ) | ( (~ Pw4)  &  (~ n628) ) ;
 assign n141 = ( Px4  &  n655 ) | ( (~ Px4)  &  (~ n655) ) ;
 assign n142 = ( Py4  &  n629 ) | ( (~ Py4)  &  (~ n629) ) ;
 assign n143 = ( Pz4  &  n336 ) | ( (~ Pz4)  &  (~ n336) ) ;
 assign n144 = ( (~ Pd5)  &  n506  &  n508 ) ;
 assign n147 = ( n182  &  n631 ) ;
 assign n145 = ( (~ Pg5)  &  (~ Pf5)  &  (~ n632) ) ;
 assign n146 = ( Pf5  &  n632 ) ;
 assign n150 = ( n147  &  Pz ) | ( n147  &  n378 ) ;
 assign n151 = ( (~ Pz)  &  (~ Pk5) ) | ( (~ Pz)  &  Pj5 ) ;
 assign n152 = ( (~ Pj5)  &  n186 ) | ( Pj5  &  (~ n186) ) ;
 assign n153 = ( (~ Pk5)  &  n359 ) | ( Pk5  &  (~ n359) ) ;
 assign n154 = ( n160  &  (~ n351)  &  n352 ) | ( n160  &  (~ n351)  &  (~ n506) ) ;
 assign n155 = ( n186  &  n339 ) | ( n186  &  (~ n506) ) ;
 assign n156 = ( Pm5  &  Pn5 ) ;
 assign n159 = ( (~ n186) ) | ( n318 ) | ( (~ n506) ) ;
 assign n160 = ( n182  &  (~ n186) ) | ( n182  &  (~ n339) ) ;
 assign n161 = ( (~ Pn5) ) | ( (~ Pm5) ) | ( (~ n503) ) ;
 assign n158 = ( n159  &  n160  &  n161  &  (~ n573) ) ;
 assign n163 = ( (~ Pr5)  &  n166  &  n291 ) | ( n166  &  n291  &  n290 ) ;
 assign n166 = ( n167  &  Pr5 ) | ( n167  &  Pp5 ) | ( n167  &  Pq5 ) ;
 assign n164 = ( n573 ) | ( Pb0 ) ;
 assign n167 = ( (~ Pz)  &  n249 ) | ( (~ Pz)  &  (~ Pq5)  &  (~ Pp5) ) ;
 assign n172 = ( Pm1 ) | ( Pn1 ) | ( n531 ) ;
 assign n169 = ( (~ Pv0)  &  n172 ) | ( n76  &  n172 ) | ( n172  &  (~ n544) ) ;
 assign n173 = ( Pv0  &  (~ Ph) ) | ( (~ Ph)  &  n76 ) | ( (~ Ph)  &  (~ n669) ) ;
 assign n176 = ( Pr4  &  (~ Pf0) ) | ( (~ Pf0)  &  n94 ) | ( (~ Pf0)  &  (~ n709) ) ;
 assign n182 = ( Pn5 ) | ( Pm5 ) | ( (~ n503) ) ;
 assign n179 = ( (~ Pr4)  &  n182 ) | ( n94  &  n182 ) | ( n182  &  (~ n206) ) ;
 assign n184 = ( (~ Pd5)  &  n510 ) ;
 assign n183 = ( (~ n94)  &  n184  &  (~ n205) ) ;
 assign n186 = ( (~ Pn5)  &  Pm5  &  n503 ) ;
 assign n185 = ( Pr5  &  n186  &  Pr4 ) ;
 assign n187 = ( (~ Pr5)  &  n184  &  (~ n205) ) | ( n184  &  (~ n186)  &  (~ n205) ) ;
 assign n191 = ( (~ Pq5) ) | ( Ph0 ) | ( (~ n186) ) ;
 assign n190 = ( n191  &  Pf3 ) | ( n191  &  Pg3 ) ;
 assign n195 = ( Pp5  &  (~ Ph0)  &  n186 ) ;
 assign n192 = ( (~ Pi3)  &  n195 ) | ( (~ Pi3)  &  (~ Ph3)  &  (~ n190) ) ;
 assign n198 = ( (~ Ph0)  &  (~ n192) ) ;
 assign n197 = ( Pp3  &  (~ Ph0) ) | ( (~ Pj3)  &  (~ Ph0) ) | ( (~ Ph0)  &  n198 ) ;
 assign n201 = ( (~ Pr5)  &  Pk5  &  (~ Pj5) ) | ( Pr4  &  Pk5  &  (~ Pj5) ) ;
 assign n206 = ( (~ Pz4)  &  (~ Ps4)  &  n517 ) ;
 assign n207 = ( (~ Pr4)  &  (~ n94) ) ;
 assign n205 = ( Pj10 ) | ( Pc5 ) ;
 assign n203 = ( (~ n184)  &  n206  &  n207 ) | ( n206  &  n207  &  n205 ) ;
 assign n208 = ( (~ Pg3)  &  n191 ) | ( (~ Pf3)  &  n191 ) ;
 assign n211 = ( Pi3  &  n195 ) | ( Pi3  &  Ph3  &  (~ n208) ) ;
 assign n214 = ( (~ Ph0)  &  (~ n211) ) ;
 assign n213 = ( (~ Pp3)  &  (~ Ph0) ) | ( (~ Pk3)  &  (~ Ph0) ) | ( (~ Ph0)  &  n214 ) ;
 assign n219 = ( n92 ) | ( n88 ) ;
 assign n217 = ( (~ Ps3)  &  n642 ) | ( Ps3  &  (~ n642) ) ;
 assign n221 = ( (~ Pq1) ) | ( Pj ) | ( n308 ) ;
 assign n220 = ( n221  &  Pq2 ) | ( n221  &  Pr2 ) ;
 assign n222 = ( (~ Pr2)  &  n221 ) | ( (~ Pq2)  &  n221 ) ;
 assign n227 = ( (~ Pf)  &  n308 ) | ( (~ Pv0)  &  Pr1  &  (~ Pf) ) ;
 assign n225 = ( Pv0  &  n227 ) | ( n76  &  n227 ) | ( n227  &  (~ n666) ) ;
 assign n229 = ( n74 ) | ( n225 ) ;
 assign n230 = ( (~ n74) ) | ( n225 ) ;
 assign n228 = ( n222  &  n220 ) | ( n229  &  n220 ) | ( n222  &  n230 ) | ( n229  &  n230 ) ;
 assign n233 = ( (~ Py0)  &  (~ Px0) ) ;
 assign n231 = ( Pp1  &  n233 ) | ( (~ Pz0)  &  Pq1  &  n233 ) ;
 assign n235 = ( (~ Pu3)  &  n671 ) | ( (~ Pp0)  &  n671 ) ;
 assign n236 = ( (~ Ps0)  &  n670 ) | ( (~ Pe4)  &  n670 ) ;
 assign n237 = ( (~ Pm0)  &  n672  &  n673 ) | ( (~ Pg3)  &  n672  &  n673 ) ;
 assign n234 = ( n235  &  n236  &  n237 ) ;
 assign n239 = ( Pq3 ) | ( n197 ) | ( n266 ) ;
 assign n240 = ( (~ Pq3) ) | ( n213 ) | ( n265 ) ;
 assign n238 = ( n239  &  n240 ) ;
 assign n241 = ( (~ Pr1)  &  (~ Pq1) ) | ( (~ Pr1)  &  (~ Pp1) ) ;
 assign n246 = ( (~ Pv3)  &  n676 ) | ( (~ Pp0)  &  n676 ) ;
 assign n247 = ( (~ Ps0)  &  n675 ) | ( (~ Pf4)  &  n675 ) ;
 assign n248 = ( (~ Pm0)  &  n677  &  n678 ) | ( (~ Ph3)  &  n677  &  n678 ) ;
 assign n245 = ( n246  &  n247  &  n248 ) ;
 assign n249 = ( (~ Pr5)  &  (~ Pq5) ) | ( (~ Pr5)  &  (~ Pp5) ) ;
 assign n253 = ( (~ Pf4) ) | ( (~ Pe4) ) | ( (~ Pd4) ) ;
 assign n252 = ( (~ Pq5)  &  n253 ) | ( Pj0  &  n253 ) ;
 assign n254 = ( (~ Pp5)  &  (~ Pj0)  &  (~ Pi4) ) | ( (~ Pp5)  &  (~ Pj0)  &  n252 ) ;
 assign n260 = ( (~ Pj4) ) | ( (~ Ph4) ) | ( n578 ) ;
 assign n257 = ( (~ Pl4)  &  (~ Pj0) ) | ( (~ Pk4)  &  (~ Pj0) ) | ( (~ Pj0)  &  n260 ) ;
 assign n263 = ( (~ Pc4) ) | ( n687 ) ;
 assign n262 = ( (~ Pq4)  &  n716 ) | ( Pq4  &  (~ n716) ) ;
 assign n265 = ( n92 ) | ( (~ n369) ) ;
 assign n266 = ( (~ n92) ) | ( (~ n369) ) ;
 assign n264 = ( n213  &  n197 ) | ( n265  &  n197 ) | ( n213  &  n266 ) | ( n265  &  n266 ) ;
 assign n267 = ( (~ Pq3)  &  n264 ) | ( Pq3  &  (~ n264) ) ;
 assign n269 = ( (~ Pw3)  &  n683 ) | ( (~ Pp0)  &  n683 ) ;
 assign n270 = ( (~ Ps0)  &  n682 ) | ( (~ Pi4)  &  n682 ) ;
 assign n271 = ( (~ Pm0)  &  n684  &  n685 ) | ( (~ Pi3)  &  n684  &  n685 ) ;
 assign n268 = ( n269  &  n270  &  n271 ) ;
 assign n273 = ( n214 ) | ( n265 ) ;
 assign n274 = ( n198 ) | ( n266 ) ;
 assign n272 = ( (~ Pk3)  &  (~ Pj3) ) | ( (~ Pj3)  &  n273 ) | ( (~ Pk3)  &  n274 ) | ( n273  &  n274 ) ;
 assign n275 = ( (~ Pp3)  &  n272 ) | ( Pp3  &  (~ n272) ) ;
 assign n277 = ( (~ Pd2) ) | ( (~ Pc2) ) | ( (~ Pb2) ) ;
 assign n276 = ( (~ Pq1)  &  n277 ) | ( Pl  &  n277 ) ;
 assign n278 = ( (~ Pp1)  &  (~ Pl)  &  (~ Pg2) ) | ( (~ Pp1)  &  (~ Pl)  &  n276 ) ;
 assign n282 = ( (~ Pq1)  &  (~ Pp1) ) | ( (~ Pp1)  &  (~ n36) ) | ( (~ Pq1)  &  n568 ) | ( (~ n36)  &  n568 ) ;
 assign n284 = ( (~ Pt)  &  (~ Ps) ) | ( (~ Ps)  &  (~ Pe2) ) | ( (~ Pt)  &  n500 ) | ( (~ Pe2)  &  n500 ) ;
 assign n285 = ( (~ Pr) ) | ( (~ Pn1) ) ;
 assign n286 = ( (~ Pz0)  &  (~ Pw) ) | ( (~ Pw)  &  (~ Pv) ) | ( (~ Pz0)  &  (~ Pl1) ) | ( (~ Pv)  &  (~ Pl1) ) ;
 assign n287 = ( (~ Pu) ) | ( (~ n225) ) ;
 assign n288 = ( (~ Pw2)  &  (~ Pm) ) | ( (~ Pn)  &  (~ Pm) ) | ( (~ Pw2)  &  (~ n329) ) | ( (~ Pn)  &  (~ n329) ) ;
 assign n289 = ( (~ Po)  &  n689 ) | ( n311  &  n689 ) ;
 assign n283 = ( n284  &  n285  &  n286  &  n287  &  n288  &  n289 ) ;
 assign n291 = ( (~ Pq5)  &  (~ Pp5) ) | ( (~ Pp5)  &  (~ n164) ) | ( (~ Pq5)  &  (~ n575) ) | ( (~ n164)  &  (~ n575) ) ;
 assign n290 = ( (~ Pc0)  &  n161 ) ;
 assign n293 = ( (~ Pb4) ) | ( n687 ) ;
 assign n292 = ( (~ Po4)  &  n581 ) | ( Po4  &  (~ n581) ) ;
 assign n294 = ( (~ Po3)  &  n643 ) | ( Po3  &  (~ n643) ) ;
 assign n298 = ( (~ Ph2) ) | ( (~ Pf2) ) | ( n588 ) ;
 assign n295 = ( (~ Pl)  &  (~ Pj2) ) | ( (~ Pl)  &  (~ Pi2) ) | ( (~ Pl)  &  n298 ) ;
 assign n301 = ( (~ Pa2) ) | ( (~ n299) ) ;
 assign n299 = ( (~ n365) ) | ( (~ n500) ) ;
 assign n300 = ( (~ Po2)  &  n722 ) | ( Po2  &  (~ n722) ) ;
 assign n303 = ( (~ Pr)  &  n691 ) | ( (~ Pm1)  &  n691 ) ;
 assign n304 = ( (~ Pu)  &  n690 ) | ( (~ Pb2)  &  n690 ) ;
 assign n305 = ( (~ Pq2)  &  n692  &  n693 ) | ( (~ Po)  &  n692  &  n693 ) ;
 assign n302 = ( n303  &  n304  &  n305 ) ;
 assign n307 = ( (~ Pa4) ) | ( n687 ) ;
 assign n306 = ( (~ Pn4)  &  n723 ) | ( Pn4  &  (~ n723) ) ;
 assign n308 = ( Pn1 ) | ( (~ Pm1) ) | ( n531 ) ;
 assign n310 = ( Pf1 ) | ( (~ Pe1) ) ;
 assign n311 = ( (~ Pe3) ) | ( (~ Pd3) ) | ( (~ Pc3) ) ;
 assign n313 = ( (~ Ps1)  &  n696 ) | ( (~ Pr)  &  n696 ) ;
 assign n314 = ( (~ Pu)  &  n695 ) | ( (~ Pc2)  &  n695 ) ;
 assign n315 = ( (~ Pr2)  &  n697  &  n698 ) | ( (~ Po)  &  n697  &  n698 ) ;
 assign n312 = ( n313  &  n314  &  n315 ) ;
 assign n318 = ( (~ Pt3) ) | ( (~ Ps3) ) | ( (~ Pr3) ) | ( (~ Pq3) ) | ( (~ Pp3) ) ;
 assign n320 = ( (~ Pz3) ) | ( n687 ) ;
 assign n319 = ( (~ Pm4)  &  n257 ) | ( Pm4  &  (~ n257) ) ;
 assign n322 = ( (~ Pz1) ) | ( (~ n299) ) ;
 assign n321 = ( (~ Pm2)  &  n617 ) | ( Pm2  &  (~ n617) ) ;
 assign n324 = ( (~ Ph1)  &  n541 ) ;
 assign n323 = ( (~ Pr1)  &  n324  &  (~ n543) ) | ( n308  &  n324  &  (~ n543) ) ;
 assign n326 = ( (~ Pc1) ) | ( n626 ) ;
 assign n325 = ( (~ Pd1)  &  (~ Pc) ) | ( Pr1  &  (~ Pc)  &  n326 ) ;
 assign n329 = ( (~ Pz2)  &  Py2  &  (~ Pe3)  &  (~ Pd3)  &  (~ Pc3)  &  (~ Pb3)  &  (~ Pa3) ) ;
 assign n332 = ( (~ Pt1)  &  n701 ) | ( (~ Pr)  &  n701 ) ;
 assign n333 = ( (~ Pu)  &  n700 ) | ( (~ Pd2)  &  n700 ) ;
 assign n334 = ( (~ Ps2)  &  n702  &  n703 ) | ( (~ Po)  &  n702  &  n703 ) ;
 assign n331 = ( n332  &  n333  &  n334 ) ;
 assign n336 = ( (~ Py4) ) | ( n629 ) ;
 assign n335 = ( (~ Pz4)  &  (~ Pa0) ) | ( Pr5  &  (~ Pa0)  &  n336 ) ;
 assign n339 = ( (~ Pt3)  &  (~ Ps3)  &  (~ Pr3)  &  (~ Pq3)  &  (~ Pp3)  &  (~ Po3)  &  Pn3 ) ;
 assign n341 = ( (~ Py3) ) | ( n687 ) ;
 assign n340 = ( (~ Pl4)  &  n725 ) | ( Pl4  &  (~ n725) ) ;
 assign n343 = ( (~ Py1) ) | ( (~ n299) ) ;
 assign n342 = ( (~ Pl2)  &  n726 ) | ( Pl2  &  (~ n726) ) ;
 assign n344 = ( (~ n308)  &  n310 ) | ( (~ n308)  &  n311 ) ;
 assign n345 = ( Pn1 ) | ( (~ Pm1) ) | ( Pl1 ) | ( Pb ) ;
 assign n348 = ( (~ Pu1)  &  n706 ) | ( (~ Pr)  &  n706 ) ;
 assign n349 = ( (~ Pu)  &  n705 ) | ( (~ Pg2)  &  n705 ) ;
 assign n350 = ( (~ Pt2)  &  n707  &  n708 ) | ( (~ Po)  &  n707  &  n708 ) ;
 assign n347 = ( n348  &  n349  &  n350 ) ;
 assign n351 = ( n186  &  n318 ) | ( n186  &  (~ n506) ) ;
 assign n352 = ( Pz ) | ( Pn5 ) | ( (~ Pm5) ) | ( Pl5 ) ;
 assign n355 = ( (~ Px3) ) | ( n687 ) ;
 assign n354 = ( (~ Pk4)  &  n260 ) | ( Pk4  &  (~ n260) ) ;
 assign n357 = ( (~ Px1) ) | ( (~ n299) ) ;
 assign n356 = ( (~ Pk2)  &  n295 ) | ( Pk2  &  (~ n295) ) ;
 assign n359 = ( Pj5  &  n186 ) ;
 assign n361 = ( (~ Pw3) ) | ( n687 ) ;
 assign n360 = ( (~ Pj4)  &  n727 ) | ( Pj4  &  (~ n727) ) ;
 assign n363 = ( (~ Pw1) ) | ( (~ n299) ) ;
 assign n362 = ( (~ Pj2)  &  n729 ) | ( Pj2  &  (~ n729) ) ;
 assign n365 = ( (~ Pn1) ) | ( Pm1 ) | ( n531 ) ;
 assign n364 = ( (~ Pj1)  &  n500 ) | ( Pj1  &  (~ n500) ) ;
 assign n369 = ( Pd0 ) | ( n201 ) | ( n203 ) ;
 assign n367 = ( (~ Ph3)  &  n92  &  (~ n190) ) ;
 assign n368 = ( Ph3  &  (~ n92)  &  (~ n208) ) ;
 assign n366 = ( n369  &  n367 ) | ( n369  &  n368 ) | ( n369  &  n195 ) ;
 assign n370 = ( Pi3  &  n366 ) | ( (~ Pi3)  &  (~ n366) ) ;
 assign n372 = ( (~ Pv1) ) | ( (~ n299) ) ;
 assign n371 = ( (~ Pi2)  &  n298 ) | ( Pi2  &  (~ n298) ) ;
 assign n374 = ( (~ Pv3) ) | ( n687 ) ;
 assign n373 = ( (~ Ph4)  &  n578 ) | ( Ph4  &  (~ n578) ) ;
 assign n375 = ( n208  &  n190 ) | ( n265  &  n190 ) | ( n208  &  n266 ) | ( n265  &  n266 ) ;
 assign n377 = ( (~ Pu1) ) | ( (~ n299) ) ;
 assign n376 = ( (~ Ph2)  &  n733 ) | ( Ph2  &  (~ n733) ) ;
 assign n378 = ( (~ Ph5)  &  n501 ) | ( Ph5  &  (~ n501) ) ;
 assign n380 = ( (~ Pu3) ) | ( n687 ) ;
 assign n379 = ( (~ Pg4)  &  n254 ) | ( Pg4  &  (~ n254) ) ;
 assign n381 = ( Pd4  &  Pe4 ) ;
 assign n383 = ( (~ Pt1) ) | ( (~ n299) ) ;
 assign n382 = ( (~ Pf2)  &  n588 ) | ( Pf2  &  (~ n588) ) ;
 assign n387 = ( Pp1  &  (~ Pj)  &  (~ n308) ) ;
 assign n384 = ( (~ Pt2)  &  n387 ) | ( (~ Pt2)  &  (~ Ps2)  &  (~ n220) ) ;
 assign n390 = ( (~ Pj)  &  (~ n384) ) ;
 assign n389 = ( (~ Pu2)  &  (~ Pj) ) | ( (~ Pj)  &  Pa3 ) | ( (~ Pj)  &  n390 ) ;
 assign n393 = ( Pt2  &  n387 ) | ( Pt2  &  Ps2  &  (~ n222) ) ;
 assign n396 = ( (~ Pj)  &  (~ n393) ) ;
 assign n395 = ( (~ Pv2)  &  (~ Pj) ) | ( (~ Pj)  &  (~ Pa3) ) | ( (~ Pj)  &  n396 ) ;
 assign n401 = ( n74 ) | ( n70 ) ;
 assign n399 = ( (~ Pe3)  &  n644 ) | ( Pe3  &  (~ n644) ) ;
 assign n403 = ( (~ Ps1) ) | ( (~ n299) ) ;
 assign n402 = ( (~ Pe2)  &  n278 ) | ( Pe2  &  (~ n278) ) ;
 assign n404 = ( (~ Pd3)  &  n645 ) | ( Pd3  &  (~ n645) ) ;
 assign n405 = ( Pc2  &  Pb2 ) ;
 assign n406 = ( (~ n76)  &  n324  &  (~ n543) ) ;
 assign n407 = ( Pv0  &  Pr1  &  (~ n308) ) ;
 assign n410 = ( (~ Pu4)  &  (~ Pt4) ) ;
 assign n408 = ( Pp5  &  n410 ) | ( (~ Pv4)  &  Pq5  &  n410 ) ;
 assign n411 = ( Pw3  &  (~ Pi0) ) | ( Pv3  &  (~ Pi0) ) | ( Pu3  &  (~ Pi0) ) ;
 assign n414 = ( Px3 ) | ( n411 ) ;
 assign n413 = ( Pz3  &  (~ Pi0) ) | ( Py3  &  (~ Pi0) ) | ( (~ Pi0)  &  n414 ) ;
 assign n415 = ( (~ Pw3)  &  (~ Pi0) ) | ( (~ Pv3)  &  (~ Pi0) ) | ( (~ Pu3)  &  (~ Pi0) ) ;
 assign n422 = ( (~ Px3) ) | ( n415 ) ;
 assign n419 = ( (~ Pz3)  &  (~ Pi0) ) | ( (~ Py3)  &  (~ Pi0) ) | ( (~ Pi0)  &  n422 ) ;
 assign n424 = ( (~ Pt3) ) | ( n179 ) ;
 assign n423 = ( (~ Pc4)  &  n646 ) | ( Pc4  &  (~ n646) ) ;
 assign n426 = ( Pb3 ) | ( n389 ) | ( n230 ) ;
 assign n427 = ( (~ Pb3) ) | ( n229 ) | ( n395 ) ;
 assign n425 = ( n426  &  n427 ) ;
 assign n429 = ( (~ Ps3) ) | ( n179 ) ;
 assign n428 = ( (~ Pb4)  &  n647 ) | ( Pb4  &  (~ n647) ) ;
 assign n430 = ( n395  &  n389 ) | ( n229  &  n389 ) | ( n395  &  n230 ) | ( n229  &  n230 ) ;
 assign n431 = ( (~ Pb3)  &  n430 ) | ( Pb3  &  (~ n430) ) ;
 assign n433 = ( n413 ) | ( n460 ) ;
 assign n434 = ( n419 ) | ( n459 ) ;
 assign n432 = ( n433  &  n434 ) ;
 assign n436 = ( n396 ) | ( n229 ) ;
 assign n437 = ( n390 ) | ( n230 ) ;
 assign n435 = ( (~ Pv2)  &  (~ Pu2) ) | ( (~ Pu2)  &  n436 ) | ( (~ Pv2)  &  n437 ) | ( n436  &  n437 ) ;
 assign n438 = ( (~ Pa3)  &  n435 ) | ( Pa3  &  (~ n435) ) ;
 assign n439 = ( Pu1  &  (~ Pk) ) | ( Pt1  &  (~ Pk) ) | ( Ps1  &  (~ Pk) ) ;
 assign n442 = ( Pv1 ) | ( n439 ) ;
 assign n441 = ( Px1  &  (~ Pk) ) | ( Pw1  &  (~ Pk) ) | ( (~ Pk)  &  n442 ) ;
 assign n443 = ( (~ Pu1)  &  (~ Pk) ) | ( (~ Pt1)  &  (~ Pk) ) | ( (~ Ps1)  &  (~ Pk) ) ;
 assign n450 = ( (~ Pv1) ) | ( n443 ) ;
 assign n447 = ( (~ Px1)  &  (~ Pk) ) | ( (~ Pw1)  &  (~ Pk) ) | ( (~ Pk)  &  n450 ) ;
 assign n452 = ( (~ Pe3) ) | ( n169 ) ;
 assign n451 = ( (~ Pa2)  &  n649 ) | ( Pa2  &  (~ n649) ) ;
 assign n454 = ( (~ Pq3) ) | ( n179 ) ;
 assign n453 = ( (~ Pz3)  &  n650 ) | ( Pz3  &  (~ n650) ) ;
 assign n455 = ( (~ Pz2)  &  n651 ) | ( Pz2  &  (~ n651) ) ;
 assign n457 = ( (~ Pd3) ) | ( n169 ) ;
 assign n456 = ( (~ Pz1)  &  n652 ) | ( Pz1  &  (~ n652) ) ;
 assign n459 = ( n176 ) | ( (~ n636) ) ;
 assign n460 = ( n176 ) | ( n636 ) ;
 assign n458 = ( n422  &  n414 ) | ( n459  &  n414 ) | ( n422  &  n460 ) | ( n459  &  n460 ) ;
 assign n462 = ( (~ Pp3) ) | ( n179 ) ;
 assign n461 = ( (~ Py3)  &  n458 ) | ( Py3  &  (~ n458) ) ;
 assign n464 = ( n441 ) | ( n477 ) ;
 assign n465 = ( n447 ) | ( n476 ) ;
 assign n463 = ( n464  &  n465 ) ;
 assign n466 = ( n415  &  n411 ) | ( n459  &  n411 ) | ( n415  &  n460 ) | ( n459  &  n460 ) ;
 assign n468 = ( (~ Po3) ) | ( n179 ) ;
 assign n467 = ( (~ Px3)  &  n466 ) | ( Px3  &  (~ n466) ) ;
 assign n470 = ( Pw2 ) | ( n437 ) ;
 assign n471 = ( (~ Pw2) ) | ( n436 ) ;
 assign n469 = ( n470  &  n471 ) ;
 assign n473 = ( (~ Pb3) ) | ( n169 ) ;
 assign n472 = ( (~ Px1)  &  n654 ) | ( Px1  &  (~ n654) ) ;
 assign n474 = ( n437  &  n436 ) ;
 assign n476 = ( n173 ) | ( (~ n638) ) ;
 assign n477 = ( n173 ) | ( n638 ) ;
 assign n475 = ( n450  &  n442 ) | ( n476  &  n442 ) | ( n450  &  n477 ) | ( n476  &  n477 ) ;
 assign n479 = ( (~ Pa3) ) | ( n169 ) ;
 assign n478 = ( (~ Pw1)  &  n475 ) | ( Pw1  &  (~ n475) ) ;
 assign n480 = ( n443  &  n439 ) | ( n476  &  n439 ) | ( n443  &  n477 ) | ( n476  &  n477 ) ;
 assign n482 = ( (~ Pz2) ) | ( n169 ) ;
 assign n481 = ( (~ Pv1)  &  n480 ) | ( Pv1  &  (~ n480) ) ;
 assign n484 = ( (~ Pr0)  &  (~ Pq0) ) | ( (~ Pq0)  &  (~ Pg4) ) | ( (~ Pr0)  &  n501 ) | ( (~ Pg4)  &  n501 ) ;
 assign n485 = ( (~ Pp0) ) | ( (~ Pn5) ) ;
 assign n486 = ( (~ Pv4)  &  (~ Pu0) ) | ( (~ Pu0)  &  (~ Pt0) ) | ( (~ Pv4)  &  (~ Pl5) ) | ( (~ Pt0)  &  (~ Pl5) ) ;
 assign n487 = ( (~ Ps0) ) | ( n369 ) ;
 assign n488 = ( (~ Pl3)  &  (~ Pk0) ) | ( (~ Pl0)  &  (~ Pk0) ) | ( (~ Pl3)  &  (~ n339) ) | ( (~ Pl0)  &  (~ n339) ) ;
 assign n489 = ( (~ Pm0)  &  n710 ) | ( n318  &  n710 ) ;
 assign n483 = ( n484  &  n485  &  n486  &  n487  &  n488  &  n489 ) ;
 assign n490 = ( (~ Pt3)  &  n657 ) | ( Pt3  &  (~ n657) ) ;
 assign n492 = ( (~ Ps2)  &  n74  &  (~ n220) ) ;
 assign n493 = ( Ps2  &  (~ n74)  &  (~ n222) ) ;
 assign n491 = ( (~ n225)  &  n387 ) | ( (~ n225)  &  n492 ) | ( (~ n225)  &  n493 ) ;
 assign n495 = ( Pt2  &  n491 ) | ( (~ Pt2)  &  (~ n491) ) ;
 assign n497 = ( (~ Pp0)  &  n712 ) | ( (~ Pm5)  &  n712 ) ;
 assign n498 = ( (~ Ps0)  &  n711 ) | ( (~ Pd4)  &  n711 ) ;
 assign n499 = ( (~ Pm0)  &  n713  &  n714 ) | ( (~ Pf3)  &  n713  &  n714 ) ;
 assign n496 = ( n497  &  n498  &  n499 ) ;
 assign n500 = ( (~ Pn2) ) | ( n588 ) ;
 assign n501 = ( (~ Pp4) ) | ( n578 ) ;
 assign n503 = ( (~ Pz)  &  Pl5 ) ;
 assign n506 = ( (~ Pb5)  &  Pa5 ) ;
 assign n508 = ( (~ Po5) ) | ( Pi5 ) | ( (~ Pg5) ) ;
 assign n510 = ( Pe5 ) | ( n506 ) | ( n508 ) ;
 assign n514 = ( (~ Pr4) ) | ( n187 ) ;
 assign n515 = ( Pz ) | ( n183 ) | ( n185 ) | ( (~ n631) ) ;
 assign n517 = ( (~ Py4)  &  (~ Px4)  &  (~ Pw4)  &  (~ Pv4)  &  (~ Pu4)  &  (~ Pt4) ) ;
 assign n531 = ( (~ Pl1) ) | ( Pb ) ;
 assign n532 = ( (~ Pz0)  &  (~ Py0)  &  (~ Px0)  &  (~ Pc1)  &  (~ Pb1)  &  (~ Pa1) ) ;
 assign n538 = ( (~ Po1) ) | ( Pk1 ) | ( (~ Pj1) ) ;
 assign n541 = ( Pi1 ) | ( (~ n310) ) | ( n538 ) ;
 assign n543 = ( Pn6 ) | ( Pg1 ) ;
 assign n544 = ( (~ Pw0)  &  (~ Pd1)  &  n532 ) ;
 assign n566 = ( Pe ) | ( (~ n33) ) ;
 assign n568 = ( n36 ) | ( n566 ) ;
 assign n573 = ( (~ Pz)  &  Pn5  &  (~ Pm5)  &  (~ Pl5) ) ;
 assign n575 = ( (~ n164)  &  n290 ) ;
 assign n578 = ( (~ Pg4) ) | ( n254 ) ;
 assign n581 = ( (~ Pn4) ) | ( (~ Pm4) ) | ( n257 ) ;
 assign n588 = ( (~ Pe2) ) | ( n278 ) ;
 assign n609 = ( (~ Pl3) ) | ( n273 ) ;
 assign n611 = ( Pl3 ) | ( n274 ) ;
 assign n617 = ( (~ Pl2) ) | ( (~ Pk2) ) | ( n295 ) ;
 assign n624 = ( (~ Py0) ) | ( (~ Px0) ) | ( (~ Pw0) ) | ( (~ Pv0) ) | ( n323 ) ;
 assign n625 = ( (~ Pz0) ) | ( n624 ) ;
 assign n626 = ( (~ Pb1) ) | ( (~ Pa1) ) | ( n625 ) ;
 assign n627 = ( (~ Pu4) ) | ( (~ Pt4) ) | ( (~ Ps4) ) | ( (~ Pr4) ) | ( n187 ) ;
 assign n628 = ( (~ Pv4) ) | ( n627 ) ;
 assign n629 = ( (~ Px4) ) | ( (~ Pw4) ) | ( n628 ) ;
 assign n631 = ( (~ Pn5) ) | ( Pm5 ) | ( (~ n503) ) ;
 assign n632 = ( Ph5 ) | ( n150 ) ;
 assign n633 = ( Pb ) | ( (~ n365) ) | ( n406 ) | ( n407 ) ;
 assign n636 = ( Pg0 ) | ( n205 ) ;
 assign n638 = ( Pi ) | ( n543 ) ;
 assign n639 = ( (~ Pv0) ) | ( n323 ) ;
 assign n640 = ( (~ Pw0) ) | ( n639 ) ;
 assign n641 = ( (~ Ps4) ) | ( n514 ) ;
 assign n642 = ( (~ Pr3)  &  n239 ) | ( Pr3  &  n240 ) | ( n239  &  n240 ) ;
 assign n643 = ( (~ Pn3)  &  n720 ) | ( (~ Pm3)  &  n720 ) | ( n609  &  n720 ) ;
 assign n644 = ( (~ Pd3)  &  n738 ) | ( (~ Pc3)  &  n738 ) | ( n427  &  n738 ) ;
 assign n645 = ( (~ Pc3)  &  n426 ) | ( Pc3  &  n427 ) | ( n426  &  n427 ) ;
 assign n646 = ( (~ Pb4)  &  n742 ) | ( (~ Pa4)  &  n742 ) | ( n434  &  n742 ) ;
 assign n647 = ( (~ Pa4)  &  n433 ) | ( Pa4  &  n434 ) | ( n433  &  n434 ) ;
 assign n648 = ( (~ Pa1) ) | ( n625 ) ;
 assign n649 = ( (~ Pz1)  &  n743 ) | ( (~ Py1)  &  n743 ) | ( n465  &  n743 ) ;
 assign n650 = ( (~ Py3)  &  n744 ) | ( n422  &  n744 ) | ( n459  &  n744 ) ;
 assign n651 = ( (~ Py2)  &  n745 ) | ( (~ Px2)  &  n745 ) | ( n471  &  n745 ) ;
 assign n652 = ( (~ Py1)  &  n464 ) | ( Py1  &  n465 ) | ( n464  &  n465 ) ;
 assign n653 = ( (~ Px0) ) | ( n640 ) ;
 assign n654 = ( (~ Pw1)  &  n747 ) | ( n450  &  n747 ) | ( n476  &  n747 ) ;
 assign n655 = ( (~ Pw4) ) | ( n628 ) ;
 assign n656 = ( (~ Pt4) ) | ( n641 ) ;
 assign n657 = ( (~ Ps3)  &  n754 ) | ( (~ Pr3)  &  n754 ) | ( n240  &  n754 ) ;
 assign n658 = ( (~ Pp2)  &  Pa ) | ( (~ Pp2)  &  n717 ) | ( Pa  &  (~ n717) ) ;
 assign n659 = ( (~ n88)  &  (~ n92) ) | ( n88  &  n728 ) | ( (~ n92)  &  n728 ) ;
 assign n660 = ( Pi1  &  (~ n763) ) | ( (~ n23)  &  (~ n763) ) ;
 assign n661 = ( n734  &  Ph1 ) | ( n734  &  n541 ) ;
 assign n662 = ( (~ Pg5)  &  (~ Pf5) ) | ( (~ Pg5)  &  n632 ) | ( (~ Pf5)  &  (~ n632) ) ;
 assign n663 = ( Pe5  &  (~ n764) ) | ( (~ n144)  &  (~ n764) ) ;
 assign n664 = ( n741  &  Pd5 ) | ( n741  &  n510 ) ;
 assign n665 = ( (~ n70)  &  (~ n74) ) | ( n70  &  n751 ) | ( (~ n74)  &  n751 ) ;
 assign n666 = ( (~ n324)  &  n544 ) | ( n543  &  n544 ) ;
 assign n669 = ( Pw0  &  n231 ) | ( Pw0  &  n532  &  Pr1 ) ;
 assign n670 = ( (~ Px4)  &  (~ Pu0) ) | ( (~ Pu0)  &  (~ Pt0) ) | ( (~ Px4)  &  (~ Ps4) ) | ( (~ Pt0)  &  (~ Ps4) ) ;
 assign n671 = ( (~ Pr0)  &  (~ Pq0) ) | ( (~ Pr0)  &  (~ Pn4) ) | ( (~ Pq0)  &  (~ Pj4) ) | ( (~ Pn4)  &  (~ Pj4) ) ;
 assign n672 = ( (~ Px3)  &  (~ Pn0) ) | ( (~ Po0)  &  (~ Pn0) ) | ( (~ Px3)  &  (~ Pa4) ) | ( (~ Po0)  &  (~ Pa4) ) ;
 assign n673 = ( (~ Pr3)  &  (~ Pn3) ) | ( (~ Pr3)  &  (~ Pl0) ) | ( (~ Pn3)  &  (~ Pk0) ) | ( (~ Pl0)  &  (~ Pk0) ) ;
 assign n674 = ( (~ Pr1)  &  (~ Pq1) ) | ( (~ Pr1)  &  (~ n566) ) | ( (~ Pq1)  &  n568 ) | ( (~ n566)  &  n568 ) ;
 assign n675 = ( (~ Py4)  &  (~ Pu0) ) | ( (~ Py4)  &  (~ Pt4) ) | ( (~ Pu0)  &  (~ Pt0) ) | ( (~ Pt4)  &  (~ Pt0) ) ;
 assign n676 = ( (~ Pr0)  &  (~ Pq0) ) | ( (~ Pr0)  &  (~ Po4) ) | ( (~ Pq0)  &  (~ Pk4) ) | ( (~ Po4)  &  (~ Pk4) ) ;
 assign n677 = ( (~ Py3)  &  (~ Pn0) ) | ( (~ Po0)  &  (~ Pn0) ) | ( (~ Py3)  &  (~ Pb4) ) | ( (~ Po0)  &  (~ Pb4) ) ;
 assign n678 = ( (~ Ps3)  &  (~ Po3) ) | ( (~ Ps3)  &  (~ Pl0) ) | ( (~ Po3)  &  (~ Pk0) ) | ( (~ Pl0)  &  (~ Pk0) ) ;
 assign n679 = ( (~ Pr5)  &  (~ Pq5) ) | ( (~ Pr5)  &  n290 ) | ( (~ Pq5)  &  (~ n575) ) | ( n290  &  (~ n575) ) ;
 assign n681 = ( (~ Pq1)  &  (~ Pp1) ) | ( (~ Pq1)  &  (~ n566) ) | ( (~ Pp1)  &  n568 ) | ( (~ n566)  &  n568 ) ;
 assign n682 = ( (~ Pz4)  &  (~ Pu4) ) | ( (~ Pz4)  &  (~ Pu0) ) | ( (~ Pu4)  &  (~ Pt0) ) | ( (~ Pu0)  &  (~ Pt0) ) ;
 assign n683 = ( (~ Pr0)  &  (~ Pq4) ) | ( (~ Pr0)  &  (~ Pq0) ) | ( (~ Pq4)  &  (~ Pl4) ) | ( (~ Pq0)  &  (~ Pl4) ) ;
 assign n684 = ( (~ Pz3)  &  (~ Pn0) ) | ( (~ Po0)  &  (~ Pn0) ) | ( (~ Pz3)  &  (~ Pc4) ) | ( (~ Po0)  &  (~ Pc4) ) ;
 assign n685 = ( (~ Pt3)  &  (~ Pp3) ) | ( (~ Pt3)  &  (~ Pl0) ) | ( (~ Pp3)  &  (~ Pk0) ) | ( (~ Pl0)  &  (~ Pk0) ) ;
 assign n686 = ( (~ Pq5)  &  (~ Pp5) ) | ( (~ Pq5)  &  n290 ) | ( (~ Pp5)  &  (~ n575) ) | ( n290  &  (~ n575) ) ;
 assign n687 = ( n631  &  n501 ) ;
 assign n689 = ( (~ Pq1)  &  (~ Pq) ) | ( (~ Pq)  &  (~ Pp) ) | ( (~ Pq1)  &  n70 ) | ( (~ Pp)  &  n70 ) ;
 assign n690 = ( (~ Pw)  &  (~ Pv) ) | ( (~ Pv0)  &  (~ Pv) ) | ( (~ Pw)  &  (~ Pa1) ) | ( (~ Pv0)  &  (~ Pa1) ) ;
 assign n691 = ( (~ Pt)  &  (~ Ps) ) | ( (~ Pt)  &  (~ Pk2) ) | ( (~ Ps)  &  (~ Pf2) ) | ( (~ Pk2)  &  (~ Pf2) ) ;
 assign n692 = ( (~ Pr1)  &  (~ Pp1) ) | ( (~ Pq)  &  (~ Pp1) ) | ( (~ Pr1)  &  (~ Pp) ) | ( (~ Pq)  &  (~ Pp) ) ;
 assign n693 = ( (~ Px2)  &  (~ Pm) ) | ( (~ Pn)  &  (~ Pm) ) | ( (~ Px2)  &  (~ Pb3) ) | ( (~ Pn)  &  (~ Pb3) ) ;
 assign n695 = ( (~ Pw0)  &  (~ Pv) ) | ( (~ Pw)  &  (~ Pv) ) | ( (~ Pw0)  &  (~ Pb1) ) | ( (~ Pw)  &  (~ Pb1) ) ;
 assign n696 = ( (~ Pt)  &  (~ Ps) ) | ( (~ Pt)  &  (~ Pl2) ) | ( (~ Ps)  &  (~ Ph2) ) | ( (~ Pl2)  &  (~ Ph2) ) ;
 assign n697 = ( (~ Py1)  &  (~ Pv1) ) | ( (~ Py1)  &  (~ Pq) ) | ( (~ Pv1)  &  (~ Pp) ) | ( (~ Pq)  &  (~ Pp) ) ;
 assign n698 = ( (~ Py2)  &  (~ Pm) ) | ( (~ Pn)  &  (~ Pm) ) | ( (~ Py2)  &  (~ Pc3) ) | ( (~ Pn)  &  (~ Pc3) ) ;
 assign n699 = ( n34  &  n345  &  n76 ) | ( n34  &  n345  &  n325 ) ;
 assign n700 = ( (~ Px0)  &  (~ Pv) ) | ( (~ Pw)  &  (~ Pv) ) | ( (~ Px0)  &  (~ Pc1) ) | ( (~ Pw)  &  (~ Pc1) ) ;
 assign n701 = ( (~ Pt)  &  (~ Ps) ) | ( (~ Pt)  &  (~ Pm2) ) | ( (~ Ps)  &  (~ Pi2) ) | ( (~ Pm2)  &  (~ Pi2) ) ;
 assign n702 = ( (~ Pz1)  &  (~ Pw1) ) | ( (~ Pz1)  &  (~ Pq) ) | ( (~ Pw1)  &  (~ Pp) ) | ( (~ Pq)  &  (~ Pp) ) ;
 assign n703 = ( (~ Pz2)  &  (~ Pm) ) | ( (~ Pn)  &  (~ Pm) ) | ( (~ Pz2)  &  (~ Pd3) ) | ( (~ Pn)  &  (~ Pd3) ) ;
 assign n704 = ( n94  &  n352  &  (~ n573) ) | ( n335  &  n352  &  (~ n573) ) ;
 assign n705 = ( (~ Py0)  &  (~ Pv) ) | ( (~ Pw)  &  (~ Pv) ) | ( (~ Py0)  &  (~ Pd1) ) | ( (~ Pw)  &  (~ Pd1) ) ;
 assign n706 = ( (~ Pt)  &  (~ Ps) ) | ( (~ Pt)  &  (~ Po2) ) | ( (~ Ps)  &  (~ Pj2) ) | ( (~ Po2)  &  (~ Pj2) ) ;
 assign n707 = ( (~ Px1)  &  (~ Pp) ) | ( (~ Pq)  &  (~ Pp) ) | ( (~ Px1)  &  (~ Pa2) ) | ( (~ Pq)  &  (~ Pa2) ) ;
 assign n708 = ( (~ Pn)  &  (~ Pm) ) | ( (~ Pn)  &  (~ Pe3) ) | ( (~ Pm)  &  (~ Pa3) ) | ( (~ Pe3)  &  (~ Pa3) ) ;
 assign n709 = ( Ps4  &  n408 ) | ( Ps4  &  n517  &  Pr5 ) ;
 assign n710 = ( (~ Pq5)  &  (~ Po0) ) | ( (~ Po0)  &  (~ Pn0) ) | ( (~ Pq5)  &  n88 ) | ( (~ Pn0)  &  n88 ) ;
 assign n711 = ( (~ Pw4)  &  (~ Pu0) ) | ( (~ Pu0)  &  (~ Pt0) ) | ( (~ Pw4)  &  (~ Pr4) ) | ( (~ Pt0)  &  (~ Pr4) ) ;
 assign n712 = ( (~ Pr0)  &  (~ Pq0) ) | ( (~ Pr0)  &  (~ Pm4) ) | ( (~ Pq0)  &  (~ Ph4) ) | ( (~ Pm4)  &  (~ Ph4) ) ;
 assign n713 = ( (~ Pr5)  &  (~ Pp5) ) | ( (~ Pp5)  &  (~ Po0) ) | ( (~ Pr5)  &  (~ Pn0) ) | ( (~ Po0)  &  (~ Pn0) ) ;
 assign n714 = ( (~ Pq3)  &  (~ Pm3) ) | ( (~ Pq3)  &  (~ Pl0) ) | ( (~ Pm3)  &  (~ Pk0) ) | ( (~ Pl0)  &  (~ Pk0) ) ;
 assign n715 = ( Pq2  &  n229 ) | ( (~ Pq2)  &  n230 ) | ( n229  &  n230 ) ;
 assign n716 = ( (~ Po4) ) | ( n581 ) ;
 assign n717 = ( (~ Pj1) ) | ( n500 ) ;
 assign n720 = ( Pn3 ) | ( n611 ) | ( Pm3 ) ;
 assign n722 = ( (~ Pm2) ) | ( n617 ) ;
 assign n723 = ( (~ Pm4) ) | ( n257 ) ;
 assign n724 = ( Pm3  &  n609 ) | ( (~ Pm3)  &  n611 ) | ( n609  &  n611 ) ;
 assign n725 = ( (~ Pk4) ) | ( n260 ) ;
 assign n726 = ( (~ Pk2) ) | ( n295 ) ;
 assign n727 = ( (~ Ph4) ) | ( n578 ) ;
 assign n728 = ( Pn3 ) | ( Po3 ) | ( Pl3 ) | ( Pm3 ) ;
 assign n729 = ( (~ Pi2) ) | ( n298 ) ;
 assign n733 = ( (~ Pf2) ) | ( n588 ) ;
 assign n734 = ( (~ Ph1) ) | ( Pb ) | ( (~ n310) ) | ( (~ n365) ) ;
 assign n735 = ( Pf3  &  n265 ) | ( (~ Pf3)  &  n266 ) | ( n265  &  n266 ) ;
 assign n738 = ( Pc3 ) | ( n426 ) | ( Pd3 ) ;
 assign n741 = ( Pz ) | ( (~ Pd5) ) | ( n506 ) | ( (~ n631) ) ;
 assign n742 = ( Pb4 ) | ( n433 ) | ( Pa4 ) ;
 assign n743 = ( Pz1 ) | ( n464 ) | ( Py1 ) ;
 assign n744 = ( n414 ) | ( n460 ) | ( Py3 ) ;
 assign n745 = ( Py2 ) | ( n470 ) | ( Px2 ) ;
 assign n746 = ( (~ Px2)  &  n470 ) | ( Px2  &  n471 ) | ( n470  &  n471 ) ;
 assign n747 = ( n442 ) | ( n477 ) | ( Pw1 ) ;
 assign n749 = ( Pv3 ) | ( n460 ) | ( Pu3 ) ;
 assign n748 = ( (~ Pv3)  &  n749 ) | ( (~ Pu3)  &  n749 ) | ( n459  &  n749 ) ;
 assign n750 = ( Pu3  &  n459 ) | ( (~ Pu3)  &  n460 ) | ( n459  &  n460 ) ;
 assign n751 = ( Py2 ) | ( Pz2 ) | ( Pw2 ) | ( Px2 ) ;
 assign n753 = ( Pt1 ) | ( n477 ) | ( Ps1 ) ;
 assign n752 = ( (~ Pt1)  &  n753 ) | ( (~ Ps1)  &  n753 ) | ( n476  &  n753 ) ;
 assign n754 = ( Ps3 ) | ( n239 ) | ( Pr3 ) ;
 assign n755 = ( Ps1  &  n476 ) | ( (~ Ps1)  &  n477 ) | ( n476  &  n477 ) ;
 assign n759 = ( n609  &  n611 ) ;
 assign n760 = ( n273  &  n274 ) ;
 assign n763 = ( Pi1  &  (~ Pb)  &  n365  &  n538 ) ;
 assign n764 = ( (~ Pz)  &  Pe5  &  n508  &  n631 ) ;
 assign Pr6 = ( Pj1 ) ;
 assign Pp10 = ( Pg5 ) ;
 assign Pm6 = ( Pe1 ) ;
 assign Pl6 = ( Pa ) ;
 assign Pi10 = ( Pa5 ) ;
 assign Ph10 = ( Py ) ;


endmodule

