module table3 (
	i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, 
	i_8_, i_9_, i_10_, i_11_, i_12_, i_13_, o_0_, o_1_, o_2_, o_3_, 
	o_4_, o_5_, o_6_, o_7_, o_8_, o_9_, o_10_, o_11_, o_12_, o_13_);

input i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, i_8_, i_9_, i_10_, i_11_, i_12_, i_13_;

output o_0_, o_1_, o_2_, o_3_, o_4_, o_5_, o_6_, o_7_, o_8_, o_9_, o_10_, o_11_, o_12_, o_13_;

wire n1, n3, n4, n5, n6, n7, n8, n9, n2, n11, n12, n13, n14, n15, n16, n17, n10, n19, n20, n21, n22, n18, n24, n25, n23, n27, n28, n29, n30, n31, n32, n26, n34, n35, n36, n37, n38, n33, n40, n41, n42, n43, n44, n45, n46, n39, n48, n49, n50, n51, n52, n53, n54, n47, n56, n57, n58, n59, n60, n61, n62, n63, n55, n65, n66, n67, n68, n64, n69, n71, n72, n70, n75, n76, n73, n74, n80, n81, n78, n77, n82, n83, n84, n85, n86, n88, n91, n87, n92, n93, n94, n97, n95, n96, n100, n99, n98, n102, n101, n103, n105, n106, n104, n110, n107, n114, n111, n119, n118, n116, n120, n121, n122, n123, n124, n125, n127, n128, n126, n129, n130, n133, n131, n138, n136, n141, n142, n139, n140, n144, n145, n143, n149, n146, n154, n151, n152, n150, n156, n157, n155, n160, n159, n158, n163, n164, n161, n162, n165, n169, n170, n168, n174, n175, n173, n177, n178, n179, n176, n181, n182, n183, n180, n185, n184, n186, n193, n190, n195, n194, n198, n196, n201, n200, n199, n203, n204, n202, n205, n206, n207, n208, n212, n213, n215, n216, n214, n217, n218, n221, n222, n220, n219, n224, n225, n226, n223, n227, n231, n229, n230, n228, n233, n232, n237, n235, n241, n243, n246, n247, n245, n248, n251, n252, n254, n255, n253, n259, n257, n258, n256, n260, n261, n262, n263, n264, n266, n267, n265, n268, n270, n271, n272, n269, n273, n276, n277, n278, n280, n282, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n338, n339, n340, n335, n341, n342, n343, n344, n345, n346, n347, n348, n350, n351, n352, n353, n354, n355, n357, n358, n359, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371;

assign o_0_ = ( (~ n70) ) ;
 assign o_1_ = ( (~ n69) ) ;
 assign o_2_ = ( (~ n64) ) ;
 assign o_3_ = ( (~ n55) ) ;
 assign o_4_ = ( (~ n47) ) ;
 assign o_5_ = ( (~ n39) ) ;
 assign o_6_ = ( (~ n33) ) ;
 assign o_7_ = ( (~ n26) ) ;
 assign o_8_ = ( (~ n23) ) ;
 assign o_9_ = ( (~ n18) ) ;
 assign o_10_ = ( (~ n10) ) ;
 assign o_11_ = ( (~ n269) ) ;
 assign o_12_ = ( (~ n2) ) ;
 assign o_13_ = ( (~ n1) ) ;
 assign n1 = ( n260  &  n62  &  n261  &  n262  &  n263  &  n264 ) ;
 assign n3 = ( n320  &  n98 ) ;
 assign n4 = ( n120  &  n121  &  n122  &  n123  &  n124  &  n125 ) ;
 assign n5 = ( n277 ) | ( n179 ) | ( n106 ) ;
 assign n6 = ( n170 ) | ( n152 ) ;
 assign n7 = ( n203  &  n204  &  n202 ) | ( n203  &  n204  &  n195 ) ;
 assign n8 = ( n350  &  n60  &  n85  &  n351 ) ;
 assign n9 = ( n343  &  n339  &  n25  &  n314  &  n84  &  n83  &  n344  &  n352 ) ;
 assign n2 = ( n3  &  n4  &  n5  &  n6  &  n7  &  n8  &  n9 ) ;
 assign n11 = ( n353  &  n77  &  n347  &  n354 ) ;
 assign n12 = ( n314  &  n25 ) ;
 assign n13 = ( n4  &  n129  &  n130 ) ;
 assign n14 = ( n179 ) | ( n177 ) | ( n95 ) | ( n229 ) ;
 assign n15 = ( n97  &  n95 ) | ( n97  &  n96 ) ;
 assign n16 = ( n280 ) | ( n151 ) ;
 assign n17 = ( n341  &  n342 ) ;
 assign n10 = ( n8  &  n11  &  n12  &  n13  &  n14  &  n15  &  n16  &  n17 ) ;
 assign n19 = ( n71  &  n15  &  n29 ) ;
 assign n20 = ( n82  &  n83  &  n84  &  n85  &  n86  &  n77 ) ;
 assign n21 = ( n75  &  n76  &  n73 ) | ( n75  &  n76  &  n74 ) ;
 assign n22 = ( n286 ) | ( n92 ) ;
 assign n18 = ( n19  &  n20  &  n21  &  n16  &  n22  &  n12 ) ;
 assign n24 = ( n179 ) | ( n181 ) | ( n266 ) ;
 assign n25 = ( n298 ) | ( n313 ) | ( n202 ) ;
 assign n23 = ( n24  &  n19  &  n25  &  n16 ) ;
 assign n27 = ( n6  &  n37  &  n38 ) ;
 assign n28 = ( i_7_ ) | ( n319 ) ;
 assign n29 = ( n87  &  n93 ) | ( n92  &  n93 ) | ( n87  &  n94 ) | ( n92  &  n94 ) ;
 assign n30 = ( (~ i_8_) ) | ( n266 ) | ( n317 ) ;
 assign n31 = ( i_8_ ) | ( n319 ) ;
 assign n32 = ( n222 ) | ( n106 ) ;
 assign n26 = ( n27  &  n3  &  n28  &  n29  &  n30  &  n31  &  n16  &  n32 ) ;
 assign n34 = ( (~ i_6_) ) | ( i_7_ ) | ( (~ i_8_) ) | ( n92 ) | ( n170 ) | ( n276 ) ;
 assign n35 = ( n32  &  n16  &  n103 ) ;
 assign n36 = ( n170 ) | ( n178 ) | ( n230 ) ;
 assign n37 = ( n246 ) | ( n170 ) | ( n311 ) ;
 assign n38 = ( n170 ) | ( n312 ) | ( n178 ) | ( i_7_ ) | ( i_8_ ) | ( i_9_ ) ;
 assign n33 = ( n34  &  n19  &  n35  &  n36  &  n37  &  n38 ) ;
 assign n40 = ( (~ i_11_) ) | ( n156 ) | ( n246 ) | ( n299 ) | ( n304 ) ;
 assign n41 = ( n106 ) | ( n324 ) ;
 assign n42 = ( (~ i_8_) ) | ( n317 ) | ( n321 ) ;
 assign n43 = ( (~ i_3_) ) | ( (~ i_5_) ) | ( (~ i_13_) ) | ( n165 ) ;
 assign n44 = ( n92 ) | ( n128 ) | ( (~ n133) ) ;
 assign n45 = ( n163  &  n164  &  n161 ) | ( n163  &  n164  &  n162 ) ;
 assign n46 = ( n252  &  n13  &  n333  &  n158  &  n270  &  n150 ) ;
 assign n39 = ( n40  &  n41  &  n42  &  n5  &  n43  &  n44  &  n45  &  n46 ) ;
 assign n48 = ( n141  &  n142  &  n139 ) | ( n141  &  n142  &  n140 ) ;
 assign n49 = ( n212  &  n213  &  n182 ) | ( n212  &  n213  &  n152 ) ;
 assign n50 = ( n333  &  n345  &  n34  &  n27  &  n332  &  n346  &  n5  &  n331 ) ;
 assign n51 = ( n7  &  n21  &  n205  &  n20  &  n206  &  n207 ) ;
 assign n52 = ( n196  &  n335  &  n150  &  n72  &  n61  &  n129  &  n347  &  n348 ) ;
 assign n53 = ( n92 ) | ( n110 ) | ( n128 ) ;
 assign n54 = ( n351  &  n350  &  n31 ) ;
 assign n47 = ( n48  &  n49  &  n50  &  n51  &  n52  &  n53  &  n3  &  n54 ) ;
 assign n56 = ( n93 ) | ( n165 ) ;
 assign n57 = ( i_0_ ) | ( (~ i_2_) ) | ( i_3_ ) | ( n159 ) ;
 assign n58 = ( n179  &  (~ n235)  &  n241 ) | ( n228  &  (~ n235)  &  n241 ) ;
 assign n59 = ( n223  &  n136  &  n227 ) ;
 assign n60 = ( n65  &  n49  &  n218  &  n29 ) ;
 assign n61 = ( n102 ) | ( n127 ) | ( n128 ) ;
 assign n62 = ( n182 ) | ( n305 ) ;
 assign n63 = ( n354  &  n353  &  n142 ) ;
 assign n55 = ( n56  &  n57  &  n58  &  n59  &  n60  &  n61  &  n62  &  n63 ) ;
 assign n65 = ( n217  &  n110 ) | ( n217  &  n174 ) ;
 assign n66 = ( n41  &  n53  &  n56  &  n158  &  n245  &  (~ n248) ) ;
 assign n67 = ( n320  &  n50  &  n58 ) ;
 assign n68 = ( n31  &  n98 ) ;
 assign n64 = ( n65  &  n59  &  n40  &  n52  &  n66  &  n67  &  n68 ) ;
 assign n69 = ( n66  &  n223  &  n251  &  n252 ) ;
 assign n71 = ( n286 ) | ( n298 ) ;
 assign n72 = ( n334  &  n22  &  n28 ) ;
 assign n70 = ( n51  &  n67  &  n68  &  n71  &  n29  &  n72 ) ;
 assign n75 = ( n293 ) | ( n102 ) | ( n259 ) | ( n292 ) ;
 assign n76 = ( n288 ) | ( n289 ) ;
 assign n73 = ( i_4_ ) | ( n259 ) | ( n246 ) ;
 assign n74 = ( i_10_ ) | ( (~ i_11_) ) | ( (~ i_12_) ) | ( (~ i_13_) ) ;
 assign n80 = ( n118 ) | ( (~ n237) ) ;
 assign n81 = ( n287 ) | ( n301 ) | ( n306 ) ;
 assign n78 = ( n246 ) | ( n300 ) ;
 assign n77 = ( n80  &  n81  &  n78 ) | ( n80  &  n81  &  (~ n193) ) ;
 assign n82 = ( i_10_ ) | ( n297 ) | ( n298 ) | ( n170 ) | ( n304 ) ;
 assign n83 = ( n302 ) | ( n303 ) ;
 assign n84 = ( n157 ) | ( n301 ) ;
 assign n85 = ( n139 ) | ( n298 ) | ( n182 ) ;
 assign n86 = ( n355  &  n300 ) | ( n355  &  n185 ) | ( n355  &  n307 ) ;
 assign n88 = ( n291 ) | ( n297 ) ;
 assign n91 = ( i_6_ ) | ( n299 ) | ( n308 ) ;
 assign n87 = ( n88  &  n91 ) | ( n91  &  (~ n133) ) | ( n88  &  (~ n237) ) | ( (~ n133)  &  (~ n237) ) ;
 assign n92 = ( (~ i_2_) ) | ( n282 ) ;
 assign n93 = ( (~ i_3_) ) | ( (~ i_4_) ) ;
 assign n94 = ( (~ i_10_) ) | ( n246 ) | ( n309 ) ;
 assign n97 = ( (~ i_13_) ) | ( n88 ) | ( n127 ) | ( n170 ) ;
 assign n95 = ( i_4_ ) | ( i_3_ ) ;
 assign n96 = ( (~ i_10_) ) | ( n127 ) | ( n233 ) ;
 assign n100 = ( (~ i_10_) ) | ( n93 ) | ( n293 ) | ( n309 ) ;
 assign n99 = ( n308 ) | ( n144 ) ;
 assign n98 = ( n100  &  n99 ) | ( n100  &  (~ n237) ) ;
 assign n102 = ( i_5_ ) | ( n93 ) ;
 assign n101 = ( n102  &  n93 ) | ( n88  &  n93 ) | ( n102  &  n91 ) | ( n88  &  n91 ) ;
 assign n103 = ( n101  &  n179 ) | ( n298  &  n179 ) | ( n101  &  n322 ) | ( n298  &  n322 ) ;
 assign n105 = ( i_7_ ) | ( (~ i_9_) ) ;
 assign n106 = ( (~ i_5_) ) | ( (~ n149) ) ;
 assign n104 = ( n105 ) | ( n106 ) | ( n74 ) | ( i_6_ ) ;
 assign n110 = ( i_5_ ) | ( (~ n149) ) ;
 assign n107 = ( (~ i_8_) ) | ( n110 ) | ( (~ n114) ) ;
 assign n114 = ( (~ i_9_)  &  (~ n161) ) ;
 assign n111 = ( n114  &  (~ n266) ) | ( (~ n229)  &  (~ n266)  &  (~ n267) ) ;
 assign n119 = ( i_9_ ) | ( n326 ) | ( n169 ) ;
 assign n118 = ( n298 ) | ( n303 ) ;
 assign n116 = ( (~ i_13_)  &  n119 ) | ( n119  &  n118 ) ;
 assign n120 = ( n139 ) | ( n298 ) | ( n106 ) ;
 assign n121 = ( (~ n193) ) | ( n287 ) | ( n306 ) ;
 assign n122 = ( n183 ) | ( n74 ) | ( n259 ) | ( n93 ) ;
 assign n123 = ( n161 ) | ( n105 ) | ( n92 ) | ( n182 ) ;
 assign n124 = ( n358  &  n359  &  n289 ) | ( n358  &  n359  &  n156 ) ;
 assign n125 = ( n357  &  n288 ) | ( n278  &  n288 ) | ( n357  &  n118 ) | ( n278  &  n118 ) ;
 assign n127 = ( i_2_ ) | ( n282 ) ;
 assign n128 = ( n304 ) | ( n230 ) ;
 assign n126 = ( n110 ) | ( n127 ) | ( n128 ) ;
 assign n129 = ( n328  &  n329  &  n126 ) ;
 assign n130 = ( n346  &  n339  &  n93 ) | ( n346  &  n339  &  n327 ) ;
 assign n133 = ( (~ i_5_)  &  n237 ) ;
 assign n131 = ( (~ n298)  &  (~ n322) ) | ( n133  &  (~ n298)  &  (~ n313) ) ;
 assign n138 = ( (~ n131)  &  n170 ) | ( (~ n131)  &  n280  &  n324 ) ;
 assign n136 = ( n96  &  n138 ) | ( n138  &  (~ n149) ) ;
 assign n141 = ( n278 ) | ( n300 ) | ( n301 ) ;
 assign n142 = ( (~ n133) ) | ( n174 ) ;
 assign n139 = ( n296 ) | ( n297 ) ;
 assign n140 = ( n151 ) | ( n298 ) ;
 assign n144 = ( i_6_ ) | ( n299 ) | ( n127 ) ;
 assign n145 = ( i_11_ ) | ( n229 ) ;
 assign n143 = ( n144 ) | ( n145 ) | ( i_5_ ) | ( i_3_ ) ;
 assign n149 = ( i_3_  &  (~ i_4_) ) ;
 assign n146 = ( (~ n99)  &  n149 ) | ( n149  &  (~ n165) ) ;
 assign n154 = ( n94  &  n96 ) | ( n95  &  n96 ) | ( n94  &  (~ n237) ) | ( n95  &  (~ n237) ) ;
 assign n151 = ( (~ i_5_) ) | ( n95 ) ;
 assign n152 = ( n179 ) | ( n313 ) ;
 assign n150 = ( (~ n146)  &  n154  &  n151 ) | ( (~ n146)  &  n154  &  n152 ) ;
 assign n156 = ( (~ i_6_) ) | ( n93 ) ;
 assign n157 = ( n300 ) | ( n179 ) ;
 assign n155 = ( n156 ) | ( n157 ) ;
 assign n160 = ( n139 ) | ( n170 ) | ( n327 ) ;
 assign n159 = ( n299 ) | ( n307 ) | ( n145 ) ;
 assign n158 = ( n160  &  n92 ) | ( n160  &  n159 ) ;
 assign n163 = ( n151 ) | ( n139 ) | ( n327 ) ;
 assign n164 = ( n246 ) | ( n202 ) | ( n259 ) | ( n292 ) ;
 assign n161 = ( i_10_ ) | ( n284 ) ;
 assign n162 = ( n95 ) | ( n92 ) ;
 assign n165 = ( n290 ) | ( n144 ) ;
 assign n169 = ( i_6_ ) | ( n296 ) ;
 assign n170 = ( (~ i_5_) ) | ( (~ n237) ) ;
 assign n168 = ( (~ i_7_) ) | ( (~ i_9_) ) | ( n169 ) | ( n170 ) ;
 assign n174 = ( n246 ) | ( n313 ) ;
 assign n175 = ( n92 ) | ( n297 ) | ( i_10_ ) | ( n229 ) ;
 assign n173 = ( n174  &  n175 ) ;
 assign n177 = ( (~ i_7_) ) | ( n267 ) ;
 assign n178 = ( n229 ) | ( n246 ) ;
 assign n179 = ( i_1_ ) | ( n294 ) ;
 assign n176 = ( n177  &  n179 ) | ( n178  &  n179 ) | ( n177  &  n161 ) | ( n178  &  n161 ) ;
 assign n181 = ( n284 ) | ( n315 ) ;
 assign n182 = ( (~ i_5_) ) | ( n93 ) ;
 assign n183 = ( i_0_ ) | ( i_1_ ) ;
 assign n180 = ( n181 ) | ( n182 ) | ( n183 ) | ( i_7_ ) ;
 assign n185 = ( (~ i_13_) ) | ( n278 ) ;
 assign n184 = ( n88 ) | ( n185 ) | ( n110 ) ;
 assign n186 = ( (~ n168)  &  (~ n278) ) | ( (~ n102)  &  (~ n278)  &  (~ n313) ) ;
 assign n193 = ( n237  &  i_6_ ) ;
 assign n190 = ( (~ n157)  &  n193 ) | ( n193  &  (~ n289) ) ;
 assign n195 = ( (~ i_6_) ) | ( n282 ) | ( n296 ) ;
 assign n194 = ( (~ n133) ) | ( n195 ) ;
 assign n198 = ( i_3_ ) | ( n276 ) | ( n326 ) ;
 assign n196 = ( (~ i_6_)  &  n198 ) | ( n78  &  n198 ) | ( (~ n149)  &  n198 ) ;
 assign n201 = ( n246 ) | ( n181 ) | ( n106 ) ;
 assign n200 = ( n284 ) | ( n325 ) ;
 assign n199 = ( n201  &  n127 ) | ( n201  &  n200 ) ;
 assign n203 = ( n278 ) | ( n313 ) | ( n110 ) ;
 assign n204 = ( n127  &  n151 ) | ( n231  &  n151 ) | ( n127  &  n222 ) | ( n231  &  n222 ) ;
 assign n202 = ( i_5_ ) | ( n95 ) ;
 assign n205 = ( n341  &  n342  &  n343  &  n344  &  n199 ) ;
 assign n206 = ( n95 ) | ( n293 ) ;
 assign n207 = ( n14  &  (~ n149) ) | ( n14  &  n327 ) ;
 assign n208 = ( (~ n91)  &  (~ n162) ) | ( (~ i_6_)  &  (~ n162)  &  (~ n300) ) ;
 assign n212 = ( n106  &  (~ n208) ) | ( (~ n208)  &  n277 ) | ( (~ n208)  &  n298 ) ;
 assign n213 = ( n93  &  n94 ) | ( n94  &  n96 ) | ( n93  &  (~ n149) ) | ( n96  &  (~ n149) ) ;
 assign n215 = ( i_6_ ) | ( (~ i_7_) ) | ( i_8_ ) ;
 assign n216 = ( i_6_ ) | ( i_7_ ) | ( (~ i_8_) ) ;
 assign n214 = ( n215  &  n216  &  i_6_ ) | ( n215  &  n216  &  n105 ) ;
 assign n217 = ( n170 ) | ( n327 ) | ( n214 ) | ( n296 ) ;
 assign n218 = ( n366  &  n127 ) | ( n366  &  n311 ) | ( n366  &  n110 ) ;
 assign n221 = ( i_7_ ) | ( n220 ) ;
 assign n222 = ( n278 ) | ( n316 ) | ( n215 ) ;
 assign n220 = ( n298 ) | ( n309 ) | ( i_6_ ) | ( i_10_ ) ;
 assign n219 = ( n221  &  n222  &  i_8_ ) | ( n221  &  n222  &  n220 ) ;
 assign n224 = ( n219  &  n93 ) | ( n182  &  n93 ) | ( n219  &  n99 ) | ( n182  &  n99 ) ;
 assign n225 = ( n362  &  n276 ) | ( n362  &  n92 ) | ( n362  &  n321 ) ;
 assign n226 = ( n94  &  n363 ) | ( (~ n237)  &  n363 ) ;
 assign n223 = ( n224  &  n225  &  n226 ) ;
 assign n227 = ( (~ n237)  &  n364  &  n365 ) | ( n293  &  n364  &  n365 ) ;
 assign n231 = ( n102 ) | ( n311 ) ;
 assign n229 = ( (~ i_12_) ) | ( (~ i_13_) ) ;
 assign n230 = ( (~ i_6_) ) | ( n295 ) ;
 assign n228 = ( n231  &  n229 ) | ( n231  &  n182 ) | ( n231  &  n230 ) ;
 assign n233 = ( i_11_ ) | ( i_12_ ) | ( (~ i_13_) ) ;
 assign n232 = ( (~ i_10_) ) | ( (~ n193) ) | ( n233 ) ;
 assign n237 = ( (~ i_3_)  &  i_4_ ) ;
 assign n235 = ( (~ n232)  &  (~ n327) ) | ( (~ n161)  &  n237  &  (~ n327) ) ;
 assign n241 = ( (~ n133) ) | ( n246 ) | ( n310 ) ;
 assign n243 = ( (~ n91)  &  (~ n95) ) ;
 assign n246 = ( (~ i_2_) ) | ( n183 ) ;
 assign n247 = ( i_8_  &  i_7_ ) ;
 assign n245 = ( n74 ) | ( n246 ) | ( n95 ) | ( n247 ) ;
 assign n248 = ( n243  &  (~ n327) ) | ( (~ n88)  &  (~ n202)  &  (~ n327) ) ;
 assign n251 = ( n61  &  n78 ) | ( n61  &  n156 ) ;
 assign n252 = ( n143  &  n48  &  n136 ) ;
 assign n254 = ( n183  &  (~ n237) ) | ( (~ n193)  &  (~ n237) ) | ( n183  &  n298 ) | ( (~ n193)  &  n298 ) ;
 assign n255 = ( i_3_  &  n302 ) | ( (~ i_6_)  &  n302 ) | ( n179  &  n302 ) ;
 assign n253 = ( n254  &  n255 ) ;
 assign n259 = ( (~ i_7_) ) | ( (~ i_8_) ) ;
 assign n257 = ( n368  &  n369  &  n370 ) ;
 assign n258 = ( (~ i_10_)  &  n367 ) | ( n301  &  n367 ) | ( n306  &  n367 ) ;
 assign n256 = ( n76  &  n259 ) | ( n76  &  n257  &  n258 ) ;
 assign n260 = ( n307 ) | ( n310 ) | ( i_3_ ) | ( n183 ) ;
 assign n261 = ( (~ i_7_) ) | ( n253 ) | ( n290 ) | ( n315 ) ;
 assign n262 = ( (~ i_9_)  &  n73 ) | ( n73  &  n256 ) | ( (~ i_9_)  &  n276 ) | ( n256  &  n276 ) ;
 assign n263 = ( (~ n237) ) | ( n293 ) ;
 assign n264 = ( n205  &  n335  &  n345  &  n12  &  n29  &  n196 ) ;
 assign n266 = ( (~ i_7_) ) | ( (~ n149) ) ;
 assign n267 = ( (~ i_8_) ) | ( i_10_ ) | ( (~ i_11_) ) ;
 assign n265 = ( n266 ) | ( n267 ) | ( n178 ) ;
 assign n268 = ( (~ i_3_) ) | ( n76 ) ;
 assign n270 = ( n330  &  n155  &  n331  &  n332 ) ;
 assign n271 = ( (~ i_3_)  &  n95 ) | ( (~ i_3_)  &  n293 ) | ( n95  &  n327 ) | ( n293  &  n327 ) ;
 assign n272 = ( n371  &  n365  &  n329  &  n328  &  n355  &  n82  &  n334  &  n36 ) ;
 assign n269 = ( n9  &  n199  &  n11  &  n270  &  n19  &  n271  &  n272 ) ;
 assign n273 = ( (~ i_9_) ) | ( i_10_ ) ;
 assign n276 = ( (~ i_11_) ) | ( n229 ) | ( n273 ) ;
 assign n277 = ( n276 ) | ( n216 ) ;
 assign n278 = ( (~ i_0_) ) | ( i_1_ ) | ( (~ i_2_) ) ;
 assign n280 = ( n277 ) | ( n278 ) ;
 assign n282 = ( i_0_ ) | ( (~ i_1_) ) ;
 assign n284 = ( (~ i_11_) ) | ( n229 ) ;
 assign n285 = ( i_8_ ) | ( n273 ) | ( n284 ) ;
 assign n286 = ( i_7_ ) | ( (~ n237) ) | ( n285 ) ;
 assign n287 = ( (~ i_10_) ) | ( n259 ) ;
 assign n288 = ( i_4_ ) | ( (~ i_6_) ) ;
 assign n289 = ( n92 ) | ( n287 ) | ( n233 ) ;
 assign n290 = ( (~ i_11_) ) | ( i_12_ ) ;
 assign n291 = ( i_10_ ) | ( n290 ) ;
 assign n292 = ( (~ i_6_) ) | ( i_13_ ) | ( n291 ) ;
 assign n293 = ( i_2_ ) | ( n183 ) ;
 assign n294 = ( (~ i_0_) ) | ( i_2_ ) ;
 assign n295 = ( i_11_ ) | ( i_10_ ) ;
 assign n296 = ( i_12_ ) | ( i_13_ ) | ( n295 ) ;
 assign n297 = ( i_6_ ) | ( n259 ) ;
 assign n298 = ( (~ i_1_) ) | ( n294 ) ;
 assign n299 = ( i_10_ ) | ( n259 ) ;
 assign n300 = ( n290 ) | ( n299 ) ;
 assign n301 = ( (~ i_6_) ) | ( n95 ) ;
 assign n302 = ( n278 ) | ( n93 ) ;
 assign n303 = ( i_12_ ) | ( n177 ) ;
 assign n304 = ( i_12_ ) | ( i_13_ ) ;
 assign n305 = ( n278 ) | ( n139 ) ;
 assign n306 = ( n233 ) | ( n179 ) ;
 assign n307 = ( (~ i_4_) ) | ( i_5_ ) | ( i_6_ ) ;
 assign n308 = ( (~ i_11_) ) | ( i_13_ ) ;
 assign n309 = ( i_11_ ) | ( n304 ) ;
 assign n310 = ( i_10_ ) | ( n145 ) ;
 assign n311 = ( n297 ) | ( n310 ) ;
 assign n312 = ( i_6_ ) | ( n295 ) ;
 assign n313 = ( n304 ) | ( n312 ) ;
 assign n314 = ( n246 ) | ( n231 ) ;
 assign n315 = ( (~ i_8_) ) | ( n273 ) ;
 assign n316 = ( n273 ) | ( n309 ) ;
 assign n317 = ( (~ n114) ) | ( n179 ) ;
 assign n318 = ( (~ i_4_) ) | ( (~ i_5_) ) | ( i_6_ ) ;
 assign n319 = ( i_3_ ) | ( i_10_ ) | ( n294 ) | ( n309 ) | ( n318 ) ;
 assign n320 = ( n88 ) | ( n127 ) | ( (~ n133) ) ;
 assign n321 = ( i_7_ ) | ( (~ n149) ) ;
 assign n322 = ( n285 ) | ( n321 ) ;
 assign n323 = ( (~ i_8_) ) | ( n105 ) ;
 assign n324 = ( n74 ) | ( n127 ) | ( n323 ) ;
 assign n325 = ( i_10_ ) | ( n93 ) ;
 assign n326 = ( i_7_ ) | ( i_8_ ) | ( n298 ) ;
 assign n327 = ( (~ i_0_) ) | ( (~ i_1_) ) | ( (~ i_2_) ) ;
 assign n328 = ( i_8_ ) | ( n106 ) | ( n220 ) ;
 assign n329 = ( n106 ) | ( n221 ) ;
 assign n330 = ( n92 ) | ( n311 ) | ( n110 ) ;
 assign n331 = ( n277 ) | ( n140 ) ;
 assign n332 = ( i_8_ ) | ( n266 ) | ( n317 ) ;
 assign n333 = ( n12  &  n35  &  n24  &  n30 ) ;
 assign n334 = ( n277 ) | ( n92 ) | ( n170 ) ;
 assign n338 = ( n45  &  n170 ) | ( n45  &  n305 ) ;
 assign n339 = ( n293 ) | ( n200 ) ;
 assign n340 = ( n173  &  n176 ) | ( n176  &  n202 ) | ( n173  &  (~ n237) ) | ( n202  &  (~ n237) ) ;
 assign n335 = ( n180  &  n184  &  (~ n186)  &  (~ n190)  &  n194  &  n338  &  n339  &  n340 ) ;
 assign n341 = ( n293 ) | ( n102 ) | ( n313 ) ;
 assign n342 = ( i_7_ ) | ( n285 ) | ( n302 ) ;
 assign n343 = ( n74 ) | ( n179 ) | ( i_7_ ) | ( n95 ) ;
 assign n344 = ( i_8_ ) | ( n95 ) | ( n317 ) ;
 assign n345 = ( n42  &  n36  &  n15 ) ;
 assign n346 = ( n151 ) | ( n324 ) ;
 assign n347 = ( n95 ) | ( n246 ) | ( n310 ) ;
 assign n348 = ( n361  &  n330 ) ;
 assign n350 = ( (~ i_6_) ) | ( (~ n149) ) | ( n157 ) ;
 assign n351 = ( n305 ) | ( n106 ) ;
 assign n352 = ( n265  &  n268  &  n150  &  n361  &  n16  &  n241 ) ;
 assign n353 = ( n151 ) | ( n221 ) ;
 assign n354 = ( n169 ) | ( n140 ) | ( i_8_ ) | ( i_9_ ) ;
 assign n355 = ( n151 ) | ( n305 ) ;
 assign n357 = ( n104  &  n107  &  (~ n111)  &  n322 ) ;
 assign n358 = ( (~ i_4_) ) | ( n276 ) | ( n326 ) ;
 assign n359 = ( i_5_ ) | ( n116 ) | ( i_4_ ) ;
 assign n361 = ( n280 ) | ( n182 ) ;
 assign n362 = ( (~ i_1_) ) | ( i_2_ ) | ( i_3_ ) | ( n74 ) | ( n318 ) | ( n323 ) ;
 assign n363 = ( n179  &  n106 ) | ( n200  &  n106 ) | ( n179  &  n152 ) | ( n200  &  n152 ) ;
 assign n364 = ( n127 ) | ( n311 ) | ( n202 ) ;
 assign n365 = ( n293 ) | ( n145 ) | ( n325 ) ;
 assign n366 = ( n316 ) | ( n215 ) | ( n140 ) ;
 assign n367 = ( n291 ) | ( n185 ) | ( n307 ) ;
 assign n368 = ( i_3_ ) | ( (~ i_5_) ) | ( n169 ) | ( n278 ) ;
 assign n369 = ( (~ i_4_) ) | ( i_5_ ) | ( n292 ) | ( n293 ) ;
 assign n370 = ( n296 ) | ( n298 ) | ( n318 ) ;
 assign n371 = ( n296 ) | ( n127 ) | ( i_5_ ) | ( n288 ) ;


endmodule

