module e64 (
	i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, 
	i_8_, i_9_, i_10_, i_11_, i_12_, i_13_, i_14_, i_15_, i_16_, i_17_, 
	i_18_, i_19_, i_20_, i_21_, i_22_, i_23_, i_24_, i_25_, i_26_, i_27_, 
	i_28_, i_29_, i_30_, i_31_, i_32_, i_33_, i_34_, i_35_, i_36_, i_37_, 
	i_38_, i_39_, i_40_, i_41_, i_42_, i_43_, i_44_, i_45_, i_46_, i_47_, 
	i_48_, i_49_, i_50_, i_51_, i_52_, i_53_, i_54_, i_55_, i_56_, i_57_, 
	i_58_, i_59_, i_60_, i_61_, i_62_, i_63_, i_64_, o_0_, o_1_, o_2_, 
	o_3_, o_4_, o_5_, o_6_, o_7_, o_8_, o_9_, o_10_, o_11_, o_12_, 
	o_13_, o_14_, o_15_, o_16_, o_17_, o_18_, o_19_, o_20_, o_21_, o_22_, 
	o_23_, o_24_, o_25_, o_26_, o_27_, o_28_, o_29_, o_30_, o_31_, o_32_, 
	o_33_, o_34_, o_35_, o_36_, o_37_, o_38_, o_39_, o_40_, o_41_, o_42_, 
	o_43_, o_44_, o_45_, o_46_, o_47_, o_48_, o_49_, o_50_, o_51_, o_52_, 
	o_53_, o_54_, o_55_, o_56_, o_57_, o_58_, o_59_, o_60_, o_61_, o_62_, 
	o_63_, o_64_);

input i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, i_8_, i_9_, i_10_, i_11_, i_12_, i_13_, i_14_, i_15_, i_16_, i_17_, i_18_, i_19_, i_20_, i_21_, i_22_, i_23_, i_24_, i_25_, i_26_, i_27_, i_28_, i_29_, i_30_, i_31_, i_32_, i_33_, i_34_, i_35_, i_36_, i_37_, i_38_, i_39_, i_40_, i_41_, i_42_, i_43_, i_44_, i_45_, i_46_, i_47_, i_48_, i_49_, i_50_, i_51_, i_52_, i_53_, i_54_, i_55_, i_56_, i_57_, i_58_, i_59_, i_60_, i_61_, i_62_, i_63_, i_64_;

output o_0_, o_1_, o_2_, o_3_, o_4_, o_5_, o_6_, o_7_, o_8_, o_9_, o_10_, o_11_, o_12_, o_13_, o_14_, o_15_, o_16_, o_17_, o_18_, o_19_, o_20_, o_21_, o_22_, o_23_, o_24_, o_25_, o_26_, o_27_, o_28_, o_29_, o_30_, o_31_, o_32_, o_33_, o_34_, o_35_, o_36_, o_37_, o_38_, o_39_, o_40_, o_41_, o_42_, o_43_, o_44_, o_45_, o_46_, o_47_, o_48_, o_49_, o_50_, o_51_, o_52_, o_53_, o_54_, o_55_, o_56_, o_57_, o_58_, o_59_, o_60_, o_61_, o_62_, o_63_, o_64_;

wire n4, n5, n6, n7, n8, n10, n12, n13, n14, n16, n18, n20, n22, n19, n26, n31, n32, n33, n35, n36, n37, n38, n30, n45, n46, n48, n44, n50, n51, n52, n53, n54, n55, n49, n61, n64, n65, n66, n67, n60, n70, n71, n72, n73, n68, n76, n77, n78, n79, n80, n74, n82, n83, n81, n86, n87, n85, n89, n88, n91, n98, n99, n101, n97, n104, n105, n106, n102, n108, n110, n112, n117, n118, n115, n121, n125, n127, n124, n129, n132, n135, n133, n137, n138, n139, n136, n142, n143, n144, n141, n149, n148, n151, n154, n160, n161, n158, n163, n164, n165, n167, n162, n170, n171, n168, n174, n175, n172, n179, n180, n181, n178, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n195, n196, n197, n198, n199, n200, n202, n203, n204, n205, n208, n212, n214, n215, n216, n219, n221, n222, n223, n224, n225, n226, n227, n228, n229, n231, n232;

assign o_0_ = ( (~ n178) ) ;
 assign o_1_ = ( i_5_  &  (~ n71)  &  (~ n83)  &  (~ n181) ) ;
 assign o_2_ = ( (~ n172) ) ;
 assign o_3_ = ( (~ n168) ) ;
 assign o_4_ = ( i_15_  &  i_29_ ) ;
 assign o_6_ = ( i_14_  &  (~ i_15_)  &  n112 ) ;
 assign o_7_ = ( (~ i_15_)  &  i_43_  &  n129 ) ;
 assign o_8_ = ( (~ n162) ) ;
 assign o_9_ = ( (~ n158) ) ;
 assign o_10_ = ( (~ i_15_)  &  i_28_  &  i_29_  &  (~ i_37_) ) ;
 assign o_11_ = ( (~ i_15_)  &  i_29_  &  i_37_ ) ;
 assign o_12_ = ( i_6_  &  (~ i_15_)  &  (~ i_24_)  &  n14  &  (~ n144)  &  (~ n195) ) ;
 assign o_13_ = ( i_41_  &  n151  &  n18  &  n132 ) ;
 assign o_14_ = ( i_50_  &  n154 ) ;
 assign o_15_ = ( i_10_  &  (~ i_58_)  &  n112  &  (~ n198) ) ;
 assign o_16_ = ( (~ i_3_)  &  i_26_  &  n10  &  n151 ) ;
 assign o_17_ = ( i_3_  &  n6  &  n8  &  (~ n71)  &  n151 ) ;
 assign o_18_ = ( (~ n148) ) ;
 assign o_19_ = ( i_64_  &  (~ n223)  &  (~ n229) ) ;
 assign o_20_ = ( i_51_  &  (~ n143)  &  (~ n144)  &  (~ n226) ) ;
 assign o_21_ = ( (~ n141) ) ;
 assign o_22_ = ( (~ n136) ) ;
 assign o_23_ = ( (~ n133) ) ;
 assign o_24_ = ( (~ i_10_)  &  i_11_  &  (~ i_14_)  &  n7  &  n129  &  n132  &  (~ n183) ) ;
 assign o_25_ = ( i_24_  &  (~ i_25_)  &  n4  &  n121 ) ;
 assign o_26_ = ( (~ n124) ) ;
 assign o_27_ = ( i_13_  &  (~ i_16_)  &  (~ i_20_)  &  (~ i_52_)  &  (~ n232) ) ;
 assign o_28_ = ( n121  &  n4  &  i_25_ ) ;
 assign o_29_ = ( (~ i_46_)  &  i_60_  &  n12  &  (~ n183) ) ;
 assign o_30_ = ( i_52_  &  (~ n232) ) ;
 assign o_31_ = ( (~ n115) ) ;
 assign o_32_ = ( i_46_  &  n12  &  (~ n183) ) ;
 assign o_33_ = ( i_39_  &  (~ i_40_)  &  n12 ) ;
 assign o_34_ = ( i_58_  &  n112  &  (~ n198) ) ;
 assign o_35_ = ( (~ i_0_)  &  i_4_  &  (~ i_41_)  &  n110  &  (~ n187)  &  (~ n231) ) ;
 assign o_36_ = ( (~ i_60_)  &  i_61_  &  (~ i_62_)  &  n26  &  n108 ) ;
 assign o_37_ = ( (~ n102) ) ;
 assign o_38_ = ( (~ n97) ) ;
 assign o_39_ = ( (~ i_40_)  &  (~ i_41_)  &  i_42_  &  (~ i_50_)  &  (~ n101)  &  (~ n187)  &  (~ n214) ) ;
 assign o_40_ = ( i_54_  &  (~ n45)  &  (~ n46)  &  (~ n66)  &  n91 ) ;
 assign o_41_ = ( (~ n88) ) ;
 assign o_42_ = ( (~ n85) ) ;
 assign o_43_ = ( (~ n81) ) ;
 assign o_44_ = ( (~ n74) ) ;
 assign o_45_ = ( (~ n68) ) ;
 assign o_46_ = ( (~ n60) ) ;
 assign o_47_ = ( i_17_  &  (~ i_35_)  &  (~ n46)  &  (~ n76) ) ;
 assign o_48_ = ( (~ n49) ) ;
 assign o_49_ = ( (~ n44) ) ;
 assign o_50_ = ( i_57_  &  (~ n66)  &  (~ n229) ) ;
 assign o_51_ = ( i_48_  &  (~ i_49_)  &  (~ i_50_)  &  (~ n55)  &  (~ n228) ) ;
 assign o_52_ = ( (~ n30) ) ;
 assign o_53_ = ( i_63_  &  (~ i_64_)  &  (~ n223)  &  (~ n229) ) ;
 assign o_54_ = ( i_55_  &  (~ i_62_)  &  n26  &  (~ n214) ) ;
 assign o_55_ = ( i_35_  &  (~ i_62_)  &  (~ n214)  &  (~ n227) ) ;
 assign o_56_ = ( (~ n19) ) ;
 assign o_57_ = ( i_18_  &  n13  &  n18  &  (~ n221) ) ;
 assign o_58_ = ( i_22_  &  n6  &  n13  &  n14  &  n16  &  (~ n193) ) ;
 assign o_59_ = ( i_40_  &  n12 ) ;
 assign o_60_ = ( i_7_  &  (~ n149) ) ;
 assign o_61_ = ( i_8_  &  n10 ) ;
 assign o_62_ = ( i_47_  &  n6  &  n8  &  (~ n180) ) ;
 assign o_63_ = ( i_56_  &  n6  &  n5  &  n7 ) ;
 assign o_64_ = ( n4  &  n5  &  i_30_ ) ;
 assign n4 = ( n7  &  n185  &  (~ n205) ) ;
 assign n5 = ( n132  &  (~ n208) ) ;
 assign n6 = ( n185  &  (~ n186) ) ;
 assign n7 = ( (~ i_50_)  &  (~ i_58_)  &  (~ i_60_)  &  (~ n180) ) ;
 assign n8 = ( (~ i_60_)  &  n5  &  (~ n99) ) ;
 assign n10 = ( (~ i_40_)  &  n8  &  (~ n71)  &  (~ n205)  &  (~ n212) ) ;
 assign n12 = ( (~ i_50_)  &  n154 ) ;
 assign n13 = ( (~ i_15_)  &  (~ i_41_)  &  (~ i_62_)  &  (~ n197) ) ;
 assign n14 = ( (~ i_3_)  &  (~ n208) ) ;
 assign n16 = ( (~ i_60_)  &  (~ n71)  &  (~ n99) ) ;
 assign n18 = ( n110  &  (~ n212)  &  (~ n219) ) ;
 assign n20 = ( i_36_ ) | ( n170 ) | ( n224 ) ;
 assign n22 = ( n222 ) | ( n135 ) | ( n77 ) ;
 assign n19 = ( i_16_ ) | ( (~ i_20_) ) | ( i_21_ ) | ( n20 ) | ( n22 ) ;
 assign n26 = ( (~ i_35_)  &  (~ n227) ) ;
 assign n31 = ( i_45_ ) | ( n180 ) ;
 assign n32 = ( i_47_ ) | ( i_48_ ) | ( i_49_ ) ;
 assign n33 = ( i_33_ ) | ( n72 ) | ( n70 ) | ( i_31_ ) | ( i_17_ ) | ( i_34_ ) ;
 assign n35 = ( i_15_ ) | ( n222 ) ;
 assign n36 = ( i_5_ ) | ( n65 ) | ( i_2_ ) | ( i_1_ ) ;
 assign n37 = ( i_9_ ) | ( n61 ) ;
 assign n38 = ( i_14_ ) | ( i_50_ ) | ( n190 ) ;
 assign n30 = ( (~ i_12_) ) | ( n31 ) | ( n32 ) | ( n33 ) | ( n35 ) | ( n36 ) | ( n37 ) | ( n38 ) ;
 assign n45 = ( n52 ) | ( n89 ) | ( n54 ) ;
 assign n46 = ( i_42_ ) | ( n180 ) | ( n179 ) ;
 assign n48 = ( i_59_ ) | ( n98 ) | ( n203 ) ;
 assign n44 = ( (~ i_53_) ) | ( i_54_ ) | ( i_55_ ) | ( n45 ) | ( n46 ) | ( n48 ) ;
 assign n50 = ( i_51_ ) | ( n202 ) ;
 assign n51 = ( n78 ) | ( (~ n185) ) ;
 assign n52 = ( i_35_ ) | ( i_34_ ) | ( i_33_ ) ;
 assign n53 = ( i_41_ ) | ( n175 ) ;
 assign n54 = ( n65 ) | ( n37 ) | ( n64 ) ;
 assign n55 = ( i_62_ ) | ( (~ n108) ) | ( n204 ) ;
 assign n49 = ( (~ i_31_) ) | ( n50 ) | ( n51 ) | ( n52 ) | ( n53 ) | ( n54 ) | ( n55 ) ;
 assign n61 = ( i_11_ ) | ( i_10_ ) ;
 assign n64 = ( n198 ) | ( n104 ) | ( i_17_ ) | ( n106 ) ;
 assign n65 = ( n196 ) | ( n197 ) ;
 assign n66 = ( i_56_ ) | ( i_55_ ) ;
 assign n67 = ( i_51_ ) | ( i_35_ ) | ( n53 ) ;
 assign n60 = ( (~ i_9_) ) | ( n51 ) | ( n61 ) | ( n64 ) | ( n65 ) | ( n66 ) | ( n67 ) | ( (~ n91) ) ;
 assign n70 = ( i_35_ ) | ( n163 ) ;
 assign n71 = ( i_47_ ) | ( n180 ) ;
 assign n72 = ( i_40_ ) | ( i_42_ ) | ( i_41_ ) ;
 assign n73 = ( i_51_ ) | ( i_50_ ) ;
 assign n68 = ( (~ i_34_) ) | ( i_55_ ) | ( n48 ) | ( n54 ) | ( n70 ) | ( n71 ) | ( n72 ) | ( n73 ) ;
 assign n76 = ( n65 ) | ( n208 ) | ( i_15_ ) | ( i_30_ ) | ( n55 ) | ( n89 ) | ( n125 ) ;
 assign n77 = ( i_45_ ) | ( n175 ) ;
 assign n78 = ( i_50_ ) | ( n184 ) ;
 assign n79 = ( i_31_ ) | ( n52 ) ;
 assign n80 = ( i_9_ ) | ( i_17_ ) ;
 assign n74 = ( (~ i_2_) ) | ( i_5_ ) | ( n50 ) | ( n76 ) | ( n77 ) | ( n78 ) | ( n79 ) | ( n80 ) ;
 assign n82 = ( n53 ) | ( n174 ) | ( (~ n185) ) ;
 assign n83 = ( i_53_ ) | ( n73 ) | ( (~ n91) ) | ( n189 ) ;
 assign n81 = ( (~ i_1_) ) | ( i_2_ ) | ( i_5_ ) | ( n54 ) | ( n79 ) | ( n82 ) | ( n83 ) ;
 assign n86 = ( n36 ) | ( n64 ) | ( n79 ) | ( n37 ) ;
 assign n87 = ( i_55_ ) | ( n202 ) ;
 assign n85 = ( (~ i_49_) ) | ( n48 ) | ( n73 ) | ( n82 ) | ( n86 ) | ( n87 ) ;
 assign n89 = ( i_37_ ) | ( n224 ) ;
 assign n88 = ( (~ i_33_) ) | ( i_34_ ) | ( i_35_ ) | ( n46 ) | ( n54 ) | ( n55 ) | ( n89 ) ;
 assign n91 = ( (~ i_58_)  &  (~ i_59_)  &  (~ i_60_)  &  (~ n187) ) ;
 assign n98 = ( i_60_ ) | ( n187 ) ;
 assign n99 = ( i_50_ ) | ( n203 ) ;
 assign n101 = ( n71 ) | ( n231 ) | ( n196 ) | ( n208 ) ;
 assign n97 = ( (~ i_59_) ) | ( n72 ) | ( n98 ) | ( n99 ) | ( n101 ) ;
 assign n104 = ( n225 ) | ( n143 ) ;
 assign n105 = ( i_16_ ) | ( n199 ) | ( n36 ) | ( i_20_ ) | ( i_21_ ) | ( i_13_ ) ;
 assign n106 = ( (~ i_29_) ) | ( i_30_ ) ;
 assign n102 = ( (~ i_19_) ) | ( i_32_ ) | ( n20 ) | ( n77 ) | ( n79 ) | ( n104 ) | ( n105 ) | ( n106 ) ;
 assign n108 = ( (~ i_58_)  &  (~ n66) ) ;
 assign n110 = ( (~ i_40_)  &  (~ i_43_)  &  n14  &  (~ n78)  &  (~ n214) ) ;
 assign n112 = ( (~ i_43_)  &  n129 ) ;
 assign n117 = ( n82 ) | ( n135 ) | ( n125 ) | ( i_30_ ) | ( i_36_ ) | ( n191 ) ;
 assign n118 = ( (~ n91) ) | ( n188 ) | ( n223 ) ;
 assign n115 = ( (~ i_21_) ) | ( n50 ) | ( n117 ) | ( n118 ) ;
 assign n121 = ( (~ i_10_)  &  (~ n198) ) ;
 assign n125 = ( i_18_ ) | ( n219 ) | ( n221 ) ;
 assign n127 = ( i_36_ ) | ( n165 ) | ( n212 ) ;
 assign n124 = ( (~ i_32_) ) | ( n79 ) | ( n105 ) | ( n125 ) | ( n127 ) ;
 assign n129 = ( (~ i_37_)  &  (~ n205) ) ;
 assign n132 = ( (~ i_15_)  &  n192 ) ;
 assign n135 = ( n79 ) | ( n199 ) | ( n36 ) ;
 assign n133 = ( (~ i_16_) ) | ( i_21_ ) | ( (~ i_29_) ) | ( n104 ) | ( n127 ) | ( n135 ) ;
 assign n137 = ( i_48_ ) | ( n184 ) ;
 assign n138 = ( i_49_ ) | ( n73 ) ;
 assign n139 = ( i_57_ ) | ( i_62_ ) | ( n188 ) | ( n203 ) | ( n204 ) ;
 assign n136 = ( (~ i_36_) ) | ( n22 ) | ( n87 ) | ( n89 ) | ( n137 ) | ( n138 ) | ( n139 ) ;
 assign n142 = ( i_10_ ) | ( n197 ) | ( n215 ) ;
 assign n143 = ( i_22_ ) | ( i_18_ ) | ( i_24_ ) ;
 assign n144 = ( i_62_ ) | ( (~ n16) ) | ( n89 ) | ( n106 ) | ( n225 ) ;
 assign n141 = ( (~ i_0_) ) | ( i_3_ ) | ( n142 ) | ( n143 ) | ( n144 ) ;
 assign n149 = ( i_28_ ) | ( i_43_ ) | ( n51 ) | ( n106 ) | ( (~ n192) ) | ( n214 ) | ( n215 ) | ( n216 ) ;
 assign n148 = ( i_7_ ) | ( (~ i_62_) ) | ( n149 ) ;
 assign n151 = ( (~ i_62_)  &  (~ n195) ) ;
 assign n154 = ( (~ i_58_)  &  n112  &  n121 ) ;
 assign n160 = ( n164 ) | ( n191 ) | ( i_52_ ) | ( n190 ) ;
 assign n161 = ( i_19_ ) | ( n105 ) | ( n200 ) ;
 assign n158 = ( (~ i_23_) ) | ( n82 ) | ( n160 ) | ( n161 ) ;
 assign n163 = ( i_37_ ) | ( i_39_ ) ;
 assign n164 = ( n79 ) | ( n186 ) | ( i_32_ ) | ( i_36_ ) ;
 assign n165 = ( n139 ) | ( n87 ) | ( i_52_ ) | ( n73 ) | ( n32 ) | ( n31 ) | ( n72 ) ;
 assign n167 = ( i_23_ ) | ( n161 ) ;
 assign n162 = ( (~ i_38_) ) | ( n163 ) | ( n164 ) | ( n165 ) | ( n167 ) ;
 assign n170 = ( n118 ) | ( n138 ) | ( n137 ) | ( i_37_ ) | ( i_52_ ) | ( n202 ) ;
 assign n171 = ( i_38_ ) | ( i_39_ ) ;
 assign n168 = ( i_43_ ) | ( (~ i_44_) ) | ( i_45_ ) | ( n72 ) | ( n164 ) | ( n167 ) | ( n170 ) | ( n171 ) ;
 assign n174 = ( i_45_ ) | ( n184 ) ;
 assign n175 = ( i_42_ ) | ( i_43_ ) ;
 assign n172 = ( (~ i_27_) ) | ( i_38_ ) | ( i_44_ ) | ( n89 ) | ( n160 ) | ( n167 ) | ( n174 ) | ( n175 ) ;
 assign n179 = ( i_47_ ) | ( n73 ) ;
 assign n180 = ( i_46_ ) | ( i_43_ ) ;
 assign n181 = ( i_9_ ) | ( n196 ) | ( n222 ) | ( n142 ) | ( n33 ) ;
 assign n178 = ( i_5_ ) | ( (~ i_45_) ) | ( n48 ) | ( n87 ) | ( n179 ) | ( n180 ) | ( n181 ) ;
 assign n183 = ( i_40_ ) | ( i_39_ ) ;
 assign n184 = ( i_47_ ) | ( i_46_ ) ;
 assign n185 = ( (~ i_37_)  &  (~ n183) ) ;
 assign n186 = ( i_28_ ) | ( n106 ) ;
 assign n187 = ( i_61_ ) | ( i_62_ ) ;
 assign n188 = ( i_63_ ) | ( i_64_ ) ;
 assign n189 = ( i_54_ ) | ( n66 ) ;
 assign n190 = ( n98 ) | ( n189 ) | ( i_51_ ) | ( n188 ) | ( i_59_ ) | ( i_58_ ) | ( i_57_ ) | ( i_53_ ) ;
 assign n191 = ( i_48_ ) | ( i_49_ ) | ( i_50_ ) ;
 assign n192 = ( (~ i_24_)  &  (~ i_25_) ) ;
 assign n193 = ( i_26_ ) | ( (~ n192) ) ;
 assign n195 = ( i_8_ ) | ( i_7_ ) ;
 assign n196 = ( i_4_ ) | ( i_0_ ) | ( i_3_ ) ;
 assign n197 = ( i_6_ ) | ( n195 ) ;
 assign n198 = ( i_15_ ) | ( i_14_ ) ;
 assign n199 = ( n198 ) | ( n37 ) | ( i_12_ ) | ( i_17_ ) ;
 assign n200 = ( i_22_ ) | ( i_18_ ) | ( n193 ) ;
 assign n202 = ( i_53_ ) | ( i_54_ ) ;
 assign n203 = ( i_56_ ) | ( i_58_ ) ;
 assign n204 = ( i_59_ ) | ( i_61_ ) | ( i_60_ ) ;
 assign n205 = ( i_28_ ) | ( (~ i_29_) ) ;
 assign n208 = ( i_14_ ) | ( n61 ) ;
 assign n212 = ( i_30_ ) | ( n163 ) ;
 assign n214 = ( i_60_ ) | ( n203 ) ;
 assign n215 = ( i_11_ ) | ( n198 ) ;
 assign n216 = ( i_8_ ) | ( i_10_ ) ;
 assign n219 = ( i_26_ ) | ( n205 ) ;
 assign n221 = ( i_22_ ) | ( (~ n192) ) ;
 assign n222 = ( n186 ) | ( n200 ) ;
 assign n223 = ( i_57_ ) | ( n66 ) ;
 assign n224 = ( i_41_ ) | ( n183 ) ;
 assign n225 = ( i_25_ ) | ( i_26_ ) | ( i_28_ ) ;
 assign n226 = ( i_0_ ) | ( i_3_ ) | ( n142 ) ;
 assign n227 = ( i_41_ ) | ( n104 ) | ( n106 ) | ( n179 ) | ( n180 ) | ( (~ n185) ) | ( n226 ) ;
 assign n228 = ( n82 ) | ( n86 ) | ( n50 ) ;
 assign n229 = ( (~ n91) ) | ( n191 ) | ( n228 ) ;
 assign n231 = ( i_55_ ) | ( i_51_ ) | ( n197 ) | ( n70 ) | ( n35 ) ;
 assign n232 = ( i_21_ ) | ( n190 ) | ( n117 ) ;
 assign o_5_ = ( i_29_ ) ;


endmodule

