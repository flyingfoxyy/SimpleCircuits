module misex3_mapped (
	a, b, c, d, e, f, g, h, 
	i, j, k, l, m, n, r2, s2, p2, q2, 
	t2, u2, j2, k2, h2, i2, n2, o2, l2, m2);

input a, b, c, d, e, f, g, h, i, j, k, l, m, n;

output r2, s2, p2, q2, t2, u2, j2, k2, h2, i2, n2, o2, l2, m2;

wire wire5098, wire5099, wire5139, wire5175, n_n1344, wire5264, wire5265, wire5268, wire5305, wire5306, wire5307, wire5333, wire5399, wire5400, wire5448, wire5449, n_n1425, wire5521, n_n1495, wire5619, wire5649, wire5650, wire5654, n_n2493, wire753, wire5668, wire5672, n_n1874, wire5722, wire5726, wire5809, wire5810, wire5811, n_n1573, wire5828, wire5829, wire5873, wire5936, wire5937, wire5938, wire6303, wire6304, wire6306, n_n1939, wire6322, wire6323, n_n1089, n_n842, n_n840, n_n1161, n_n1207, n_n711, n_n713, n_n709, n_n1188, n_n886, n_n920, wire38, n_n942, wire20, wire46, n_n893, wire75, wire84, wire148, n_n1261, wire1145, wire153, wire172, wire175, wire202, wire224, wire229, wire233, wire393, n_n1177, n_n1165, n_n904, n_n626, n_n671, n_n1101, n_n1229, n_n1193, wire5207, wire5208, wire5209, wire5210, wire22, wire31, wire58, wire45, wire54, wire71, wire65, wire101, wire113, n_n1228, n_n766, wire138, wire195, wire232, wire258, wire371, n_n1217, n_n1201, n_n1220, n_n918, wire15, wire41, wire1012, wire29, n_n1104, wire98, wire228, wire265, wire25, wire32, wire220, wire390, n_n861, wire417, n_n1187, n_n996, n_n1155, n_n1171, n_n698, n_n617, n_n730, n_n618, n_n857, n_n933, n_n821, n_n700, n_n824, wire928, wire929, wire5406, wire5407, n_n1792, wire30, wire34, n_n747, wire179, wire210, wire255, wire291, wire309, wire380, n_n1069, n_n1203, n_n876, n_n1166, wire871, wire5474, wire5475, wire74, wire76, n_n1233, wire5499, wire92, wire112, wire120, wire183, wire184, wire196, wire223, wire230, n_n841, n_n1194, wire5583, wire5584, wire5585, wire33, wire93, n_n971, wire106, wire156, wire203, n_n1195, wire219, n_n1138, n_n1159, wire283, n_n1253, n_n978, n_n1249, n_n2507, n_n1080, n_n973, wire118, wire188, n_n2494, n_n1142, n_n989, wire780, wire5639, wire116, n_n2602, wire777, wire199, wire775, wire776, n_n1190, n_n1202, n_n1039, n_n987, n_n988, n_n2511, n_n975, n_n1260, n_n992, wire765, wire5659, wire157, n_n1215, wire762, wire5629, wire5633, wire267, n_n949, n_n761, n_n1231, n_n997, wire751, wire5685, wire5686, wire5687, wire190, wire44, wire57, n_n1219, n_n822, wire94, n_n1083, n_n912, wire108, n_n825, wire200, wire254, wire379, n_n1082, wire407, n_n864, wire413, n_n872, n_n838, n_n977, n_n1252, wire5731, wire5732, n_n1920, wire700, wire703, wire5740, wire5743, n_n1919, n_n1210, wire5774, wire5775, wire39, wire77, wire89, n_n1036, n_n1056, n_n823, wire117, n_n1137, n_n817, wire135, wire159, wire5751, wire160, wire164, wire165, wire5752, wire5753, wire167, wire386, n_n1022, wire5848, wire5849, wire5850, wire5851, n_n820, n_n1264, n_n3060, wire14, wire40, wire146, wire208, n_n859, wire80, wire351, n_n1085, n_n1053, n_n619, wire5905, wire5906, n_n816, wire21, wire36, wire50, wire207, n_n623, wire209, wire290, wire70, wire5814, wire320, wire6168, wire6169, wire6170, wire6171, n_n2023, wire114, wire127, wire263, wire268, wire404, n_n1204, n_n1072, n_n1028, wire37, wire384, n_n1160, n_n662, wire282, wire373, n_n1180, n_n1196, wire204, wire227, n_n1121, n_n1164, n_n1222, n_n1095, wire221, wire234, wire285, wire286, wire301, n_n1148, n_n1191, n_n1133, n_n819, n_n1131, wire79, wire158, wire170, wire194, n_n1243, n_n1227, n_n1091, wire95, wire226, wire395, n_n818, n_n529, n_n670, wire23, wire59, wire96, wire134, wire398, n_n387, n_n694, wire72, wire47, wire211, wire231, wire137, n_n1118, n_n1216, n_n868, n_n1094, wire249, n_n628, wire396, n_n1146, wire121, n_n1116, n_n940, n_n765, wire248, wire55, wire149, wire18, n_n874, n_n605, n_n1084, n_n875, n_n871, n_n235, n_n2572, wire5830, n_n2953, n_n1167, n_n1189, n_n703, wire197, wire161, wire305, wire399, wire414, wire369, n_n2660, n_n982, n_n919, n_n844, wire35, wire6251, wire6252, wire6256, wire56, wire142, wire216, wire260, wire181, wire104, wire293, wire43, wire24, wire49, wire109, wire206, wire105, wire152, wire299, wire388, wire162, wire198, wire377, wire385, wire16, wire60, wire69, wire81, wire85, wire115, wire368, wire6310, wire42, wire61, wire63, wire66, wire6287, wire140, wire6289, wire150, wire163, wire173, wire177, wire178, wire180, wire6257, wire6258, wire252, wire6262, wire6263, wire253, wire6264, wire269, wire6266, wire271, wire6268, wire272, wire274, wire276, wire6272, wire278, wire280, wire281, wire6211, wire6216, wire6217, wire307, wire6225, wire6226, wire6227, wire316, wire6230, wire317, wire6233, wire318, wire6236, wire322, wire328, wire330, wire6177, wire333, wire6180, wire334, wire6185, wire336, wire6187, wire6188, wire337, wire338, wire339, wire340, wire341, wire342, wire6151, wire352, wire353, wire354, wire355, wire357, wire362, wire389, wire6109, wire429, wire6112, wire430, wire431, wire6115, wire432, wire6118, wire433, wire6119, wire434, wire435, wire440, wire441, wire442, wire6072, wire443, wire444, wire445, wire6078, wire446, wire447, wire6082, wire448, wire449, wire6085, wire450, wire451, wire452, wire453, wire454, wire455, wire456, wire457, wire458, wire459, wire460, wire6042, wire461, wire6047, wire463, wire465, wire466, wire467, wire6054, wire469, wire6005, wire480, wire6006, wire481, wire482, wire6010, wire483, wire6012, wire484, wire6014, wire485, wire486, wire487, wire6020, wire488, wire6022, wire489, wire490, wire491, wire492, wire493, wire494, wire495, wire496, wire5971, wire499, wire500, wire501, wire5979, wire504, wire505, wire508, wire509, wire510, wire512, wire513, wire516, wire520, wire5958, wire521, wire5959, wire522, wire523, wire5964, wire527, wire5941, wire528, wire5946, wire532, wire533, wire534, wire535, wire536, wire537, wire539, wire540, wire541, wire542, wire543, wire544, wire545, wire546, wire547, wire548, wire549, wire550, wire551, wire552, wire554, wire565, wire566, wire567, wire568, wire569, wire5884, wire570, wire571, wire5886, wire572, wire573, wire575, wire576, wire577, wire5813, wire580, wire1016, wire583, wire585, wire586, wire587, wire5857, wire588, wire590, wire593, wire594, wire598, wire610, wire5839, wire611, wire617, wire618, wire619, wire626, wire627, wire628, wire629, wire630, wire631, wire632, wire633, wire635, wire643, wire644, wire5781, wire645, wire646, wire647, wire649, wire650, wire651, wire652, wire653, wire5694, wire655, wire743, wire1116, wire663, wire664, wire670, wire671, wire672, wire679, wire680, wire681, wire682, wire683, wire684, wire699, wire701, wire702, wire704, wire708, wire709, wire1112, wire1113, wire5690, wire713, wire716, wire5699, wire718, wire719, wire724, wire1068, wire5253, wire725, wire726, wire727, wire729, wire731, wire732, wire736, wire739, wire5674, wire745, wire749, wire750, wire5663, wire5664, wire754, wire766, wire767, wire5640, wire781, wire782, wire5587, wire783, wire5590, wire784, wire5592, wire785, wire786, wire787, wire5598, wire788, wire789, wire5600, wire790, wire5601, wire791, wire796, wire797, wire5557, wire798, wire799, wire802, wire5526, wire808, wire5529, wire809, wire5532, wire810, wire5534, wire811, wire812, wire813, wire814, wire815, wire816, wire817, wire818, wire821, wire822, wire823, wire826, wire827, wire828, wire829, wire830, wire831, wire832, wire833, wire834, wire835, wire836, wire837, wire5480, wire843, wire5486, wire845, wire849, wire5498, wire850, wire853, wire854, wire858, wire859, wire869, wire5454, wire879, wire880, wire884, wire886, wire895, wire898, wire900, wire901, wire902, wire5422, wire903, wire904, wire906, wire907, wire908, wire909, wire911, wire912, wire914, wire923, wire924, wire925, wire926, wire5313, wire931, wire5367, wire932, wire934, wire935, wire938, wire939, wire940, wire941, wire942, wire943, wire945, wire948, wire952, wire960, wire961, wire962, wire965, wire966, wire967, wire968, wire969, wire970, wire971, wire972, wire973, wire974, wire975, wire976, wire977, wire978, wire5309, wire982, wire983, wire985, wire5314, wire986, wire5317, wire989, wire5318, wire990, wire991, wire992, wire993, wire994, wire995, wire5289, wire997, wire1039, wire5270, wire5271, wire1018, wire5274, wire1019, wire5277, wire1020, wire5279, wire1021, wire1022, wire1023, wire1024, wire1027, wire1030, wire1031, wire1032, wire1033, wire1034, wire1036, wire5246, wire1051, wire1052, wire1053, wire1054, wire5220, wire1055, wire1057, wire1058, wire1059, wire5088, wire1060, wire1061, wire5252, wire1062, wire5213, wire1070, wire1071, wire1074, wire1075, wire1076, wire1077, wire1078, wire1079, wire1080, wire1081, wire1082, wire1083, wire1096, wire1100, wire1102, wire1106, wire5140, wire1123, wire5144, wire1147, wire1148, wire1128, wire1129, wire1130, wire1131, wire1135, wire1137, wire1198, wire1200, wire1138, wire1139, wire5116, wire1140, wire1155, wire1156, wire1157, wire1158, wire1162, wire1163, wire1166, wire1167, wire1168, wire1169, wire1170, wire1171, wire1172, wire1173, wire1175, wire1176, wire1185, wire1186, wire1187, wire1188, wire1189, wire1192, wire1193, wire1194, wire1195, wire1196, wire1197, wire5091, wire5093, wire5094, wire5095, wire5108, wire5117, wire5120, wire5125, wire5126, wire5127, wire5128, wire5129, wire5130, wire5136, wire5137, wire5146, wire5156, wire5159, wire5160, wire5161, wire5162, wire5163, wire5169, wire5170, wire5171, wire5172, wire5176, wire5177, wire5179, wire5181, wire5183, wire5184, wire5187, wire5188, wire5190, wire5191, wire5192, wire5194, wire5197, wire5198, wire5199, wire5201, wire5204, wire5205, wire5215, wire5216, wire5226, wire5227, wire5228, wire5232, wire5233, wire5237, wire5238, wire5241, wire5243, wire5244, wire5251, wire5255, wire5256, wire5257, wire5266, wire5290, wire5291, wire5293, wire5297, wire5298, wire5299, wire5300, wire5316, wire5321, wire5323, wire5325, wire5327, wire5328, wire5329, wire5330, wire5356, wire5357, wire5358, wire5359, wire5360, wire5364, wire5368, wire5379, wire5382, wire5386, wire5387, wire5388, wire5389, wire5391, wire5395, wire5396, wire5397, wire5413, wire5414, wire5415, wire5416, wire5418, wire5424, wire5431, wire5432, wire5433, wire5435, wire5436, wire5437, wire5443, wire5444, wire5446, wire5451, wire5453, wire5456, wire5457, wire5459, wire5460, wire5461, wire5462, wire5463, wire5467, wire5469, wire5477, wire5479, wire5485, wire5489, wire5490, wire5493, wire5495, wire5505, wire5507, wire5508, wire5509, wire5513, wire5515, wire5517, wire5520, wire5561, wire5570, wire5572, wire5573, wire5574, wire5575, wire5576, wire5578, wire5579, wire5602, wire5603, wire5605, wire5611, wire5613, wire5615, wire5618, wire5621, wire5637, wire5652, wire5677, wire5678, wire5679, wire5681, wire5693, wire5695, wire5703, wire5704, wire5705, wire5708, wire5709, wire5710, wire5711, wire5715, wire5718, wire5719, wire5720, wire5721, wire5727, wire5744, wire5758, wire5759, wire5760, wire5761, wire5762, wire5763, wire5766, wire5792, wire5793, wire5795, wire5797, wire5798, wire5806, wire5824, wire5825, wire5826, wire5831, wire5833, wire5835, wire5836, wire5837, wire5842, wire5846, wire5847, wire5858, wire5860, wire5864, wire5865, wire5866, wire5867, wire5870, wire5871, wire5875, wire5876, wire5877, wire5888, wire5897, wire5898, wire5899, wire5901, wire5925, wire5927, wire5928, wire5929, wire5930, wire5934, wire5943, wire5944, wire5945, wire5951, wire5954, wire5955, wire5961, wire5962, wire5963, wire5967, wire5969, wire5970, wire5981, wire5982, wire5986, wire5990, wire5998, wire5999, wire6035, wire6036, wire6037, wire6038, wire6041, wire6045, wire6057, wire6062, wire6064, wire6065, wire6066, wire6067, wire6070, wire6071, wire6100, wire6101, wire6102, wire6103, wire6106, wire6123, wire6125, wire6132, wire6133, wire6135, wire6138, wire6139, wire6141, wire6142, wire6143, wire6144, wire6145, wire6147, wire6156, wire6158, wire6159, wire6160, wire6161, wire6165, wire6176, wire6183, wire6184, wire6194, wire6195, wire6200, wire6203, wire6204, wire6205, wire6206, wire6207, wire6210, wire6213, wire6220, wire6222, wire6224, wire6238, wire6239, wire6240, wire6241, wire6245, wire6246, wire6248, wire6249, wire6250, wire6281, wire6282, wire6283, wire6285, wire6286, wire6290, wire6292, wire6298, wire6300, wire6301, wire6307, wire6309, wire6317, wire6318, _36, _37, _38, _70, _119, _120, _122, _126, _182, _183, _202, _203, _217, _218, _224, _225, _226, _227, _255, _256, _274, _275, _294, _298, _300, _313, _314, _331, _333, _334, _335, _336, _373, _378, _379, _405, _446, _493, _494, _497, _507, _508, _513, _559, _560, _561, _566, _576, _577, _589, _594, _595, _611, _612, _621, _624, _665, _666, _670, _679, _680, _763, _803, _804, _814, _843, _860, _861, _877, _905, _7270, _7308, _7373, _7387, _7390, _7433, _7437, _7453, _7462, _7467, _7479, _7481, _7503, _7511, _7524, _7528, _7541, _7556, _7569, _7632, _7649, _7662, _7671, _7743, _7745, _7751, _7757, _7759, _7776, _7780, _7783, _7794, _7798, _7815, _7833, _7862, _7877, _7920, _7925, _7927, _8063, _8076, _8084, _8097, _8115, _8116, _8202, _8227, _8242, _8243, _8290, _8318, _8344, _8362, _8370, _8385, _8388, _8391, _8394, _8427, _8439, _8469, _8474, _8487, _8504, _8515, _8524, _8533, _8543, _8553, _8574, _8577, _8608, _8619, _8636, _8639, _8646, _8668, _8701, _8711, _8715, _8731, _8732, _8742, _8746, _8747, _8748, _8750, _8769, _8771, _8772, _8776, _8786, _8794, _8801, _8819, _8820, _8823, _8830, _8835, _8851, _8855, _8868, _8878, _8880, _8882, _8890, _8939, _8940, _8970, _8976, _8993, _8998, _9007, _9018, _9020, _9021, _9051, _9054, _9055, _9062, _9064, _9065, _9067, _9075, _9076, _9092, _9094, _9128, _9142, _9143, _9161, _9163, _9164, _9184, _9185, _9186, _9190, _9192, _9203, _9209;

assign r2 = ( wire5098 ) | ( wire5099 ) | ( wire5139 ) | ( wire5175 ) ;
 assign s2 = ( n_n1344 ) | ( wire5264 ) | ( wire5265 ) | ( wire5268 ) ;
 assign p2 = ( wire5305 ) | ( wire5306 ) | ( wire5307 ) | ( wire5333 ) ;
 assign q2 = ( wire5399 ) | ( wire5400 ) | ( wire5448 ) | ( wire5449 ) ;
 assign t2 = ( wire5521 ) | ( wire5520 ) | ( _8115 ) | ( _8116 ) ;
 assign u2 = ( n_n1495 ) | ( wire5621 ) | ( _8242 ) | ( _8243 ) ;
 assign j2 = ( wire5649 ) | ( wire5650 ) | ( wire5654 ) ;
 assign k2 = ( n_n2493 ) | ( wire753 ) | ( wire5668 ) | ( wire5672 ) ;
 assign h2 = ( n_n1874 ) | ( wire5722 ) | ( wire5726 ) ;
 assign i2 = ( wire5809 ) | ( wire5810 ) | ( wire5811 ) ;
 assign n2 = ( n_n1573 ) | ( wire5828 ) | ( wire5829 ) | ( wire5873 ) ;
 assign o2 = ( wire5936 ) | ( wire5937 ) | ( _8715 ) ;
 assign l2 = ( wire6303 ) | ( wire6304 ) | ( wire6306 ) ;
 assign m2 = ( n_n1939 ) | ( wire6322 ) | ( wire6323 ) ;
 assign wire5098 = ( wire1195 ) | ( wire1197 ) | ( wire5093 ) ;
 assign wire5099 = ( wire1196 ) | ( wire5094 ) | ( wire5095 ) ;
 assign wire5139 = ( wire5129 ) | ( wire5130 ) | ( wire5136 ) | ( wire5137 ) ;
 assign wire5175 = ( wire5169 ) | ( wire5170 ) | ( wire5171 ) | ( wire5172 ) ;
 assign n_n1344 = ( wire5207 ) | ( wire5208 ) | ( wire5209 ) | ( wire5210 ) ;
 assign wire5264 = ( wire1051 ) | ( wire1052 ) | ( wire1053 ) | ( wire1054 ) ;
 assign wire5265 = ( wire1057 ) | ( wire1058 ) | ( wire1060 ) | ( wire1061 ) ;
 assign wire5268 = ( wire5232 ) | ( wire5233 ) | ( wire5266 ) ;
 assign wire5305 = ( wire1018 ) | ( wire1027 ) | ( wire5290 ) | ( wire5297 ) ;
 assign wire5306 = ( wire1031 ) | ( wire1032 ) | ( wire1036 ) ;
 assign wire5307 = ( wire1034 ) | ( wire5298 ) | ( wire5299 ) | ( wire5300 ) ;
 assign wire5333 = ( wire5327 ) | ( wire5328 ) | ( wire5329 ) | ( wire5330 ) ;
 assign wire5399 = ( wire977 ) | ( wire5360 ) | ( wire5364 ) | ( wire5396 ) ;
 assign wire5400 = ( wire5389 ) | ( wire5395 ) | ( wire5397 ) | ( _7877 ) ;
 assign wire5448 = ( wire5446 ) | ( _576 ) | ( _577 ) | ( _7920 ) ;
 assign wire5449 = ( n_n1792 ) | ( wire5443 ) | ( wire5444 ) ;
 assign n_n1425 = ( wire871 ) | ( wire5474 ) | ( wire5475 ) ;
 assign wire5521 = ( wire5462 ) | ( wire5463 ) | ( wire5467 ) | ( wire5517 ) ;
 assign n_n1495 = ( wire5583 ) | ( wire5584 ) | ( wire5585 ) ;
 assign wire5619 = ( wire783 ) | ( wire785 ) | ( wire798 ) | ( wire799 ) ;
 assign wire5649 = ( n_n2494 ) | ( n_n1215  &  wire5629  &  wire5633 ) ;
 assign wire5650 = ( wire767 ) | ( wire781 ) | ( wire782 ) ;
 assign wire5654 = ( wire116 ) | ( n_n2602 ) | ( wire777 ) | ( wire5652 ) ;
 assign n_n2493 = ( n_n1104  &  (~ wire118)  &  wire188  &  n_n975 ) ;
 assign wire753 = ( n_n1039  &  wire5663  &  wire5664 ) ;
 assign wire5668 = ( wire754 ) | ( wire781 ) | ( wire782 ) ;
 assign wire5672 = ( wire157 ) | ( wire267 ) | ( _8318 ) ;
 assign n_n1874 = ( wire751 ) | ( wire5685 ) | ( wire5686 ) | ( wire5687 ) ;
 assign wire5722 = ( wire729 ) | ( wire731 ) | ( wire732 ) | ( wire5710 ) ;
 assign wire5726 = ( wire5718 ) | ( wire5719 ) | ( wire5720 ) | ( wire5721 ) ;
 assign wire5809 = ( n_n1919 ) | ( wire5761 ) | ( wire5762 ) | ( wire5766 ) ;
 assign wire5810 = ( n_n1939 ) | ( wire5792 ) | ( wire5793 ) | ( wire5806 ) ;
 assign wire5811 = ( n_n1920 ) | ( wire5797 ) | ( wire5798 ) | ( _8524 ) ;
 assign n_n1573 = ( wire5848 ) | ( wire5849 ) | ( wire5850 ) | ( wire5851 ) ;
 assign wire5828 = ( wire5825 ) | ( n_n1210  &  wire211 ) ;
 assign wire5829 = ( wire320 ) | ( wire5824 ) | ( wire5826 ) ;
 assign wire5873 = ( wire351 ) | ( wire5866 ) | ( wire5870 ) | ( wire5871 ) ;
 assign wire5936 = ( wire546 ) | ( wire552 ) | ( wire5925 ) | ( wire5930 ) ;
 assign wire5937 = ( wire5927 ) | ( wire5928 ) | ( _8701 ) ;
 assign wire5938 = ( wire5929 ) | ( wire5934 ) | ( n_n1220  &  wire207 ) ;
 assign wire6303 = ( wire6101 ) | ( wire6102 ) | ( wire6106 ) | ( wire6301 ) ;
 assign wire6304 = ( n_n2023 ) | ( wire6138 ) | ( wire6139 ) | ( wire6300 ) ;
 assign wire6306 = ( wire6071 ) | ( wire6286 ) | ( _9209 ) ;
 assign n_n1939 = ( n_n2493 ) | ( n_n2511 ) | ( wire5774 ) | ( wire5775 ) ;
 assign wire6322 = ( wire116 ) | ( wire781 ) | ( wire782 ) | ( wire6318 ) ;
 assign wire6323 = ( wire199 ) | ( wire157 ) | ( wire267 ) | ( wire6317 ) ;
 assign n_n1089 = ( f  &  (~ g)  &  (~ h) ) ;
 assign n_n842 = ( b  &  (~ c)  &  d ) ;
 assign n_n840 = ( b  &  d  &  (~ e) ) ;
 assign n_n1161 = ( (~ e)  &  g  &  (~ h) ) ;
 assign n_n1207 = ( f  &  g  &  (~ h) ) ;
 assign n_n711 = ( b  &  c  &  e ) ;
 assign n_n713 = ( b  &  c  &  (~ d) ) ;
 assign n_n709 = ( b  &  (~ d)  &  e ) ;
 assign n_n1188 = ( g  &  j  &  (~ k) ) ;
 assign n_n886 = ( e  &  (~ f)  &  h ) ;
 assign n_n920 = ( a  &  b  &  (~ c) ) ;
 assign wire38 = ( m  &  (~ n)  &  n_n920 ) ;
 assign n_n942 = ( h  &  (~ j)  &  l ) ;
 assign wire20 = ( (~ h)  &  i  &  l ) | ( h  &  (~ i)  &  l ) | ( h  &  j  &  (~ l) ) ;
 assign wire46 = ( (~ g)  &  n_n942 ) | ( g  &  wire20 ) ;
 assign n_n893 = ( i  &  (~ j)  &  l ) ;
 assign wire75 = ( (~ m)  &  n  &  n_n893 ) ;
 assign wire84 = ( i  &  k  &  (~ m)  &  n ) ;
 assign wire148 = ( i  &  l  &  m  &  (~ n) ) ;
 assign n_n1261 = ( a  &  b  &  c ) ;
 assign wire1145 = ( a  &  b  &  d  &  (~ e) ) ;
 assign wire153 = ( wire1145 ) | ( (~ d)  &  e  &  n_n1261 ) ;
 assign wire172 = ( (~ i)  &  k  &  (~ m)  &  n ) ;
 assign wire175 = ( (~ e)  &  f  &  (~ g) ) | ( (~ e)  &  (~ f)  &  (~ g) ) ;
 assign wire202 = ( b  &  (~ c)  &  d ) | ( b  &  (~ d)  &  e ) ;
 assign wire224 = ( a  &  b  &  (~ c)  &  f ) ;
 assign wire229 = ( e  &  f  &  g ) | ( e  &  f  &  (~ g) ) ;
 assign wire233 = ( (~ i)  &  j  &  (~ k) ) | ( (~ i)  &  j  &  l ) | ( j  &  (~ k)  &  l ) ;
 assign wire393 = ( (~ f)  &  g  &  (~ h)  &  n_n711 ) | ( (~ f)  &  (~ g)  &  (~ h)  &  n_n711 ) ;
 assign n_n1177 = ( (~ m)  &  n ) ;
 assign n_n1165 = ( (~ m)  &  (~ n) ) ;
 assign n_n904 = ( a  &  (~ c)  &  d ) ;
 assign n_n626 = ( c  &  (~ e)  &  f ) ;
 assign n_n671 = ( (~ b)  &  c  &  f ) ;
 assign n_n1101 = ( (~ c)  &  d  &  f ) ;
 assign n_n1229 = ( c  &  d  &  e ) ;
 assign n_n1193 = ( f  &  g  &  (~ i) ) ;
 assign wire5207 = ( wire5199 ) | ( wire379  &  wire5183 ) | ( wire379  &  wire5184 ) ;
 assign wire5208 = ( wire1106 ) | ( wire5201 ) | ( wire152  &  wire299 ) ;
 assign wire5209 = ( wire5197 ) | ( wire5198 ) | ( wire5204 ) ;
 assign wire5210 = ( wire5205 ) | ( wire74  &  wire388 ) | ( wire74  &  wire5194 ) ;
 assign wire22 = ( k  &  (~ l)  &  m  &  (~ n) ) ;
 assign wire31 = ( (~ i)  &  l  &  m ) | ( j  &  (~ l)  &  m ) ;
 assign wire58 = ( (~ k)  &  l  &  m  &  (~ n) ) ;
 assign wire45 = ( (~ j)  &  wire22 ) | ( j  &  wire58 ) ;
 assign wire54 = ( (~ j)  &  l  &  m  &  (~ n) ) ;
 assign wire71 = ( (~ f)  &  h ) ;
 assign wire65 = ( (~ h)  &  i  &  k ) | ( h  &  (~ i)  &  k ) | ( h  &  (~ j)  &  k ) | ( h  &  j  &  (~ k) ) ;
 assign wire101 = ( wire65 ) | ( h  &  k  &  (~ l) ) ;
 assign wire113 = ( (~ j)  &  k  &  m  &  (~ n) ) ;
 assign n_n1228 = ( f  &  g  &  i ) ;
 assign n_n766 = ( f  &  g  &  (~ j) ) ;
 assign wire138 = ( wire22  &  n_n1228 ) | ( wire113  &  n_n1228 ) | ( wire22  &  n_n766 ) ;
 assign wire195 = ( f  &  g  &  j  &  wire58 ) ;
 assign wire232 = ( (~ c) ) | ( (~ d) ) | ( e ) | ( (~ f) ) ;
 assign wire258 = ( (~ e)  &  g  &  n_n904 ) ;
 assign wire371 = ( a  &  (~ c)  &  d  &  _7927 ) ;
 assign n_n1217 = ( i  &  j  &  k ) ;
 assign n_n1201 = ( f  &  g  &  h ) ;
 assign n_n1220 = ( k  &  m  &  (~ n) ) ;
 assign n_n918 = ( a  &  b  &  d ) ;
 assign wire15 = ( a  &  (~ b)  &  c ) | ( (~ a)  &  b  &  (~ d) ) ;
 assign wire41 = ( n_n1104  &  wire14 ) | ( n_n876  &  n_n875 ) ;
 assign wire1012 = ( f  &  g  &  (~ h)  &  wire16 ) ;
 assign wire29 = ( a  &  (~ b)  &  c ) | ( a  &  b  &  (~ c) ) | ( (~ a)  &  b  &  (~ d) ) ;
 assign n_n1104 = ( (~ f)  &  g  &  (~ h) ) ;
 assign wire98 = ( n_n1207  &  wire29 ) | ( n_n918  &  n_n1104 ) ;
 assign wire228 = ( j  &  l  &  m  &  (~ n) ) ;
 assign wire265 = ( j  &  (~ k)  &  m  &  (~ n) ) ;
 assign wire25 = ( n_n1195  &  wire14 ) | ( n_n876  &  n_n1148 ) ;
 assign wire32 = ( n_n904  &  n_n1201 ) | ( n_n1201  &  n_n730 ) | ( n_n904  &  n_n1196 ) ;
 assign wire220 = ( m  &  (~ n)  &  wire25 ) | ( m  &  (~ n)  &  wire32 ) ;
 assign wire390 = ( n_n1193  &  wire228 ) | ( n_n1193  &  wire265 ) ;
 assign n_n861 = ( (~ f)  &  g  &  (~ i) ) ;
 assign wire417 = ( wire228  &  n_n861 ) | ( wire265  &  n_n861 ) ;
 assign n_n1187 = ( m  &  (~ n) ) ;
 assign n_n996 = ( (~ j)  &  k  &  l ) ;
 assign n_n1155 = ( g  &  h  &  (~ i) ) ;
 assign n_n1171 = ( b  &  e  &  (~ f) ) ;
 assign n_n698 = ( (~ a)  &  b  &  e ) ;
 assign n_n617 = ( h  &  j  &  (~ k) ) ;
 assign n_n730 = ( a  &  d  &  (~ e) ) ;
 assign n_n618 = ( h  &  (~ j)  &  k ) ;
 assign n_n857 = ( (~ f)  &  g  &  i ) ;
 assign n_n933 = ( (~ i)  &  j  &  l ) ;
 assign n_n821 = ( (~ g)  &  h  &  (~ i) ) ;
 assign n_n700 = ( (~ c)  &  d  &  (~ e) ) ;
 assign n_n824 = ( f  &  h  &  (~ i) ) ;
 assign wire928 = ( wire106  &  wire142 ) | ( wire50  &  wire142 ) | ( wire142  &  wire5313 ) ;
 assign wire929 = ( wire54  &  wire106 ) | ( wire54  &  wire50 ) | ( wire54  &  wire5313 ) ;
 assign wire5406 = ( _566 ) | ( wire54  &  wire15  &  n_n1194 ) ;
 assign wire5407 = ( wire923 ) | ( wire924 ) | ( wire925 ) | ( wire926 ) ;
 assign n_n1792 = ( wire928 ) | ( wire929 ) | ( wire5406 ) | ( wire5407 ) ;
 assign wire30 = ( b  &  d  &  f ) | ( b  &  (~ e)  &  f ) ;
 assign wire34 = ( (~ c)  &  d  &  f ) | ( c  &  (~ d)  &  f ) | ( c  &  (~ e)  &  f ) ;
 assign n_n747 = ( i  &  j  &  l ) ;
 assign wire179 = ( n_n1228  &  n_n996 ) | ( n_n1207  &  n_n747 ) ;
 assign wire210 = ( b  &  (~ c)  &  d ) | ( b  &  c  &  (~ d) ) | ( (~ b)  &  c  &  (~ e) ) ;
 assign wire255 = ( g  &  (~ h) ) ;
 assign wire291 = ( m  &  (~ n)  &  n_n1201  &  wire15 ) ;
 assign wire309 = ( (~ f)  &  h  &  n_n709 ) ;
 assign wire380 = ( g  &  h  &  (~ i)  &  wire54 ) ;
 assign n_n1069 = ( (~ c)  &  (~ d)  &  e ) ;
 assign n_n1203 = ( c  &  e  &  (~ f) ) ;
 assign n_n876 = ( a  &  c  &  (~ d) ) ;
 assign n_n1166 = ( (~ h)  &  i  &  (~ j) ) ;
 assign wire871 = ( wire390  &  wire43 ) | ( wire43  &  wire1068 ) | ( wire43  &  wire5253 ) ;
 assign wire5474 = ( wire44  &  wire5469 ) | ( (~ n_n842)  &  wire224  &  wire44 ) ;
 assign wire5475 = ( wire869 ) | ( wire138  &  wire43 ) | ( wire195  &  wire43 ) ;
 assign wire74 = ( i  &  (~ j)  &  k ) | ( (~ i)  &  j  &  (~ k) ) | ( (~ i)  &  j  &  l ) | ( j  &  (~ k)  &  l ) | ( i  &  k  &  (~ l) ) | ( (~ j)  &  k  &  (~ l) ) ;
 assign wire76 = ( (~ j)  &  l  &  (~ m)  &  n ) ;
 assign n_n1233 = ( (~ d)  &  f  &  g ) ;
 assign wire5499 = ( (~ d)  &  f  &  (~ g) ) ;
 assign wire92 = ( wire20  &  n_n1233 ) | ( n_n942  &  wire5499 ) ;
 assign wire112 = ( f  &  g ) ;
 assign wire120 = ( a  &  m  &  (~ n) ) ;
 assign wire183 = ( i  &  (~ j)  &  k ) | ( (~ i)  &  j  &  l ) | ( j  &  (~ k)  &  l ) | ( i  &  k  &  (~ l) ) | ( (~ j)  &  k  &  (~ l) ) ;
 assign wire184 = ( g  &  n_n842  &  wire71 ) | ( g  &  n_n711  &  wire71 ) | ( (~ g)  &  n_n711  &  wire71 ) ;
 assign wire196 = ( (~ b)  &  f ) ;
 assign wire223 = ( m  &  (~ n)  &  n_n920  &  n_n1233 ) ;
 assign wire230 = ( (~ f)  &  (~ h)  &  i ) | ( g  &  (~ h)  &  i ) ;
 assign n_n841 = ( g  &  (~ h)  &  i ) ;
 assign n_n1194 = ( f  &  (~ g)  &  h ) ;
 assign wire5583 = ( wire836 ) | ( wire5578 ) | ( wire93  &  wire135 ) ;
 assign wire5584 = ( wire833 ) | ( wire834 ) | ( wire5572 ) | ( wire5579 ) ;
 assign wire5585 = ( wire5573 ) | ( wire5574 ) | ( wire5575 ) | ( wire5576 ) ;
 assign wire33 = ( wire22 ) | ( wire113 ) ;
 assign wire93 = ( (~ b)  &  c  &  (~ e) ) | ( (~ b)  &  c  &  f ) | ( b  &  e  &  (~ f) ) ;
 assign n_n971 = ( (~ f)  &  (~ g)  &  h ) ;
 assign wire106 = ( n_n920  &  n_n1194 ) | ( n_n918  &  n_n971 ) ;
 assign wire156 = ( n_n1207  &  n_n920 ) | ( n_n918  &  n_n1104 ) ;
 assign wire203 = ( n_n920  &  n_n1228 ) | ( n_n918  &  n_n857 ) ;
 assign n_n1195 = ( (~ f)  &  g  &  h ) ;
 assign wire219 = ( m  &  (~ n)  &  n_n918  &  n_n1195 ) ;
 assign n_n1138 = ( (~ c)  &  (~ d)  &  (~ f) ) ;
 assign n_n1159 = ( (~ j)  &  (~ k)  &  (~ l) ) ;
 assign wire283 = ( (~ h)  &  (~ i)  &  j ) ;
 assign n_n1253 = ( b  &  c  &  d ) ;
 assign n_n978 = ( k  &  l  &  (~ m)  &  n ) ;
 assign n_n1249 = ( (~ e)  &  (~ f)  &  g ) ;
 assign n_n2507 = ( wire283  &  n_n1253  &  n_n978  &  n_n1249 ) ;
 assign n_n1080 = ( (~ c)  &  (~ d)  &  (~ e) ) ;
 assign n_n973 = ( c  &  d  &  (~ e) ) ;
 assign wire118 = ( i ) | ( (~ j) ) ;
 assign wire188 = ( k  &  l  &  (~ m)  &  (~ n) ) ;
 assign n_n2494 = ( n_n1104  &  n_n973  &  (~ wire118)  &  wire188 ) ;
 assign n_n1142 = ( (~ g)  &  h  &  i ) ;
 assign n_n989 = ( j  &  (~ k)  &  l ) ;
 assign wire780 = ( n_n1104  &  n_n975  &  n_n1204  &  wire5640 ) ;
 assign wire5639 = ( m  &  (~ n)  &  n_n997  &  wire5637 ) ;
 assign wire116 = ( wire780 ) | ( n_n1142  &  n_n989  &  wire5639 ) ;
 assign n_n2602 = ( n_n1207  &  n_n1069  &  (~ wire118)  &  wire188 ) ;
 assign wire777 = ( n_n987  &  n_n988  &  wire398  &  n_n982 ) ;
 assign wire199 = ( n_n2602 ) | ( wire777 ) ;
 assign wire775 = ( n_n1253  &  n_n1249  &  n_n1085  &  n_n982 ) ;
 assign wire776 = ( n_n1195  &  n_n973  &  n_n1204  &  n_n1180 ) ;
 assign n_n1190 = ( (~ l)  &  (~ m)  &  (~ n) ) ;
 assign n_n1202 = ( (~ k)  &  (~ m)  &  (~ n) ) ;
 assign n_n1039 = ( (~ f)  &  (~ g)  &  (~ h) ) ;
 assign n_n987 = ( e  &  (~ f)  &  g ) ;
 assign n_n988 = ( (~ b)  &  c  &  d ) ;
 assign n_n2511 = ( wire283  &  n_n978  &  n_n987  &  n_n988 ) ;
 assign n_n975 = ( (~ c)  &  d  &  e ) ;
 assign n_n1260 = ( d  &  e  &  f ) ;
 assign n_n992 = ( g  &  h  &  i ) ;
 assign wire765 = ( n_n1253  &  n_n978  &  n_n1252  &  n_n1264 ) ;
 assign wire5659 = ( m  &  (~ n)  &  n_n1261  &  n_n1146 ) ;
 assign wire157 = ( wire765 ) | ( n_n1260  &  n_n992  &  wire5659 ) ;
 assign n_n1215 = ( l  &  m  &  (~ n) ) ;
 assign wire762 = ( n_n1229  &  n_n1217  &  n_n1201  &  n_n1204 ) ;
 assign wire5629 = ( d  &  f  &  (~ j) ) ;
 assign wire5633 = ( (~ n_n1260)  &  n_n992  &  n_n997  &  n_n1222 ) ;
 assign wire267 = ( wire762 ) | ( n_n1215  &  wire5629  &  wire5633 ) ;
 assign n_n949 = ( a  &  (~ b)  &  c ) ;
 assign n_n761 = ( a  &  c  &  e ) ;
 assign n_n1231 = ( (~ e)  &  f  &  g ) ;
 assign n_n997 = ( (~ a)  &  b  &  c ) ;
 assign wire751 = ( m  &  (~ n)  &  wire92  &  n_n997 ) ;
 assign wire5685 = ( n_n2602 ) | ( wire749 ) | ( wire181  &  wire5677 ) ;
 assign wire5686 = ( wire745 ) | ( wire46  &  wire5679 ) ;
 assign wire5687 = ( wire750 ) | ( wire46  &  wire5681 ) ;
 assign wire190 = ( h  &  k  &  m  &  (~ n) ) ;
 assign wire44 = ( h  &  wire22 ) | ( (~ g)  &  wire190 ) ;
 assign wire57 = ( (~ c) ) | ( (~ d) ) ;
 assign n_n1219 = ( (~ l)  &  m  &  (~ n) ) ;
 assign n_n822 = ( f  &  h  &  k ) ;
 assign wire94 = ( n_n1220  &  n_n1194 ) | ( n_n1219  &  n_n822 ) ;
 assign n_n1083 = ( (~ e)  &  f  &  h ) ;
 assign n_n912 = ( (~ e)  &  f  &  (~ g) ) ;
 assign wire108 = ( wire22  &  n_n1083 ) | ( wire190  &  n_n912 ) ;
 assign n_n825 = ( (~ f)  &  h  &  k ) ;
 assign wire200 = ( n_n1220  &  n_n971 ) | ( n_n1219  &  n_n825 ) ;
 assign wire254 = ( (~ k)  &  (~ l)  &  (~ m)  &  (~ n) ) ;
 assign wire379 = ( g  &  (~ j)  &  wire22 ) | ( g  &  j  &  wire58 ) ;
 assign n_n1082 = ( e  &  (~ g)  &  h ) ;
 assign wire407 = ( (~ g)  &  (~ h)  &  (~ i) ) ;
 assign n_n864 = ( e  &  g  &  (~ i) ) ;
 assign wire413 = ( e  &  g  &  (~ i)  &  _8391 ) ;
 assign n_n872 = ( a  &  (~ d)  &  e ) ;
 assign n_n838 = ( b  &  d  &  f ) ;
 assign n_n977 = ( (~ i)  &  j  &  (~ k) ) ;
 assign n_n1252 = ( e  &  f  &  g ) ;
 assign wire5731 = ( wire223  &  wire149 ) | ( wire149  &  wire388 ) ;
 assign wire5732 = ( wire708 ) | ( wire709 ) | ( wire46  &  wire5727 ) ;
 assign n_n1920 = ( wire5731 ) | ( wire5732 ) | ( wire38  &  wire92 ) ;
 assign wire700 = ( wire20  &  n_n904  &  n_n1187  &  n_n1252 ) ;
 assign wire703 = ( n_n920  &  n_n1187  &  n_n1233  &  wire55 ) ;
 assign wire5740 = ( wire701 ) | ( wire702 ) | ( wire704 ) ;
 assign wire5743 = ( wire699 ) | ( wire55  &  wire388 ) | ( wire18  &  wire388 ) ;
 assign n_n1919 = ( wire700 ) | ( wire703 ) | ( wire5740 ) | ( wire5743 ) ;
 assign n_n1210 = ( k  &  (~ m)  &  n ) ;
 assign wire5774 = ( wire670 ) | ( wire671 ) | ( wire672 ) ;
 assign wire5775 = ( n_n2507 ) | ( n_n2494 ) | ( wire775 ) | ( wire776 ) ;
 assign wire39 = ( i  &  (~ j)  &  k ) | ( (~ i)  &  j  &  l ) | ( i  &  k  &  (~ l) ) | ( (~ j)  &  k  &  (~ l) ) ;
 assign wire77 = ( k  &  (~ l)  &  (~ m)  &  n ) ;
 assign wire89 = ( f  &  (~ h)  &  i ) | ( f  &  h  &  (~ i) ) | ( f  &  h  &  (~ j) ) ;
 assign n_n1036 = ( (~ k)  &  (~ m)  &  n ) ;
 assign n_n1056 = ( (~ l)  &  (~ m)  &  n ) ;
 assign n_n823 = ( f  &  h  &  j ) ;
 assign wire117 = ( n_n822  &  n_n1056 ) | ( n_n1036  &  n_n823 ) ;
 assign n_n1137 = ( g  &  h  &  j ) ;
 assign n_n817 = ( g  &  h  &  k ) ;
 assign wire135 = ( n_n1036  &  n_n1137 ) | ( n_n1056  &  n_n817 ) ;
 assign wire159 = ( n_n876  &  n_n864 ) | ( n_n861  &  n_n872 ) ;
 assign wire5751 = ( b  &  d  &  e ) ;
 assign wire160 = ( n_n1253  &  n_n1082 ) | ( n_n1195  &  wire5751 ) ;
 assign wire164 = ( g  &  (~ h)  &  i ) | ( g  &  h  &  (~ i) ) | ( g  &  h  &  (~ j) ) ;
 assign wire165 = ( i  &  (~ j)  &  k ) | ( (~ i)  &  j  &  (~ k) ) | ( (~ i)  &  j  &  l ) | ( i  &  k  &  (~ l) ) ;
 assign wire5752 = ( e  &  (~ g)  &  (~ h) ) ;
 assign wire5753 = ( b  &  d  &  e ) ;
 assign wire167 = ( n_n1253  &  wire5752 ) | ( n_n1104  &  wire5753 ) ;
 assign wire386 = ( (~ i)  &  (~ k) ) ;
 assign n_n1022 = ( f  &  h  &  (~ j) ) ;
 assign wire5848 = ( wire617 ) | ( wire5842 ) | ( _298 ) | ( _8543 ) ;
 assign wire5849 = ( wire611 ) | ( wire220  &  wire81 ) | ( wire220  &  wire5831 ) ;
 assign wire5850 = ( wire618 ) | ( _274 ) | ( _275 ) ;
 assign wire5851 = ( wire5846 ) | ( wire5847 ) ;
 assign n_n820 = ( g  &  h  &  (~ j) ) ;
 assign n_n1264 = ( h  &  i  &  j ) ;
 assign n_n3060 = ( n_n904  &  wire113  &  _8608 ) ;
 assign wire14 = ( a  &  c  &  e ) | ( a  &  (~ d)  &  e ) ;
 assign wire40 = ( h  &  (~ i)  &  k ) | ( h  &  (~ j)  &  k ) ;
 assign wire146 = ( h  &  (~ j) ) ;
 assign wire208 = ( g  &  n_n1171  &  wire146 ) | ( (~ g)  &  wire30  &  wire146 ) ;
 assign n_n859 = ( e  &  g  &  i ) ;
 assign wire80 = ( n_n857  &  wire14 ) | ( n_n1228  &  wire16 ) ;
 assign wire351 = ( wire113  &  wire80 ) | ( wire113  &  n_n876  &  n_n859 ) ;
 assign n_n1085 = ( h  &  i  &  (~ j) ) ;
 assign n_n1053 = ( (~ b)  &  c  &  (~ e) ) ;
 assign n_n619 = ( (~ h)  &  i  &  k ) ;
 assign wire5905 = ( wire570 ) | ( wire573 ) | ( wire5897 ) | ( wire5901 ) ;
 assign wire5906 = ( wire572 ) | ( wire580 ) ;
 assign n_n816 = ( (~ g)  &  h  &  k ) ;
 assign wire21 = ( (~ j)  &  k  &  (~ m) ) | ( j  &  (~ k)  &  (~ m) ) ;
 assign wire36 = ( b  &  (~ c)  &  d ) | ( b  &  c  &  (~ d) ) ;
 assign wire50 = ( n_n876  &  n_n1082 ) | ( n_n971  &  wire14 ) ;
 assign wire207 = ( wire29  &  n_n1194 ) | ( n_n918  &  n_n971 ) ;
 assign n_n623 = ( c  &  f  &  (~ g) ) ;
 assign wire209 = ( n_n1203  &  n_n1202 ) | ( n_n1202  &  n_n623 ) | ( n_n1036  &  n_n623 ) ;
 assign wire290 = ( g  &  h  &  i  &  (~ n) ) ;
 assign wire70 = ( j  &  (~ k)  &  (~ m)  &  n ) ;
 assign wire5814 = ( n_n709  &  n_n992  &  wire70 ) | ( n_n1171  &  n_n992  &  wire70 ) ;
 assign wire320 = ( wire5814 ) | ( _255 ) | ( _256 ) ;
 assign wire6168 = ( wire353 ) | ( n_n1072  &  wire161 ) ;
 assign wire6169 = ( wire352 ) | ( wire354 ) | ( wire355 ) | ( wire389 ) ;
 assign wire6170 = ( wire357 ) | ( wire6165 ) | ( n_n1028  &  _8830 ) ;
 assign wire6171 = ( wire362 ) | ( wire6159 ) | ( wire6160 ) | ( wire6161 ) ;
 assign n_n2023 = ( wire6168 ) | ( wire6169 ) | ( wire6170 ) | ( wire6171 ) ;
 assign wire114 = ( (~ g)  &  (~ h) ) ;
 assign wire127 = ( (~ i)  &  (~ m)  &  (~ n) ) ;
 assign wire263 = ( (~ b)  &  (~ m)  &  n ) ;
 assign wire268 = ( (~ c)  &  e  &  (~ f) ) | ( c  &  (~ e)  &  (~ f) ) ;
 assign wire404 = ( (~ b)  &  m  &  (~ n) ) ;
 assign n_n1204 = ( l  &  (~ m)  &  (~ n) ) ;
 assign n_n1072 = ( (~ d)  &  (~ e)  &  (~ f) ) ;
 assign n_n1028 = ( (~ e)  &  (~ f)  &  (~ g) ) ;
 assign wire37 = ( h ) | ( i ) ;
 assign wire384 = ( h  &  (~ i)  &  (~ j) ) ;
 assign n_n1160 = ( (~ e)  &  f  &  (~ h) ) ;
 assign n_n662 = ( (~ f)  &  (~ h)  &  i ) ;
 assign wire282 = ( j  &  (~ k)  &  (~ m)  &  (~ n) ) ;
 assign wire373 = ( (~ h)  &  (~ i)  &  (~ j)  &  l ) ;
 assign n_n1180 = ( i  &  (~ j)  &  (~ k) ) ;
 assign n_n1196 = ( (~ e)  &  g  &  h ) ;
 assign wire204 = ( f ) | ( (~ m) ) | ( n ) ;
 assign wire227 = ( j  &  (~ k)  &  (~ m)  &  n ) ;
 assign n_n1121 = ( (~ b)  &  e  &  (~ f) ) ;
 assign n_n1164 = ( c  &  (~ e)  &  (~ f) ) ;
 assign n_n1222 = ( (~ k)  &  m  &  (~ n) ) ;
 assign n_n1095 = ( f  &  (~ h)  &  i ) ;
 assign wire221 = ( (~ j)  &  k  &  (~ m)  &  n ) ;
 assign wire234 = ( h ) | ( i ) | ( j ) ;
 assign wire285 = ( (~ i)  &  (~ k)  &  (~ m)  &  n ) ;
 assign wire286 = ( (~ h)  &  (~ i)  &  (~ m)  &  n ) ;
 assign wire301 = ( (~ k)  &  (~ l)  &  (~ m)  &  n ) ;
 assign n_n1148 = ( e  &  g  &  h ) ;
 assign n_n1191 = ( k  &  (~ m)  &  (~ n) ) ;
 assign n_n1133 = ( i  &  (~ j)  &  k ) ;
 assign n_n819 = ( (~ g)  &  h  &  (~ j) ) ;
 assign n_n1131 = ( g  &  i  &  k ) ;
 assign wire79 = ( (~ c)  &  d  &  (~ e) ) | ( c  &  e  &  (~ f) ) ;
 assign wire158 = ( (~ c)  &  g  &  h ) | ( (~ f)  &  g  &  h ) ;
 assign wire170 = ( (~ j)  &  (~ m)  &  (~ n) ) ;
 assign wire194 = ( (~ g)  &  h ) ;
 assign n_n1243 = ( (~ i)  &  (~ k)  &  (~ m) ) ;
 assign n_n1227 = ( j  &  (~ k)  &  (~ m) ) ;
 assign n_n1091 = ( (~ c)  &  (~ f)  &  (~ g) ) ;
 assign wire95 = ( c  &  (~ f) ) | ( (~ c)  &  g ) ;
 assign wire226 = ( (~ h)  &  (~ i)  &  (~ m)  &  (~ n) ) ;
 assign wire395 = ( (~ c)  &  (~ d) ) | ( (~ c)  &  (~ f) ) ;
 assign n_n818 = ( (~ g)  &  h  &  j ) ;
 assign n_n529 = ( g  &  (~ i)  &  j ) ;
 assign n_n670 = ( h  &  (~ i)  &  j ) ;
 assign wire23 = ( g  &  (~ h)  &  i ) | ( g  &  h  &  (~ i) ) ;
 assign wire59 = ( f  &  (~ h)  &  i ) | ( f  &  h  &  (~ i) ) ;
 assign wire96 = ( (~ k)  &  m  &  (~ n) ) | ( l  &  m  &  (~ n) ) ;
 assign wire134 = ( (~ g)  &  (~ h)  &  i ) | ( (~ g)  &  h  &  (~ i) ) ;
 assign wire398 = ( (~ h)  &  i  &  j ) ;
 assign n_n387 = ( g  &  (~ j)  &  k ) ;
 assign n_n694 = ( g  &  i  &  (~ j) ) ;
 assign wire72 = ( n_n1219  &  n_n387 ) | ( n_n1220  &  n_n694 ) ;
 assign wire47 = ( b  &  (~ c)  &  d ) | ( b  &  c  &  (~ d) ) | ( b  &  (~ d)  &  e ) ;
 assign wire211 = ( (~ g)  &  n_n711  &  wire146 ) | ( g  &  wire146  &  wire47 ) ;
 assign wire231 = ( (~ f)  &  h  &  (~ i) ) | ( (~ f)  &  h  &  (~ j) ) ;
 assign wire137 = ( (~ g) ) | ( (~ j) ) ;
 assign n_n1118 = ( (~ k)  &  (~ l)  &  (~ m) ) ;
 assign n_n1216 = ( l  &  (~ m)  &  n ) ;
 assign n_n868 = ( j  &  (~ l)  &  m ) ;
 assign n_n1094 = ( (~ g)  &  (~ h)  &  i ) ;
 assign wire249 = ( c  &  (~ d) ) ;
 assign n_n628 = ( c  &  (~ d)  &  f ) ;
 assign wire396 = ( b  &  (~ c) ) ;
 assign n_n1146 = ( j  &  k  &  l ) ;
 assign wire121 = ( h  &  k ) ;
 assign n_n1116 = ( i  &  k  &  (~ m) ) ;
 assign n_n940 = ( e  &  f  &  (~ g) ) ;
 assign n_n765 = ( f  &  g  &  j ) ;
 assign wire248 = ( (~ m)  &  n  &  n_n1253  &  n_n1252 ) ;
 assign wire55 = ( j  &  (~ k)  &  l ) | ( (~ j)  &  k  &  (~ l) ) ;
 assign wire149 = ( (~ i)  &  j  &  (~ k) ) | ( (~ i)  &  j  &  l ) ;
 assign wire18 = ( i  &  (~ j)  &  k ) | ( i  &  k  &  (~ l) ) ;
 assign n_n874 = ( i  &  l  &  m ) ;
 assign n_n605 = ( j  &  (~ k)  &  (~ l) ) ;
 assign n_n1084 = ( (~ f)  &  h  &  (~ j) ) ;
 assign n_n875 = ( e  &  g  &  (~ h) ) ;
 assign n_n871 = ( (~ i)  &  l  &  m ) ;
 assign n_n235 = ( h  &  k  &  (~ l) ) ;
 assign n_n2572 = ( wire113  &  n_n876  &  n_n859 ) ;
 assign wire5830 = ( (~ k)  &  (~ l)  &  m  &  (~ n) ) ;
 assign n_n2953 = ( n_n698  &  n_n1137  &  wire5830 ) ;
 assign n_n1167 = ( (~ c)  &  e  &  (~ f) ) ;
 assign n_n1189 = ( (~ a)  &  d  &  (~ e) ) ;
 assign n_n703 = ( b  &  (~ e)  &  f ) ;
 assign wire197 = ( g  &  (~ j) ) ;
 assign wire161 = ( (~ k)  &  m  &  (~ n) ) | ( (~ l)  &  m  &  (~ n) ) ;
 assign wire305 = ( (~ c)  &  (~ d)  &  i ) ;
 assign wire399 = ( (~ g)  &  (~ k)  &  m  &  (~ n) ) ;
 assign wire414 = ( e  &  g  &  i  &  _7925 ) ;
 assign wire369 = ( a  &  c  &  (~ d)  &  e ) ;
 assign n_n2660 = ( g  &  j  &  wire58  &  wire369 ) ;
 assign n_n982 = ( (~ k)  &  l  &  (~ m)  &  n ) ;
 assign n_n919 = ( d  &  (~ e)  &  g ) ;
 assign n_n844 = ( k  &  (~ l)  &  (~ m) ) ;
 assign wire35 = ( c  &  e  &  (~ f) ) | ( c  &  f  &  (~ g) ) ;
 assign wire6251 = ( wire322 ) | ( wire6245 ) | ( _8939  &  _8940 ) ;
 assign wire6252 = ( wire328 ) | ( wire330 ) | ( wire6246 ) ;
 assign wire6256 = ( wire307 ) | ( wire6248 ) | ( wire6249 ) | ( wire6250 ) ;
 assign wire56 = ( (~ h)  &  i  &  k ) | ( h  &  j  &  (~ k) ) ;
 assign wire142 = ( k  &  l  &  m  &  (~ n) ) ;
 assign wire216 = ( (~ g)  &  h  &  (~ j) ) | ( (~ g)  &  h  &  k ) | ( g  &  j  &  (~ k) ) ;
 assign wire260 = ( (~ j)  &  l  &  (~ m)  &  (~ n) ) ;
 assign wire181 = ( wire20 ) | ( (~ i)  &  j  &  (~ k) ) ;
 assign wire104 = ( (~ e)  &  g  &  h ) | ( f  &  g  &  h ) ;
 assign wire293 = ( (~ j)  &  k  &  (~ m)  &  n ) | ( j  &  (~ k)  &  (~ m)  &  n ) ;
 assign wire43 = ( (~ a)  &  b  &  (~ d) ) | ( (~ a)  &  b  &  e ) ;
 assign wire24 = ( (~ c)  &  d  &  f ) | ( c  &  (~ e)  &  f ) ;
 assign wire49 = ( (~ i)  &  k  &  (~ m) ) | ( (~ j)  &  k  &  (~ m) ) | ( j  &  (~ k)  &  (~ m) ) ;
 assign wire109 = ( (~ c)  &  d  &  (~ e) ) | ( (~ c)  &  d  &  f ) | ( c  &  (~ e)  &  f ) | ( c  &  e  &  (~ f) ) ;
 assign wire206 = ( (~ g)  &  h  &  i ) | ( g  &  i  &  (~ j) ) ;
 assign wire105 = ( (~ g)  &  h  &  (~ j) ) | ( g  &  j  &  (~ k) ) ;
 assign wire152 = ( (~ l)  &  n_n1187  &  n_n1137 ) | ( l  &  n_n1187  &  wire23 ) ;
 assign wire299 = ( a  &  (~ c)  &  d  &  _7541 ) ;
 assign wire388 = ( n_n918  &  n_n1187  &  n_n1249 ) | ( n_n918  &  n_n1187  &  n_n1231 ) ;
 assign wire162 = ( wire282 ) | ( (~ n_n1264)  &  n_n1191 ) ;
 assign wire198 = ( h  &  j  &  (~ k) ) | ( h  &  k  &  (~ l) ) ;
 assign wire377 = ( (~ f)  &  g  &  h  &  n_n711 ) | ( (~ f)  &  (~ g)  &  h  &  n_n711 ) ;
 assign wire385 = ( (~ f)  &  g  &  h  &  (~ n) ) ;
 assign wire16 = ( a  &  (~ c)  &  d ) | ( a  &  d  &  (~ e) ) ;
 assign wire60 = ( (~ b)  &  c  &  (~ e) ) | ( b  &  e  &  (~ f) ) ;
 assign wire69 = ( wire54  &  n_n1082 ) | ( wire148  &  n_n875 ) ;
 assign wire81 = ( wire265  &  n_n1155 ) | ( wire58  &  n_n1137 ) ;
 assign wire85 = ( (~ j)  &  m  &  (~ n) ) | ( k  &  m  &  (~ n) ) ;
 assign wire115 = ( n_n713  &  n_n886 ) | ( n_n1253  &  n_n1083 ) ;
 assign wire368 = ( e  &  g  &  h  &  (~ n) ) ;
 assign wire6310 = ( (~ i)  &  (~ j)  &  (~ k) ) ;
 assign wire42 = ( n_n971  &  n_n973  &  n_n1204  &  wire6310 ) ;
 assign wire61 = ( n_n1165  &  n_n1138  &  n_n1142  &  n_n1146 ) ;
 assign wire63 = ( n_n1138  &  wire254  &  wire407 ) ;
 assign wire66 = ( n_n988  &  n_n1028  &  wire384  &  n_n982 ) ;
 assign wire6287 = ( c  &  h  &  (~ j) ) | ( d  &  h  &  (~ j) ) ;
 assign wire140 = ( n_n1202  &  (~ wire268)  &  wire6287 ) ;
 assign wire6289 = ( (~ c)  &  g  &  h ) | ( (~ d)  &  g  &  h ) ;
 assign wire150 = ( m  &  (~ n)  &  n_n1180  &  wire6289 ) ;
 assign wire163 = ( (~ c)  &  (~ d)  &  n_n1155  &  wire127 ) ;
 assign wire173 = ( (~ a)  &  (~ b)  &  m  &  (~ n) ) ;
 assign wire177 = ( (~ b)  &  (~ c)  &  (~ m)  &  n ) ;
 assign wire178 = ( (~ g)  &  (~ h)  &  m  &  (~ n) ) ;
 assign wire180 = ( (~ l)  &  m  &  (~ n)  &  _8794 ) ;
 assign wire6257 = ( g ) | ( (~ f)  &  h ) ;
 assign wire6258 = ( (~ i)  &  (~ k)  &  (~ m)  &  (~ n) ) ;
 assign wire252 = ( (~ n_n861)  &  wire395  &  wire6257  &  wire6258 ) ;
 assign wire6262 = ( h  &  (~ j)  &  (~ k)  &  (~ m) ) ;
 assign wire6263 = ( (~ g)  &  (~ h) ) | ( (~ g)  &  i ) | ( g  &  (~ i) ) | ( (~ h)  &  (~ i) ) | ( g  &  j ) | ( (~ h)  &  j ) | ( i  &  j ) ;
 assign wire253 = ( wire6262  &  wire6263 ) ;
 assign wire6264 = ( (~ g)  &  (~ i)  &  (~ m)  &  (~ n) ) ;
 assign wire269 = ( wire395  &  (~ n_n1118)  &  wire6264 ) ;
 assign wire6266 = ( (~ c)  &  (~ d)  &  g ) ;
 assign wire271 = ( wire127  &  (~ n_n765)  &  wire6266 ) ;
 assign wire6268 = ( c  &  (~ g)  &  (~ h) ) | ( f  &  (~ g)  &  (~ h) ) ;
 assign wire272 = ( wire254  &  wire6268 ) ;
 assign wire274 = ( h  &  (~ j)  &  (~ wire127)  &  n_n1118 ) ;
 assign wire276 = ( wire127  &  _9185 ) | ( wire127  &  _9186 ) ;
 assign wire6272 = ( h  &  (~ i)  &  (~ m)  &  (~ n) ) ;
 assign wire278 = ( n_n1194  &  n_n1202  &  n_n819 ) ;
 assign wire280 = ( n_n1202  &  n_n1083  &  n_n694 ) ;
 assign wire281 = ( c  &  (~ e)  &  (~ f)  &  _9203 ) ;
 assign wire6211 = ( i  &  (~ m)  &  (~ n) ) ;
 assign wire6216 = ( (~ n_n857)  &  (~ n_n1260)  &  (~ wire35) ) ;
 assign wire6217 = ( (~ n_n766)  &  (~ n_n919)  &  wire6213 ) ;
 assign wire307 = ( (~ n_n912)  &  wire6211  &  wire6216  &  wire6217 ) ;
 assign wire6225 = ( i  &  j  &  (~ m)  &  (~ n) ) ;
 assign wire6226 = ( c ) | ( (~ d) ) ;
 assign wire6227 = ( c  &  (~ f) ) | ( (~ f)  &  g ) | ( c  &  (~ g) ) | ( f  &  (~ g) ) | ( c  &  (~ j) ) | ( f  &  (~ j) ) | ( g  &  (~ j) ) ;
 assign wire316 = ( (~ wire35)  &  wire6225  &  wire6226  &  wire6227 ) ;
 assign wire6230 = ( (~ c)  &  (~ f) ) ;
 assign wire317 = ( n_n1190  &  (~ wire127)  &  (~ n_n919)  &  wire6230 ) ;
 assign wire6233 = ( (~ a)  &  m  &  (~ n) ) ;
 assign wire318 = ( (~ e)  &  (~ f)  &  wire234  &  wire6233 ) ;
 assign wire6236 = ( (~ d)  &  j ) | ( e  &  j ) | ( (~ g)  &  j ) ;
 assign wire322 = ( (~ m)  &  (~ n)  &  n_n1164  &  wire6236 ) ;
 assign wire328 = ( (~ m)  &  n  &  n_n1069  &  n_n940 ) ;
 assign wire330 = ( m  &  (~ n)  &  n_n700  &  n_n1189 ) ;
 assign wire6177 = ( (~ f)  &  (~ g)  &  (~ m)  &  n ) ;
 assign wire333 = ( (~ n_n1171)  &  (~ n_n700)  &  (~ n_n973)  &  wire6177 ) ;
 assign wire6180 = ( f ) | ( (~ b)  &  e ) ;
 assign wire334 = ( (~ wire263)  &  wire286  &  n_n1216  &  wire6180 ) ;
 assign wire6185 = ( (~ b)  &  (~ f)  &  (~ m)  &  n ) ;
 assign wire336 = ( (~ n_n1249)  &  (~ n_n1216)  &  wire6185 ) ;
 assign wire6187 = ( (~ c)  &  (~ e)  &  (~ f) ) | ( d  &  (~ e)  &  (~ f) ) ;
 assign wire6188 = ( (~ a)  &  (~ f)  &  m  &  (~ n) ) ;
 assign wire337 = ( wire6187  &  wire6188 ) ;
 assign wire338 = ( (~ wire407)  &  wire170  &  wire226 ) ;
 assign wire339 = ( a  &  j  &  wire399 ) | ( (~ b)  &  j  &  wire399 ) ;
 assign wire340 = ( n_n1210  &  wire286  &  (~ n_n1216) ) ;
 assign wire341 = ( (~ e)  &  wire286  &  (~ n_n1216) ) ;
 assign wire342 = ( n_n1171  &  n_n1056  &  wire286 ) ;
 assign wire6151 = ( (~ g)  &  (~ m)  &  (~ n) ) ;
 assign wire352 = ( (~ c)  &  (~ d)  &  f  &  wire6151 ) | ( (~ c)  &  d  &  (~ f)  &  wire6151 ) ;
 assign wire353 = ( j  &  wire232  &  wire399 ) ;
 assign wire354 = ( (~ c)  &  wire286 ) | ( (~ d)  &  wire286 ) ;
 assign wire355 = ( (~ wire204)  &  _8819 ) | ( (~ wire204)  &  _8820 ) ;
 assign wire357 = ( (~ c)  &  (~ d)  &  n_n1190  &  (~ n_n1091) ) ;
 assign wire362 = ( (~ e)  &  (~ f)  &  (~ g)  &  _8835 ) ;
 assign wire389 = ( c  &  (~ e)  &  (~ f)  &  _8823 ) ;
 assign wire6109 = ( f  &  g  &  h ) ;
 assign wire429 = ( n_n1217  &  (~ n_n1260)  &  n_n1215  &  wire6109 ) ;
 assign wire6112 = ( (~ a)  &  f  &  g  &  h ) ;
 assign wire430 = ( n_n1217  &  n_n1215  &  wire6112 ) ;
 assign wire431 = ( n_n1217  &  wire196  &  n_n1264  &  n_n1216 ) ;
 assign wire6115 = ( h  &  j ) | ( i  &  j ) ;
 assign wire432 = ( n_n1253  &  wire6115  &  _8855 ) ;
 assign wire6118 = ( (~ e)  &  (~ f)  &  (~ h)  &  (~ j) ) ;
 assign wire433 = ( (~ m)  &  n  &  n_n1253  &  wire6118 ) ;
 assign wire6119 = ( c  &  d  &  e  &  (~ n) ) ;
 assign wire434 = ( n_n1228  &  n_n1227  &  wire6119 ) ;
 assign wire435 = ( n_n1253  &  n_n1249  &  _8880 ) ;
 assign wire440 = ( n_n1261  &  n_n1260  &  _8868 ) ;
 assign wire441 = ( n_n1253  &  n_n1249  &  wire285 ) ;
 assign wire442 = ( n_n1253  &  n_n1252  &  _8851 ) ;
 assign wire6072 = ( c  &  (~ i)  &  (~ k) ) ;
 assign wire443 = ( n_n1022  &  n_n1204  &  wire6072 ) ;
 assign wire444 = ( _8746  &  _8747 ) ;
 assign wire445 = ( (~ d)  &  (~ e)  &  n_n1261  &  _8748 ) ;
 assign wire6078 = ( (~ d)  &  h ) | ( (~ e)  &  h ) | ( (~ f)  &  h ) ;
 assign wire446 = ( n_n1217  &  n_n1204  &  (~ n_n1091)  &  wire6078 ) ;
 assign wire447 = ( n_n1207  &  n_n1229  &  _8750 ) ;
 assign wire6082 = ( (~ e)  &  (~ f)  &  i ) | ( (~ e)  &  (~ f)  &  (~ j) ) ;
 assign wire448 = ( n_n1253  &  n_n1210  &  wire6082 ) ;
 assign wire449 = ( n_n1203  &  n_n1202  &  wire384 ) ;
 assign wire6085 = ( a  &  (~ f)  &  m  &  (~ n) ) ;
 assign wire450 = ( wire373  &  wire6085 ) ;
 assign wire451 = ( (~ n_n1188)  &  n_n1229  &  n_n1193  &  n_n1190 ) ;
 assign wire452 = ( n_n1217  &  (~ n_n1138)  &  n_n1204  &  wire194 ) ;
 assign wire453 = ( _8731  &  _8732 ) ;
 assign wire454 = ( n_n1229  &  n_n1228  &  wire170 ) ;
 assign wire455 = ( n_n1229  &  n_n1193  &  n_n1204 ) ;
 assign wire456 = ( n_n1229  &  n_n1201  &  n_n1190 ) ;
 assign wire457 = ( n_n1217  &  n_n1215  &  wire158 ) ;
 assign wire458 = ( m  &  (~ n)  &  n_n1188  &  n_n1189 ) ;
 assign wire459 = ( n_n1253  &  n_n1252  &  _8742 ) ;
 assign wire460 = ( n_n1217  &  n_n1204  &  wire158 ) ;
 assign wire6042 = ( (~ d)  &  (~ f)  &  g  &  (~ h) ) ;
 assign wire461 = ( (~ n_n1203)  &  n_n1204  &  (~ n_n1227)  &  wire6042 ) ;
 assign wire6047 = ( (~ h)  &  i  &  (~ m)  &  (~ n) ) ;
 assign wire463 = ( (~ n_n857)  &  wire395  &  wire6047 ) ;
 assign wire465 = ( n_n1161  &  wire226  &  wire395 ) ;
 assign wire466 = ( (~ wire95)  &  wire226  &  _9007 ) ;
 assign wire467 = ( g  &  (~ h)  &  n_n1204  &  n_n1243 ) ;
 assign wire6054 = ( c  &  (~ f)  &  (~ h) ) | ( (~ c)  &  g  &  (~ h) ) ;
 assign wire469 = ( n_n1190  &  wire95  &  wire226 ) ;
 assign wire6005 = ( (~ c)  &  e  &  (~ f) ) | ( c  &  (~ e)  &  (~ f) ) ;
 assign wire480 = ( n_n1133  &  wire170  &  wire6005 ) ;
 assign wire6006 = ( c  &  (~ g)  &  h ) ;
 assign wire481 = ( n_n1159  &  wire170  &  wire6006 ) ;
 assign wire482 = ( n_n861  &  (~ n_n1080)  &  (~ wire79)  &  wire170 ) ;
 assign wire6010 = ( c  &  i ) | ( d  &  i ) | ( e  &  i ) ;
 assign wire483 = ( n_n1072  &  wire170  &  wire6010 ) ;
 assign wire6012 = ( c  &  (~ k)  &  (~ m)  &  (~ n) ) ;
 assign wire484 = ( n_n1082  &  wire170  &  wire6012 ) ;
 assign wire6014 = ( (~ f)  &  k  &  (~ m)  &  (~ n) ) ;
 assign wire485 = ( n_n1131  &  (~ wire79)  &  wire6014 ) ;
 assign wire486 = ( n_n861  &  (~ n_n1080)  &  n_n1202  &  (~ wire79) ) ;
 assign wire487 = ( n_n1165  &  n_n1195  &  n_n1137  &  (~ wire79) ) ;
 assign wire6020 = ( (~ e)  &  (~ f)  &  (~ g)  &  (~ i) ) ;
 assign wire488 = ( n_n1164  &  n_n1191  &  wire6020 ) ;
 assign wire6022 = ( (~ h)  &  (~ k)  &  m  &  (~ n) ) ;
 assign wire489 = ( m  &  (~ n)  &  n_n1189  &  wire6022 ) ;
 assign wire490 = ( (~ c)  &  d  &  n_n1202  &  n_n819 ) ;
 assign wire491 = ( n_n1159  &  wire158  &  wire170 ) ;
 assign wire492 = ( (~ n_n1260)  &  n_n1146  &  _9092 ) ;
 assign wire493 = ( n_n975  &  n_n1146  &  _9094 ) ;
 assign wire494 = ( m  &  (~ n)  &  n_n1195  &  n_n1180 ) ;
 assign wire495 = ( m  &  (~ n)  &  n_n1180  &  n_n1148 ) ;
 assign wire496 = ( (~ m)  &  n  &  n_n1142  &  n_n1146 ) ;
 assign wire5971 = ( (~ h)  &  i ) | ( (~ h)  &  (~ j) ) ;
 assign wire499 = ( n_n1121  &  wire5971  &  _9067 ) ;
 assign wire500 = ( n_n1036  &  wire146  &  (~ wire263)  &  (~ n_n1196) ) ;
 assign wire501 = ( wire54  &  (~ n_n1203)  &  (~ n_n1164)  &  (~ wire234) ) ;
 assign wire5979 = ( e  &  (~ f)  &  h  &  j ) ;
 assign wire504 = ( (~ m)  &  n  &  n_n1121  &  wire5979 ) ;
 assign wire505 = ( n_n1161  &  wire263  &  wire286 ) ;
 assign wire508 = ( (~ b)  &  wire54  &  (~ wire234) ) ;
 assign wire509 = ( n_n975  &  (~ wire204)  &  n_n1121 ) ;
 assign wire510 = ( (~ b)  &  f  &  (~ h)  &  wire70 ) ;
 assign wire512 = ( (~ m)  &  n  &  n_n1121  &  wire285 ) ;
 assign wire513 = ( (~ m)  &  n  &  n_n1121  &  wire221 ) ;
 assign wire516 = ( m  &  (~ n)  &  n_n1095  &  n_n1189 ) ;
 assign wire520 = ( (~ e)  &  h  &  wire263  &  n_n1180 ) ;
 assign wire5958 = ( d  &  (~ f)  &  m  &  (~ n) ) ;
 assign wire521 = ( wire373  &  wire5958 ) ;
 assign wire5959 = ( a  &  g  &  h ) | ( (~ b)  &  g  &  h ) ;
 assign wire522 = ( m  &  (~ n)  &  n_n1180  &  wire5959 ) ;
 assign wire523 = ( (~ b)  &  (~ j)  &  n_n1036  &  n_n1196 ) ;
 assign wire5964 = ( (~ e)  &  (~ f)  &  (~ l) ) ;
 assign wire527 = ( (~ m)  &  n  &  n_n1253  &  wire5964 ) ;
 assign wire5941 = ( (~ g)  &  (~ h)  &  (~ k) ) ;
 assign wire528 = ( (~ c)  &  d  &  n_n1190  &  wire5941 ) ;
 assign wire5946 = ( (~ d)  &  g  &  (~ h)  &  i ) ;
 assign wire532 = ( wire282  &  wire5946 ) ;
 assign wire533 = ( (~ m)  &  (~ n)  &  n_n1166  &  wire268 ) ;
 assign wire534 = ( i  &  j  &  n_n1161  &  n_n1202 ) ;
 assign wire535 = ( (~ m)  &  (~ n)  &  n_n1159  &  n_n1160 ) ;
 assign wire536 = ( n_n1220  &  n_n730  &  (~ n_n1053)  &  n_n816 ) ;
 assign wire537 = ( n_n700  &  wire21  &  wire290 ) ;
 assign wire539 = ( n_n841  &  n_n1210  &  wire36 ) ;
 assign wire540 = ( wire34  &  n_n1202  &  n_n1264 ) ;
 assign wire541 = ( n_n671  &  n_n1036  &  n_n1264 ) ;
 assign wire542 = ( n_n671  &  n_n1210  &  n_n619 ) ;
 assign wire543 = ( n_n671  &  n_n1210  &  n_n1085 ) ;
 assign wire544 = ( n_n841  &  n_n1210  &  n_n1053 ) ;
 assign wire545 = ( n_n904  &  n_n1220  &  n_n1194 ) ;
 assign wire546 = ( n_n711  &  n_n1142  &  wire70 ) | ( wire30  &  n_n1142  &  wire70 ) ;
 assign wire547 = ( wire34  &  n_n619  &  n_n1191 ) | ( n_n619  &  n_n1191  &  wire35 ) ;
 assign wire548 = ( wire34  &  n_n1085  &  n_n1191 ) | ( n_n1085  &  n_n1191  &  wire35 ) ;
 assign wire549 = ( m  &  (~ n)  &  n_n698  &  n_n816 ) ;
 assign wire550 = ( m  &  (~ n)  &  n_n698  &  n_n618 ) ;
 assign wire551 = ( n_n700  &  n_n841  &  n_n1191 ) ;
 assign wire552 = ( n_n992  &  wire36  &  wire70 ) ;
 assign wire554 = ( n_n709  &  wire230  &  n_n1210 ) ;
 assign wire565 = ( wire22  &  (~ wire29)  &  n_n730  &  wire146 ) ;
 assign wire566 = ( wire22  &  n_n918  &  (~ wire14)  &  wire146 ) ;
 assign wire567 = ( wire22  &  n_n1022  &  wire369 ) ;
 assign wire568 = ( n_n1187  &  n_n996  &  n_n1155  &  n_n698 ) ;
 assign wire569 = ( n_n992  &  n_n1053  &  wire293 ) ;
 assign wire5884 = ( (~ h)  &  (~ k) ) | ( j  &  (~ k) ) ;
 assign wire570 = ( n_n1201  &  wire15  &  n_n1187  &  wire5884 ) ;
 assign wire571 = ( n_n1171  &  n_n992  &  wire221 ) | ( n_n992  &  wire221  &  wire47 ) ;
 assign wire5886 = ( (~ h)  &  (~ k) ) | ( j  &  (~ k) ) ;
 assign wire572 = ( wire25  &  n_n1187  &  wire5886 ) | ( wire32  &  n_n1187  &  wire5886 ) ;
 assign wire573 = ( n_n1201  &  wire29  &  n_n1187  &  n_n996 ) ;
 assign wire575 = ( wire22  &  wire29  &  n_n1022 ) ;
 assign wire576 = ( wire22  &  wire14  &  n_n1084 ) ;
 assign wire577 = ( n_n904  &  wire22  &  n_n1022 ) ;
 assign wire5813 = ( f  &  h  &  i ) ;
 assign wire580 = ( wire25  &  n_n1187  &  n_n996 ) | ( wire32  &  n_n1187  &  n_n996 ) ;
 assign wire1016 = ( m  &  (~ n)  &  n_n920  &  n_n1201 ) ;
 assign wire583 = ( g  &  h  &  i  &  wire113 ) ;
 assign wire585 = ( wire22  &  wire210  &  wire14  &  wire197 ) ;
 assign wire586 = ( wire22  &  n_n987  &  wire14  &  wire197 ) ;
 assign wire587 = ( n_n904  &  wire22  &  (~ n_n987)  &  wire197 ) ;
 assign wire5857 = ( a  &  b  &  d  &  (~ e) ) ;
 assign wire588 = ( g  &  (~ j)  &  wire22  &  wire5857 ) ;
 assign wire590 = ( n_n711  &  n_n1142  &  wire70 ) ;
 assign wire593 = ( n_n920  &  wire22  &  n_n766 ) ;
 assign wire594 = ( wire210  &  n_n992  &  wire70 ) ;
 assign wire598 = ( n_n840  &  n_n1210  &  n_n1022 ) ;
 assign wire610 = ( n_n1201  &  wire29  &  n_n1187  &  n_n605 ) ;
 assign wire5839 = ( i  &  k  &  m  &  (~ n) ) ;
 assign wire611 = ( wire41  &  wire5839 ) | ( wire1012  &  wire5839 ) | ( wire299  &  wire5839 ) ;
 assign wire617 = ( n_n1220  &  n_n698  &  n_n841 ) ;
 assign wire618 = ( wire25  &  n_n1187  &  n_n605 ) | ( wire32  &  n_n1187  &  n_n605 ) ;
 assign wire619 = ( n_n918  &  n_n1187  &  n_n1195  &  n_n605 ) ;
 assign wire626 = ( n_n700  &  wire290  &  n_n1227 ) ;
 assign wire627 = ( n_n1155  &  n_n1210  &  wire47 ) | ( n_n1155  &  n_n1210  &  wire60 ) ;
 assign wire628 = ( n_n711  &  n_n821  &  n_n1210 ) | ( n_n821  &  wire30  &  n_n1210 ) ;
 assign wire629 = ( n_n671  &  n_n1036  &  n_n1264 ) ;
 assign wire630 = ( n_n1210  &  n_n820  &  n_n1053 ) ;
 assign wire631 = ( n_n1171  &  n_n1219  &  n_n387 ) ;
 assign wire632 = ( wire30  &  n_n1142  &  wire70 ) ;
 assign wire633 = ( n_n709  &  n_n1210  &  wire231 ) ;
 assign wire635 = ( n_n840  &  n_n824  &  n_n1210 ) ;
 assign wire643 = ( n_n1080  &  n_n1190  &  n_n1039  &  wire386 ) ;
 assign wire644 = ( n_n838  &  (~ n_n1252)  &  n_n1210  &  wire89 ) ;
 assign wire5781 = ( a  &  b  &  d  &  (~ e) ) ;
 assign wire645 = ( (~ g)  &  wire190  &  wire5781 ) ;
 assign wire646 = ( n_n1187  &  n_n949  &  n_n1252  &  wire165 ) ;
 assign wire647 = ( n_n842  &  n_n1210  &  wire164 ) ;
 assign wire649 = ( n_n1187  &  n_n987  &  n_n949  &  wire39 ) ;
 assign wire650 = ( n_n1187  &  n_n987  &  n_n949  &  n_n977 ) ;
 assign wire651 = ( n_n988  &  n_n1210  &  wire89 ) ;
 assign wire652 = ( n_n1217  &  n_n971  &  n_n1080  &  n_n1204 ) ;
 assign wire653 = ( (~ g)  &  wire224  &  wire190 ) ;
 assign wire5694 = ( wire54  &  n_n971 ) | ( wire31  &  wire385 ) ;
 assign wire655 = ( n_n872  &  wire5694 ) | ( wire148  &  n_n1104  &  n_n872 ) ;
 assign wire743 = ( (~ l)  &  m  &  (~ n)  &  _8344 ) ;
 assign wire1116 = ( wire31  &  wire368 ) ;
 assign wire663 = ( _331 ) | ( n_n1187  &  n_n949  &  wire69 ) ;
 assign wire664 = ( n_n876  &  wire69 ) | ( wire31  &  n_n876  &  wire368 ) ;
 assign wire670 = ( wire283  &  n_n1253  &  n_n1252  &  wire301 ) ;
 assign wire671 = ( n_n1201  &  n_n1069  &  n_n1204  &  n_n1180 ) ;
 assign wire672 = ( n_n1207  &  n_n1229  &  n_n1190  &  n_n977 ) ;
 assign wire679 = ( wire76  &  n_n838  &  _8439 ) ;
 assign wire680 = ( wire58  &  n_n857  &  n_n872  &  (~ wire137) ) ;
 assign wire681 = ( n_n1161  &  wire84  &  n_n988 ) ;
 assign wire682 = ( n_n988  &  wire77  &  n_n1196 ) ;
 assign wire683 = ( n_n842  &  wire76  &  n_n841 ) ;
 assign wire684 = ( wire22  &  n_n857  &  n_n872 ) | ( wire113  &  n_n857  &  n_n872 ) ;
 assign wire699 = ( n_n904  &  n_n1187  &  wire74  &  n_n1252 ) ;
 assign wire701 = ( n_n942  &  n_n904  &  n_n1187  &  n_n940 ) ;
 assign wire702 = ( n_n1161  &  n_n893  &  n_n1177  &  n_n988 ) ;
 assign wire704 = ( n_n920  &  n_n1187  &  n_n1233  &  wire18 ) ;
 assign wire708 = ( n_n1187  &  n_n949  &  n_n1252  &  wire55 ) ;
 assign wire709 = ( n_n1187  &  n_n989  &  n_n987  &  n_n949 ) ;
 assign wire1112 = ( wire228  &  n_n864 ) | ( wire265  &  n_n864 ) ;
 assign wire1113 = ( wire22  &  n_n859 ) | ( wire113  &  n_n859 ) ;
 assign wire5690 = ( c  &  d  &  wire120 ) ;
 assign wire713 = ( wire417  &  wire1112  &  wire5690 ) | ( wire417  &  wire1113  &  wire5690 ) ;
 assign wire716 = ( wire120  &  wire183  &  n_n1231  &  (~ wire57) ) ;
 assign wire5699 = ( a  &  b  &  c  &  d ) ;
 assign wire718 = ( n_n1165  &  n_n1138  &  n_n1142  &  n_n1146 ) ;
 assign wire719 = ( n_n1138  &  wire254  &  wire407 ) ;
 assign wire724 = ( n_n1220  &  n_n997  &  n_n1082 ) ;
 assign wire1068 = ( i  &  l  &  m  &  wire5252 ) ;
 assign wire5253 = ( wire54  &  n_n1194 ) | ( wire31  &  wire5251 ) ;
 assign wire725 = ( wire390  &  n_n949 ) | ( n_n949  &  wire1068 ) | ( n_n949  &  wire5253 ) ;
 assign wire726 = ( wire58  &  n_n949  &  n_n765 ) ;
 assign wire727 = ( _373 ) | ( wire379  &  _8370 ) ;
 assign wire729 = ( _405 ) | ( n_n1220  &  n_n876  &  n_n1082 ) ;
 assign wire731 = ( n_n997  &  wire69 ) | ( wire31  &  n_n997  &  wire368 ) ;
 assign wire732 = ( n_n876  &  wire69 ) | ( wire31  &  n_n876  &  wire368 ) ;
 assign wire736 = ( wire22  &  n_n876  &  n_n859 ) ;
 assign wire739 = ( (~ f)  &  g  &  (~ h)  &  wire148 ) ;
 assign wire5674 = ( c  &  d  &  (~ f)  &  g ) ;
 assign wire745 = ( n_n1261  &  n_n1187  &  wire74  &  wire5674 ) ;
 assign wire749 = ( n_n1201  &  n_n1069  &  n_n1204  &  n_n1180 ) ;
 assign wire750 = ( n_n1187  &  wire74  &  n_n1233  &  n_n997 ) ;
 assign wire5663 = ( (~ c)  &  (~ d)  &  (~ e)  &  (~ i) ) ;
 assign wire5664 = ( (~ k)  &  (~ l)  &  (~ m)  &  (~ n) ) ;
 assign wire754 = ( n_n1217  &  n_n1069  &  n_n971  &  n_n1204 ) ;
 assign wire766 = ( n_n1159  &  wire226  &  _8290 ) ;
 assign wire767 = ( n_n1217  &  n_n971  &  n_n1080  &  n_n1204 ) ;
 assign wire5640 = ( i  &  j  &  (~ k) ) ;
 assign wire781 = ( n_n987  &  n_n988  &  n_n1085  &  n_n982 ) ;
 assign wire782 = ( n_n1195  &  n_n975  &  n_n1204  &  n_n1180 ) ;
 assign wire5587 = ( c  &  (~ d)  &  e ) ;
 assign wire783 = ( n_n1207  &  n_n893  &  n_n1165  &  wire5587 ) ;
 assign wire5590 = ( i  &  j  &  (~ k) ) ;
 assign wire784 = ( n_n1201  &  wire29  &  n_n1187  &  wire5590 ) ;
 assign wire5592 = ( i  &  j  &  (~ k) ) ;
 assign wire785 = ( n_n1201  &  n_n1187  &  n_n698  &  wire5592 ) ;
 assign wire786 = ( n_n893  &  wire148  &  wire29  &  n_n1194 ) ;
 assign wire787 = ( n_n893  &  wire148  &  n_n698  &  n_n1194 ) ;
 assign wire5598 = ( i  &  k  &  m  &  (~ n) ) ;
 assign wire788 = ( wire15  &  n_n1194  &  wire5598 ) ;
 assign wire789 = ( n_n1207  &  wire148  &  n_n1228  &  wire15 ) ;
 assign wire5600 = ( i  &  j  &  (~ k) ) ;
 assign wire790 = ( wire25  &  n_n1187  &  wire5600 ) | ( wire32  &  n_n1187  &  wire5600 ) ;
 assign wire5601 = ( i  &  j  &  (~ k) ) ;
 assign wire791 = ( n_n918  &  n_n1187  &  n_n1195  &  wire5601 ) ;
 assign wire796 = ( wire76  &  n_n841  &  wire93 ) ;
 assign wire797 = ( wire22  &  n_n1228  &  wire15 ) | ( wire113  &  n_n1228  &  wire15 ) ;
 assign wire5557 = ( n_n1161  &  n_n713 ) | ( wire396  &  n_n875 ) ;
 assign wire798 = ( _446 ) | ( n_n893  &  n_n1177  &  wire5557 ) ;
 assign wire799 = ( wire371  &  wire33 ) | ( wire33  &  wire80 ) | ( wire33  &  wire414 ) ;
 assign wire802 = ( wire148  &  wire41 ) | ( wire148  &  wire1012 ) | ( wire148  &  wire299 ) ;
 assign wire5526 = ( c  &  (~ d)  &  e  &  (~ n) ) ;
 assign wire808 = ( n_n1201  &  wire49  &  wire5526 ) ;
 assign wire5529 = ( c  &  (~ d)  &  e  &  (~ n) ) ;
 assign wire809 = ( n_n1201  &  n_n844  &  wire5529 ) ;
 assign wire5532 = ( c  &  (~ d)  &  e  &  (~ n) ) ;
 assign wire810 = ( n_n1207  &  n_n1116  &  wire5532 ) ;
 assign wire5534 = ( g  &  i  &  j ) ;
 assign wire811 = ( wire58  &  n_n1171  &  wire5534 ) ;
 assign wire812 = ( b  &  (~ c)  &  n_n1148  &  wire293 ) ;
 assign wire813 = ( b  &  (~ c)  &  wire172  &  n_n1148 ) ;
 assign wire814 = ( b  &  (~ c)  &  wire77  &  n_n1148 ) ;
 assign wire815 = ( n_n713  &  n_n1196  &  wire293 ) ;
 assign wire816 = ( n_n840  &  n_n1201  &  wire293 ) ;
 assign wire817 = ( n_n1171  &  wire290  &  n_n868 ) ;
 assign wire818 = ( n_n841  &  wire260  &  wire109 ) ;
 assign wire821 = ( n_n713  &  wire172  &  n_n1196 ) ;
 assign wire822 = ( n_n840  &  wire172  &  n_n1201 ) ;
 assign wire823 = ( wire93  &  n_n1210  &  wire164 ) ;
 assign wire826 = ( n_n713  &  wire77  &  n_n1196 ) ;
 assign wire827 = ( n_n840  &  n_n1201  &  wire77 ) ;
 assign wire828 = ( wire54  &  n_n1171  &  n_n1142 ) ;
 assign wire829 = ( n_n1190  &  n_n817  &  wire24 ) ;
 assign wire830 = ( n_n698  &  n_n1219  &  n_n1131 ) ;
 assign wire831 = ( n_n700  &  n_n1190  &  n_n817 ) ;
 assign wire832 = ( n_n1203  &  n_n1190  &  n_n817 ) ;
 assign wire833 = ( n_n1171  &  n_n1219  &  n_n1131 ) ;
 assign wire834 = ( n_n1202  &  n_n1137  &  wire109 ) ;
 assign wire835 = ( n_n698  &  n_n841  &  n_n1215 ) ;
 assign wire836 = ( wire84  &  wire5557 ) | ( n_n840  &  n_n1207  &  wire84 ) ;
 assign wire837 = ( n_n1171  &  n_n841  &  n_n1215 ) ;
 assign wire5480 = ( c  &  e  &  f  &  g ) ;
 assign wire843 = ( (~ n_n1229)  &  wire74  &  wire120  &  wire5480 ) ;
 assign wire5486 = ( d  &  f  &  g ) ;
 assign wire845 = ( wire74  &  wire120  &  wire196  &  wire5486 ) ;
 assign wire849 = ( n_n730  &  wire112  &  wire120  &  wire183 ) ;
 assign wire5498 = ( (~ b)  &  c  &  e  &  f ) ;
 assign wire850 = ( wire76  &  n_n1095  &  wire5498 ) ;
 assign wire853 = ( n_n1165  &  wire65  &  n_n1203 ) | ( n_n1165  &  n_n1203  &  n_n235 ) ;
 assign wire854 = ( n_n842  &  wire84  &  n_n1104 ) ;
 assign wire858 = ( wire390  &  n_n730 ) | ( n_n730  &  wire1068 ) | ( n_n730  &  wire5253 ) ;
 assign wire859 = ( n_n920  &  n_n1187  &  wire74  &  n_n1233 ) ;
 assign wire869 = ( n_n842  &  n_n1177  &  n_n1252  &  n_n235 ) ;
 assign wire5454 = ( (~ b)  &  c  &  e ) ;
 assign wire879 = ( n_n1203  &  n_n1166  &  n_n1204 ) ;
 assign wire880 = ( n_n709  &  n_n1210  &  wire231 ) ;
 assign wire884 = ( n_n709  &  n_n1210  &  n_n662 ) ;
 assign wire886 = ( a  &  d  &  (~ e)  &  wire94 ) ;
 assign wire895 = ( (~ wire15)  &  wire228  &  n_n730  &  wire255 ) ;
 assign wire898 = ( n_n1165  &  n_n1155  &  n_n700  &  n_n1146 ) ;
 assign wire900 = ( n_n1207  &  n_n904  &  wire228  &  n_n1187 ) ;
 assign wire901 = ( n_n1207  &  wire29  &  wire228  &  n_n1187 ) ;
 assign wire902 = ( n_n1207  &  wire228  &  n_n1187  &  n_n698 ) ;
 assign wire5422 = ( m  &  (~ n)  &  n_n996 ) ;
 assign wire903 = ( wire371  &  wire5422 ) | ( wire80  &  wire5422 ) | ( wire414  &  wire5422 ) ;
 assign wire904 = ( n_n1177  &  n_n1155  &  wire210  &  n_n1146 ) ;
 assign wire906 = ( n_n1177  &  n_n821  &  wire30  &  n_n1146 ) ;
 assign wire907 = ( n_n711  &  n_n1177  &  n_n821  &  n_n1146 ) ;
 assign wire908 = ( n_n1177  &  n_n1155  &  n_n1171  &  n_n1146 ) ;
 assign wire909 = ( n_n918  &  n_n1187  &  n_n996  &  n_n857 ) ;
 assign wire911 = ( wire25  &  n_n1187  &  wire380 ) | ( wire32  &  n_n1187  &  wire380 ) ;
 assign wire912 = ( wire54  &  n_n1155  &  wire219 ) | ( wire54  &  n_n1155  &  wire1016 ) ;
 assign wire914 = ( wire41  &  wire228 ) | ( n_n1161  &  n_n904  &  wire228 ) ;
 assign wire923 = ( wire58  &  n_n918  &  (~ wire137)  &  (~ n_n765) ) ;
 assign wire924 = ( n_n904  &  wire58  &  (~ n_n987)  &  (~ wire137) ) ;
 assign wire925 = ( n_n698  &  n_n694  &  wire142 ) ;
 assign wire926 = ( wire15  &  n_n1194  &  wire142 ) ;
 assign wire5313 = ( n_n904  &  n_n1194 ) | ( n_n730  &  n_n1194 ) | ( n_n904  &  wire5220 ) ;
 assign wire931 = ( n_n711  &  (~ wire30)  &  n_n982  &  wire56 ) ;
 assign wire5367 = ( (~ c)  &  d  &  (~ e)  &  l ) ;
 assign wire932 = ( n_n1202  &  n_n1137  &  wire5367 ) ;
 assign wire934 = ( n_n700  &  n_n841  &  wire260 ) ;
 assign wire935 = ( n_n1171  &  n_n1215  &  wire216 ) ;
 assign wire938 = ( n_n1171  &  n_n694  &  wire142 ) ;
 assign wire939 = ( n_n1137  &  wire47  &  n_n982 ) ;
 assign wire940 = ( wire30  &  n_n818  &  n_n982 ) ;
 assign wire941 = ( n_n709  &  n_n978  &  n_n1084 ) ;
 assign wire942 = ( n_n840  &  n_n978  &  n_n1022 ) ;
 assign wire943 = ( n_n698  &  n_n1215  &  wire216 ) ;
 assign wire945 = ( n_n978  &  n_n1094  &  n_n703 ) ;
 assign wire948 = ( n_n671  &  n_n618  &  n_n1216 ) ;
 assign wire952 = ( n_n1171  &  n_n841  &  n_n978 ) ;
 assign wire960 = ( wire34  &  n_n1204 ) | ( n_n1204  &  wire35 ) ;
 assign wire961 = ( c  &  f  &  (~ g)  &  _7862 ) ;
 assign wire962 = ( g  &  (~ h)  &  wire228  &  n_n1171 ) ;
 assign wire965 = ( n_n709  &  wire76  &  n_n662 ) ;
 assign wire966 = ( n_n840  &  wire76  &  n_n1095 ) ;
 assign wire967 = ( wire76  &  n_n841  &  n_n1053 ) ;
 assign wire968 = ( n_n841  &  n_n978  &  wire47 ) ;
 assign wire969 = ( n_n709  &  n_n978  &  n_n662 ) ;
 assign wire970 = ( n_n1137  &  n_n1053  &  n_n982 ) ;
 assign wire971 = ( n_n978  &  n_n820  &  n_n1053 ) ;
 assign wire972 = ( n_n671  &  n_n978  &  n_n670 ) ;
 assign wire973 = ( n_n840  &  n_n978  &  n_n1095 ) ;
 assign wire974 = ( n_n711  &  n_n978  &  n_n1094 ) ;
 assign wire975 = ( n_n841  &  n_n978  &  n_n1053 ) ;
 assign wire976 = ( n_n978  &  n_n838  &  n_n1094 ) ;
 assign wire977 = ( _624 ) | ( n_n1171  &  wire76  &  n_n841 ) ;
 assign wire978 = ( wire58  &  n_n730  &  n_n765 ) ;
 assign wire5309 = ( j  &  k  &  m  &  (~ n) ) ;
 assign wire982 = ( wire15  &  n_n1194  &  wire5309 ) ;
 assign wire983 = ( n_n1201  &  wire15  &  wire265 ) ;
 assign wire985 = ( n_n1217  &  n_n1220  &  n_n698  &  n_n841 ) ;
 assign wire5314 = ( j  &  k  &  m  &  (~ n) ) ;
 assign wire986 = ( wire106  &  wire5314 ) | ( wire50  &  wire5314 ) | ( wire5313  &  wire5314 ) ;
 assign wire5317 = ( i  &  wire58 ) ;
 assign wire989 = ( wire41  &  wire5317 ) | ( wire1012  &  wire5317 ) | ( wire299  &  wire5317 ) ;
 assign wire5318 = ( i  &  j  &  k  &  _7798 ) ;
 assign wire990 = ( wire41  &  wire5318 ) | ( wire1012  &  wire5318 ) | ( wire299  &  wire5318 ) ;
 assign wire991 = ( n_n918  &  wire228  &  n_n861 ) | ( n_n918  &  wire265  &  n_n861 ) ;
 assign wire992 = ( n_n1193  &  wire15  &  wire228 ) | ( n_n1193  &  wire15  &  wire265 ) ;
 assign wire993 = ( n_n920  &  n_n1193  &  wire228 ) | ( n_n920  &  n_n1193  &  wire265 ) ;
 assign wire994 = ( wire265  &  n_n698  &  n_n1137 ) ;
 assign wire995 = ( wire265  &  wire25  &  n_n1187 ) | ( wire265  &  wire32  &  n_n1187 ) ;
 assign wire5289 = ( n_n876  &  n_n864 ) | ( n_n1193  &  wire16 ) ;
 assign wire997 = ( wire228  &  wire5289 ) | ( wire228  &  n_n861  &  wire14 ) ;
 assign wire1039 = ( (~ m)  &  (~ n)  &  wire34 ) | ( (~ m)  &  (~ n)  &  wire35 ) ;
 assign wire5270 = ( (~ m)  &  n  &  n_n671 ) | ( (~ m)  &  n  &  n_n623 ) ;
 assign wire5271 = ( j  &  k  &  (~ m)  &  n ) ;
 assign wire1018 = ( wire59  &  wire1039  &  wire5271 ) | ( wire59  &  wire5270  &  wire5271 ) ;
 assign wire5274 = ( j  &  k  &  (~ m)  &  n ) ;
 assign wire1019 = ( wire23  &  wire47  &  wire5274 ) | ( wire23  &  wire60  &  wire5274 ) ;
 assign wire5277 = ( (~ f)  &  (~ g)  &  (~ h)  &  i ) | ( (~ f)  &  (~ g)  &  h  &  (~ i) ) ;
 assign wire1020 = ( n_n1210  &  wire5277  &  _7751 ) ;
 assign wire5279 = ( j  &  k  &  (~ m)  &  n ) ;
 assign wire1021 = ( n_n711  &  wire134  &  wire5279 ) | ( wire30  &  wire134  &  wire5279 ) ;
 assign wire1022 = ( n_n1191  &  wire23  &  _7757 ) ;
 assign wire1023 = ( n_n1036  &  n_n1137  &  wire47 ) | ( n_n1036  &  n_n1137  &  wire60 ) ;
 assign wire1024 = ( n_n1210  &  wire59  &  _7759 ) ;
 assign wire1027 = ( n_n711  &  n_n1036  &  n_n818 ) | ( wire30  &  n_n1036  &  n_n818 ) ;
 assign wire1030 = ( n_n700  &  n_n1202  &  n_n1137 ) ;
 assign wire1031 = ( wire34  &  n_n1191  &  wire398 ) | ( n_n1191  &  wire398  &  wire35 ) ;
 assign wire1032 = ( wire34  &  n_n1191  &  n_n670 ) | ( n_n1191  &  n_n670  &  wire35 ) ;
 assign wire1033 = ( wire265  &  n_n1171  &  n_n1137 ) ;
 assign wire1034 = ( wire265  &  wire5289 ) | ( wire265  &  n_n861  &  wire14 ) ;
 assign wire1036 = ( n_n617  &  wire1039 ) | ( n_n617  &  wire5270 ) ;
 assign wire5246 = ( (~ f)  &  h  &  (~ m)  &  (~ n) ) ;
 assign wire1051 = ( n_n1229  &  wire65  &  wire5246 ) | ( n_n1229  &  n_n235  &  wire5246 ) ;
 assign wire1052 = ( n_n1165  &  wire65  &  (~ wire232) ) | ( n_n1165  &  (~ wire232)  &  n_n235 ) ;
 assign wire1053 = ( n_n1165  &  n_n1101  &  wire65 ) | ( n_n1165  &  n_n1101  &  n_n235 ) ;
 assign wire1054 = ( n_n1177  &  n_n671  &  wire65 ) | ( n_n1177  &  n_n671  &  n_n235 ) ;
 assign wire5220 = ( (~ e)  &  (~ g)  &  h ) ;
 assign wire1055 = ( n_n904  &  wire54  &  wire5220 ) ;
 assign wire1057 = ( _763 ) | ( wire84  &  n_n1253  &  n_n1160 ) ;
 assign wire1058 = ( wire172  &  wire377 ) | ( wire172  &  wire115 ) ;
 assign wire1059 = ( n_n904  &  wire58  &  n_n765 ) ;
 assign wire5088 = ( k  &  n_n1177  &  n_n819 ) | ( (~ k)  &  n_n1177  &  n_n818 ) ;
 assign wire1060 = ( n_n626  &  wire5088 ) | ( n_n626  &  n_n1056  &  n_n816 ) ;
 assign wire1061 = ( a  &  (~ c)  &  d  &  wire138 ) ;
 assign wire5252 = ( f  &  g  &  (~ h)  &  (~ n) ) ;
 assign wire1062 = ( n_n904  &  wire5253 ) | ( n_n904  &  n_n874  &  wire5252 ) ;
 assign wire5213 = ( (~ a)  &  b  &  d ) ;
 assign wire1070 = ( n_n1220  &  n_n1082  &  wire5213 ) ;
 assign wire1071 = ( n_n1166  &  n_n973  &  n_n1204  &  n_n1095 ) ;
 assign wire1074 = ( n_n626  &  n_n1210  &  wire134 ) ;
 assign wire1075 = ( n_n626  &  wire76  &  n_n1094 ) ;
 assign wire1076 = ( n_n973  &  n_n1095  &  n_n1191 ) ;
 assign wire1077 = ( n_n1229  &  n_n1166  &  n_n1204  &  n_n662 ) ;
 assign wire1078 = ( n_n1229  &  n_n662  &  n_n1191 ) ;
 assign wire1079 = ( n_n904  &  n_n1220  &  wire5220 ) ;
 assign wire1080 = ( n_n1101  &  n_n1166  &  n_n1204 ) ;
 assign wire1081 = ( n_n671  &  n_n1166  &  n_n1216 ) ;
 assign wire1082 = ( wire293  &  wire377 ) | ( wire293  &  wire115 ) ;
 assign wire1083 = ( wire77  &  wire377 ) | ( wire77  &  wire115 ) ;
 assign wire1096 = ( wire175  &  n_n918  &  n_n1187  &  n_n816 ) ;
 assign wire1100 = ( n_n949  &  n_n816  &  _7511 ) ;
 assign wire1102 = ( n_n942  &  n_n1187  &  n_n949  &  n_n912 ) ;
 assign wire1106 = ( _814 ) | ( n_n893  &  wire393  &  n_n1177 ) ;
 assign wire5140 = ( b  &  c  &  (~ d)  &  (~ h) ) ;
 assign wire1123 = ( wire224  &  wire190  &  _7467 ) ;
 assign wire5144 = ( b  &  (~ c)  &  d ) ;
 assign wire1147 = ( a  &  b  &  c  &  _7437 ) ;
 assign wire1148 = ( a  &  b  &  d  &  _7433 ) ;
 assign wire1128 = ( n_n711  &  n_n886  &  wire172 ) ;
 assign wire1129 = ( n_n709  &  n_n1188  &  wire148 ) ;
 assign wire1130 = ( n_n1089  &  n_n842  &  wire84 ) ;
 assign wire1131 = ( n_n1161  &  n_n713  &  n_n893  &  n_n1177 ) ;
 assign wire1135 = ( wire76  &  n_n1095  &  n_n1094  &  n_n703 ) ;
 assign wire1137 = ( n_n840  &  wire76  &  n_n1095 ) ;
 assign wire1198 = ( g  &  (~ i)  &  j  &  wire96 ) ;
 assign wire1200 = ( g  &  i  &  k  &  _7270 ) ;
 assign wire1138 = ( wire153  &  wire72 ) | ( wire153  &  wire1198 ) | ( wire153  &  wire1200 ) ;
 assign wire1139 = ( n_n709  &  wire72 ) | ( n_n709  &  wire1198 ) | ( n_n709  &  wire1200 ) ;
 assign wire5116 = ( n_n842  &  n_n1194 ) | ( n_n713  &  n_n1196 ) ;
 assign wire1140 = ( wire172  &  wire5116 ) | ( n_n842  &  wire172  &  n_n1201 ) ;
 assign wire1155 = ( n_n711  &  wire172  &  _7387 ) ;
 assign wire1156 = ( n_n709  &  n_n1201  &  wire293 ) ;
 assign wire1157 = ( (~ m)  &  (~ n)  &  n_n626  &  wire198 ) ;
 assign wire1158 = ( n_n709  &  wire172  &  n_n1201 ) ;
 assign wire1162 = ( n_n709  &  n_n1201  &  wire77 ) ;
 assign wire1163 = ( n_n840  &  n_n822  &  wire77 ) ;
 assign wire1166 = ( n_n1191  &  n_n628  &  n_n235 ) ;
 assign wire1167 = ( n_n1229  &  n_n662  &  n_n1191 ) ;
 assign wire1168 = ( g  &  n_n711  &  wire71  &  wire293 ) | ( (~ g)  &  n_n711  &  wire71  &  wire293 ) ;
 assign wire1169 = ( g  &  n_n711  &  wire71  &  wire77 ) | ( (~ g)  &  n_n711  &  wire71  &  wire77 ) ;
 assign wire1170 = ( m  &  (~ n)  &  n_n698  &  n_n816 ) ;
 assign wire1171 = ( n_n1229  &  n_n1190  &  n_n825 ) ;
 assign wire1172 = ( n_n713  &  n_n886  &  wire172 ) ;
 assign wire1173 = ( n_n626  &  n_n1166  &  n_n1204 ) ;
 assign wire1175 = ( wire293  &  wire5116 ) | ( n_n842  &  n_n1201  &  wire293 ) ;
 assign wire1176 = ( wire77  &  wire5116 ) | ( n_n842  &  n_n1201  &  wire77 ) ;
 assign wire1185 = ( n_n709  &  n_n1219  &  n_n825 ) ;
 assign wire1186 = ( n_n821  &  n_n1210  &  n_n703 ) ;
 assign wire1187 = ( n_n840  &  n_n1036  &  n_n823 ) ;
 assign wire1188 = ( n_n709  &  wire228  &  n_n861 ) | ( n_n709  &  wire265  &  n_n861 ) ;
 assign wire1189 = ( n_n1229  &  n_n662  &  wire260 ) ;
 assign wire1192 = ( n_n698  &  n_n1219  &  n_n1137 ) ;
 assign wire1193 = ( n_n1210  &  n_n1094  &  n_n703 ) ;
 assign wire1194 = ( n_n840  &  n_n1210  &  wire89 ) ;
 assign wire1195 = ( n_n698  &  wire72 ) | ( n_n698  &  wire1198 ) | ( n_n698  &  wire1200 ) ;
 assign wire1196 = ( _905 ) | ( wire379  &  _7308 ) ;
 assign wire1197 = ( n_n703  &  wire5088 ) | ( n_n1056  &  n_n816  &  n_n703 ) ;
 assign wire5091 = ( n_n698  &  n_n1215  &  wire23 ) | ( n_n698  &  n_n1215  &  wire105 ) ;
 assign wire5093 = ( wire1185 ) | ( wire1186 ) | ( wire1194 ) ;
 assign wire5094 = ( wire1187 ) | ( wire1189 ) | ( wire5091 ) ;
 assign wire5095 = ( wire1188 ) | ( wire1192 ) | ( wire1193 ) ;
 assign wire5108 = ( c  &  (~ e)  &  f  &  wire65 ) ;
 assign wire5117 = ( n_n709  &  n_n868  &  wire385 ) | ( n_n709  &  n_n871  &  wire385 ) ;
 assign wire5120 = ( n_n709  &  wire54  &  n_n971 ) | ( n_n709  &  n_n1220  &  n_n971 ) ;
 assign wire5125 = ( wire1156 ) | ( n_n1229  &  wire71  &  wire162 ) ;
 assign wire5126 = ( wire1168 ) | ( wire1169 ) ;
 assign wire5127 = ( wire1157 ) | ( wire1158 ) | ( wire5117 ) ;
 assign wire5128 = ( wire1162 ) | ( wire1163 ) | ( wire5120 ) ;
 assign wire5129 = ( wire1166 ) | ( wire1167 ) | ( wire1170 ) | ( wire1171 ) ;
 assign wire5130 = ( wire1172 ) | ( wire1173 ) | ( wire162  &  wire5108 ) ;
 assign wire5136 = ( wire1175 ) | ( wire1176 ) | ( _7390 ) ;
 assign wire5137 = ( wire5125 ) | ( wire5126 ) | ( wire5127 ) | ( wire5128 ) ;
 assign wire5146 = ( wire202  &  wire76  &  n_n1095 ) ;
 assign wire5156 = ( a  &  b  &  (~ c)  &  _7503 ) ;
 assign wire5159 = ( wire1123 ) | ( wire84  &  wire5140  &  _7462 ) ;
 assign wire5160 = ( _843 ) | ( wire76  &  n_n1095  &  wire5144 ) ;
 assign wire5161 = ( wire84  &  wire393 ) | ( n_n893  &  wire393  &  n_n1177 ) ;
 assign wire5162 = ( wire1135 ) | ( (~ g)  &  wire153  &  wire190 ) ;
 assign wire5163 = ( wire1128 ) | ( wire1129 ) | ( wire1137 ) ;
 assign wire5169 = ( _7453 ) | ( wire46  &  wire1147 ) | ( wire46  &  wire1148 ) ;
 assign wire5170 = ( wire1140 ) | ( wire5159 ) | ( wire5160 ) | ( wire5161 ) ;
 assign wire5171 = ( wire1138 ) | ( wire5162 ) | ( wire5163 ) ;
 assign wire5172 = ( wire1139 ) | ( wire46  &  wire5146 ) | ( wire46  &  wire5156 ) ;
 assign wire5176 = ( _803 ) | ( _804 ) ;
 assign wire5177 = ( m  &  (~ n)  &  n_n918  &  wire105 ) ;
 assign wire5179 = ( (~ m)  &  n  &  n_n713  &  n_n1231 ) ;
 assign wire5181 = ( n_n713  &  n_n893  &  n_n1177  &  n_n1231 ) ;
 assign wire5183 = ( a  &  (~ b)  &  c  &  _7524 ) ;
 assign wire5184 = ( (~ a)  &  b  &  d  &  e ) ;
 assign wire5187 = ( a  &  (~ b)  &  c  &  _7556 ) ;
 assign wire5188 = ( (~ a)  &  b  &  d  &  e ) ;
 assign wire5190 = ( m  &  (~ n)  &  n_n949  &  n_n1231 ) ;
 assign wire5191 = ( a  &  (~ b)  &  c  &  _7569 ) ;
 assign wire5192 = ( (~ a)  &  b  &  d  &  e ) ;
 assign wire5194 = ( m  &  (~ n)  &  n_n949  &  n_n1231 ) ;
 assign wire5197 = ( wire5176  &  wire5177 ) | ( wire20  &  wire5181 ) ;
 assign wire5198 = ( wire1096 ) | ( n_n1187  &  n_n949  &  wire108 ) ;
 assign wire5199 = ( wire1100 ) | ( wire1102 ) | ( wire101  &  wire5179 ) ;
 assign wire5201 = ( wire181  &  wire388 ) | ( wire152  &  wire5190 ) ;
 assign wire5204 = ( wire1112  &  wire5187 ) | ( wire1113  &  wire5187 ) | ( wire1112  &  wire5188 ) | ( wire1113  &  wire5188 ) ;
 assign wire5205 = ( wire69  &  wire5191 ) | ( wire1116  &  wire5191 ) | ( wire69  &  wire5192 ) | ( wire1116  &  wire5192 ) ;
 assign wire5215 = ( a  &  (~ c)  &  d  &  (~ e) ) ;
 assign wire5216 = ( (~ a)  &  b  &  d  &  e ) ;
 assign wire5226 = ( n_n1219  &  wire121  &  wire5215 ) | ( n_n1219  &  wire121  &  wire5216 ) ;
 assign wire5227 = ( wire1070 ) | ( wire1071 ) | ( wire1074 ) | ( wire1075 ) ;
 assign wire5228 = ( wire1076 ) | ( wire1077 ) | ( wire1078 ) | ( wire1079 ) ;
 assign wire5232 = ( wire1080 ) | ( wire1081 ) | ( wire1082 ) | ( wire5228 ) ;
 assign wire5233 = ( wire1083 ) | ( wire5227 ) | ( _7649 ) ;
 assign wire5237 = ( n_n904  &  (~ wire22)  &  _7662 ) ;
 assign wire5238 = ( a  &  (~ c)  &  d  &  (~ n) ) ;
 assign wire5241 = ( n_n1193  &  (~ wire22)  &  wire5238 ) ;
 assign wire5243 = ( m  &  (~ n)  &  n_n904  &  _7671 ) ;
 assign wire5244 = ( (~ f)  &  h  &  wire54 ) ;
 assign wire5251 = ( f  &  g  &  h  &  (~ n) ) ;
 assign wire5255 = ( wire31  &  (~ wire54)  &  wire5237 ) | ( wire31  &  (~ wire54)  &  wire5241 ) ;
 assign wire5256 = ( wire45  &  wire258 ) | ( wire31  &  wire258  &  wire5244 ) ;
 assign wire5257 = ( wire1055 ) | ( wire1059 ) | ( wire101  &  wire5243 ) ;
 assign wire5266 = ( wire1062 ) | ( wire5255 ) | ( wire5256 ) | ( wire5257 ) ;
 assign wire5290 = ( n_n1171  &  n_n529  &  wire96 ) | ( n_n698  &  n_n529  &  wire96 ) ;
 assign wire5291 = ( n_n1220  &  n_n1171  &  n_n818 ) | ( n_n1220  &  n_n698  &  n_n818 ) ;
 assign wire5293 = ( wire58  &  n_n1171  &  n_n841 ) | ( wire58  &  n_n698  &  n_n841 ) ;
 assign wire5297 = ( wire1030 ) | ( wire1033 ) | ( wire5291 ) ;
 assign wire5298 = ( wire1019 ) | ( wire5293 ) ;
 assign wire5299 = ( wire1023 ) | ( _679 ) | ( _680 ) ;
 assign wire5300 = ( wire1020 ) | ( wire1021 ) | ( wire1022 ) | ( wire1024 ) ;
 assign wire5316 = ( i  &  j  &  k  &  _7815 ) ;
 assign wire5321 = ( wire985 ) | ( wire994 ) | ( _670 ) ;
 assign wire5323 = ( wire993 ) | ( _665 ) | ( _666 ) ;
 assign wire5325 = ( wire98  &  wire5316 ) | ( i  &  wire58  &  wire98 ) ;
 assign wire5327 = ( wire982 ) | ( wire983 ) | ( wire5321 ) | ( wire5323 ) ;
 assign wire5328 = ( wire986 ) | ( wire989 ) ;
 assign wire5329 = ( wire990 ) | ( wire995 ) ;
 assign wire5330 = ( wire991 ) | ( wire992 ) | ( wire997 ) | ( wire5325 ) ;
 assign wire5356 = ( _621 ) | ( wire58  &  wire14  &  _7833 ) ;
 assign wire5357 = ( n_n2660 ) | ( wire962 ) | ( wire968 ) ;
 assign wire5358 = ( wire965 ) | ( wire966 ) | ( wire967 ) | ( wire969 ) ;
 assign wire5359 = ( wire970 ) | ( wire971 ) | ( wire972 ) | ( wire973 ) ;
 assign wire5360 = ( wire974 ) | ( wire975 ) | ( wire976 ) | ( wire978 ) ;
 assign wire5364 = ( wire5356 ) | ( wire5357 ) | ( wire5358 ) | ( wire5359 ) ;
 assign wire5368 = ( k  &  (~ m)  &  n_n670 ) ;
 assign wire5379 = ( n_n700  &  n_n841  &  wire188 ) | ( n_n700  &  wire188  &  n_n820 ) ;
 assign wire5382 = ( n_n671  &  n_n1166  &  n_n1216 ) | ( n_n671  &  n_n1216  &  wire56 ) ;
 assign wire5386 = ( wire932 ) | ( wire934 ) | ( wire943 ) ;
 assign wire5387 = ( wire938 ) | ( wire941 ) | ( wire5379 ) ;
 assign wire5388 = ( wire942 ) | ( wire945 ) | ( wire5382 ) ;
 assign wire5389 = ( wire948 ) | ( wire952 ) | ( wire380  &  wire208 ) ;
 assign wire5391 = ( wire931 ) | ( wire935 ) | ( wire939 ) | ( wire940 ) ;
 assign wire5395 = ( wire5386 ) | ( wire5387 ) | ( wire5391 ) ;
 assign wire5396 = ( n_n1166  &  wire960 ) | ( n_n1166  &  wire961 ) | ( wire960  &  wire5368 ) | ( wire961  &  wire5368 ) ;
 assign wire5397 = ( wire5388 ) | ( _589 ) | ( _594 ) | ( _595 ) ;
 assign wire5413 = ( f  &  h  &  (~ i)  &  wire30 ) ;
 assign wire5414 = ( (~ m)  &  n  &  wire34  &  n_n1146 ) ;
 assign wire5415 = ( _559 ) | ( _560 ) | ( _561 ) ;
 assign wire5416 = ( (~ m)  &  n  &  n_n824  &  n_n1146 ) ;
 assign wire5418 = ( (~ m)  &  n  &  n_n933  &  n_n1146 ) ;
 assign wire5424 = ( m  &  (~ n)  &  wire29 ) ;
 assign wire5431 = ( wire895 ) | ( wire54  &  n_n1155  &  n_n698 ) ;
 assign wire5432 = ( wire5415  &  wire5416 ) | ( wire309  &  wire5418 ) ;
 assign wire5433 = ( wire900 ) | ( wire901 ) ;
 assign wire5435 = ( wire906 ) | ( wire54  &  n_n1155  &  wire291 ) ;
 assign wire5436 = ( wire898 ) | ( wire907 ) | ( wire908 ) | ( wire909 ) ;
 assign wire5437 = ( wire5413  &  wire5414 ) | ( wire179  &  wire5424 ) ;
 assign wire5443 = ( wire912 ) | ( wire5431 ) | ( wire5432 ) | ( wire5433 ) ;
 assign wire5444 = ( wire902 ) | ( wire904 ) | ( wire911 ) | ( wire5435 ) ;
 assign wire5446 = ( wire903 ) | ( wire914 ) | ( wire5436 ) | ( wire5437 ) ;
 assign wire5451 = ( (~ c)  &  e ) | ( (~ d)  &  e ) ;
 assign wire5453 = ( n_n1166  &  n_n1204  &  wire5451 ) ;
 assign wire5456 = ( (~ b)  &  c  &  e ) ;
 assign wire5457 = ( n_n709  &  wire71  &  wire77 ) | ( n_n709  &  wire71  &  wire227 ) ;
 assign wire5459 = ( wire884 ) | ( (~ n_n1069)  &  n_n1095  &  wire5453 ) ;
 assign wire5460 = ( _513 ) | ( n_n1210  &  wire89  &  wire5454 ) ;
 assign wire5461 = ( wire879 ) | ( wire880 ) | ( wire5457 ) ;
 assign wire5462 = ( wire184  &  wire77 ) | ( wire117  &  wire5456 ) ;
 assign wire5463 = ( n_n709  &  wire135 ) | ( wire94  &  wire43 ) ;
 assign wire5467 = ( wire886 ) | ( wire5459 ) | ( wire5460 ) | ( wire5461 ) ;
 assign wire5469 = ( a  &  (~ b)  &  d  &  f ) ;
 assign wire5477 = ( b  &  (~ c) ) | ( b  &  (~ e) ) | ( (~ c)  &  (~ f) ) | ( (~ e)  &  (~ f) ) ;
 assign wire5479 = ( (~ n_n709)  &  wire229  &  wire5477 ) ;
 assign wire5485 = ( wire229  &  n_n1165  &  (~ n_n1229)  &  (~ n_n1069) ) ;
 assign wire5489 = ( _493 ) | ( _494 ) ;
 assign wire5490 = ( (~ m)  &  n  &  n_n893  &  n_n1166 ) ;
 assign wire5493 = ( (~ m)  &  n  &  n_n842  &  wire229 ) ;
 assign wire5495 = ( a  &  m  &  (~ n)  &  _8084 ) ;
 assign wire5505 = ( wire854 ) | ( wire76  &  n_n1095  &  wire5479 ) ;
 assign wire5507 = ( wire84  &  wire393 ) | ( n_n893  &  wire393  &  n_n1177 ) ;
 assign wire5508 = ( wire65  &  wire5485 ) | ( n_n235  &  wire5485 ) | ( wire65  &  wire5493 ) | ( n_n235  &  wire5493 ) ;
 assign wire5509 = ( wire853 ) | ( n  &  wire184  &  wire49 ) ;
 assign wire5513 = ( wire46  &  wire5495 ) | ( wire46  &  wire5489  &  wire5490 ) ;
 assign wire5515 = ( wire859 ) | ( n_n920  &  n_n1187  &  wire92 ) ;
 assign wire5517 = ( wire5505 ) | ( wire5507 ) | ( _8076 ) ;
 assign wire5520 = ( wire5508 ) | ( wire5509 ) | ( wire5515 ) ;
 assign wire5561 = ( n_n1220  &  n_n1171  &  wire206 ) | ( n_n1220  &  n_n698  &  wire206 ) ;
 assign wire5570 = ( n_n820  &  n_n1191  &  wire109 ) | ( n_n1191  &  wire23  &  wire109 ) ;
 assign wire5572 = ( wire809 ) | ( wire810 ) | ( wire811 ) | ( wire813 ) ;
 assign wire5573 = ( wire814 ) | ( wire817 ) | ( wire5561 ) ;
 assign wire5574 = ( wire821 ) | ( wire822 ) | ( wire826 ) | ( wire827 ) ;
 assign wire5575 = ( wire828 ) | ( wire829 ) | ( wire830 ) | ( wire831 ) ;
 assign wire5576 = ( wire823 ) | ( wire832 ) | ( wire835 ) ;
 assign wire5578 = ( wire808 ) | ( wire812 ) | ( wire815 ) | ( wire837 ) ;
 assign wire5579 = ( wire816 ) | ( wire818 ) | ( wire5570 ) ;
 assign wire5602 = ( i  &  k  &  m  &  (~ n) ) ;
 assign wire5603 = ( i  &  k  &  m  &  (~ n) ) ;
 assign wire5605 = ( (~ i)  &  wire148 ) | ( (~ j)  &  wire148 ) ;
 assign wire5611 = ( wire106  &  wire5602 ) | ( n_n893  &  wire148  &  wire106 ) ;
 assign wire5613 = ( wire148  &  wire156 ) | ( wire33  &  wire203 ) ;
 assign wire5615 = ( wire784 ) | ( wire786 ) | ( wire787 ) | ( wire788 ) ;
 assign wire5618 = ( wire50  &  wire5603 ) | ( wire5313  &  wire5603 ) | ( wire50  &  wire5605 ) | ( wire5313  &  wire5605 ) ;
 assign wire5621 = ( wire790 ) | ( wire796 ) | ( wire797 ) | ( wire5613 ) ;
 assign wire5637 = ( d  &  (~ e)  &  f ) ;
 assign wire5652 = ( n_n2507 ) | ( wire775 ) | ( wire776 ) | ( wire766 ) ;
 assign wire5677 = ( c  &  d  &  wire120  &  n_n1231 ) ;
 assign wire5678 = ( c  &  d  &  (~ f) ) ;
 assign wire5679 = ( m  &  (~ n)  &  n_n1261  &  wire5678 ) ;
 assign wire5681 = ( c  &  d  &  wire120  &  n_n912 ) ;
 assign wire5693 = ( n_n1220  &  wire120  &  (~ wire57)  &  n_n1082 ) ;
 assign wire5695 = ( c  &  d  &  wire120 ) ;
 assign wire5703 = ( (~ a)  &  b  &  c  &  e ) ;
 assign wire5704 = ( a  &  c  &  (~ d)  &  e ) ;
 assign wire5705 = ( (~ a)  &  b  &  c  &  (~ d) ) ;
 assign wire5708 = ( n_n2660 ) | ( wire736 ) | ( wire108  &  wire5705 ) ;
 assign wire5709 = ( wire718 ) | ( wire719 ) | ( wire724 ) | ( wire726 ) ;
 assign wire5710 = ( wire200  &  wire5693 ) | ( wire379  &  wire5703 ) ;
 assign wire5711 = ( wire138  &  n_n949 ) | ( wire138  &  wire5704 ) ;
 assign wire5715 = ( n_n997  &  wire1112 ) | ( wire413  &  wire1112 ) | ( n_n997  &  wire1113 ) | ( wire413  &  wire1113 ) ;
 assign wire5718 = ( wire5708 ) | ( wire5711 ) | ( n_n949  &  wire94 ) ;
 assign wire5719 = ( wire725 ) | ( _378 ) | ( _379 ) ;
 assign wire5720 = ( wire713 ) | ( wire727 ) | ( wire5709 ) ;
 assign wire5721 = ( wire5715 ) | ( _8394 ) ;
 assign wire5727 = ( a  &  b  &  d  &  _8487 ) ;
 assign wire5744 = ( (~ b)  &  c  &  d  &  _8427 ) ;
 assign wire5758 = ( n_n840  &  wire76  &  n_n1095 ) | ( wire76  &  n_n988  &  n_n1095 ) ;
 assign wire5759 = ( wire228  &  wire159 ) | ( wire22  &  wire159  &  wire197 ) ;
 assign wire5760 = ( n_n2572 ) | ( wire680 ) | ( wire84  &  wire167 ) ;
 assign wire5761 = ( wire681 ) | ( wire682 ) | ( wire683 ) | ( wire684 ) ;
 assign wire5762 = ( n  &  wire160  &  wire49 ) | ( n  &  wire49  &  wire5744 ) ;
 assign wire5763 = ( n_n2660 ) | ( wire679 ) | ( wire736 ) | ( wire5758 ) ;
 assign wire5766 = ( wire5759 ) | ( wire5760 ) | ( wire5763 ) ;
 assign wire5792 = ( wire265  &  wire159 ) | ( wire75  &  wire167 ) ;
 assign wire5793 = ( wire643 ) | ( wire645 ) | ( wire77  &  wire160 ) ;
 assign wire5795 = ( wire649 ) | ( n_n838  &  (~ n_n1252)  &  wire117 ) ;
 assign wire5797 = ( n_n988  &  wire117 ) | ( n_n842  &  wire135 ) ;
 assign wire5798 = ( wire644 ) | ( wire647 ) | ( wire651 ) | ( wire652 ) ;
 assign wire5806 = ( wire655 ) | ( wire663 ) | ( _8474 ) ;
 assign wire5824 = ( wire626 ) | ( wire629 ) | ( wire630 ) | ( wire633 ) ;
 assign wire5825 = ( wire627 ) | ( n_n698  &  wire72 ) ;
 assign wire5826 = ( wire628 ) | ( wire631 ) | ( wire632 ) | ( wire635 ) ;
 assign wire5831 = ( wire54  &  n_n1155 ) | ( n_n529  &  wire142 ) ;
 assign wire5833 = ( (~ n_n1193)  &  (~ n_n1201)  &  n_n918  &  n_n1187 ) ;
 assign wire5835 = ( m  &  (~ n)  &  n_n1207  &  wire29 ) ;
 assign wire5836 = ( m  &  (~ n)  &  n_n1201  &  wire29 ) ;
 assign wire5837 = ( i  &  k  &  m  &  (~ n) ) ;
 assign wire5842 = ( wire610 ) | ( wire156  &  wire5837 ) ;
 assign wire5846 = ( wire81  &  wire5833 ) | ( wire5831  &  wire5833 ) | ( wire81  &  wire5835 ) | ( wire5831  &  wire5835 ) ;
 assign wire5847 = ( n_n698  &  wire81 ) | ( n_n698  &  wire5831 ) | ( wire81  &  wire5836 ) | ( wire5831  &  wire5836 ) ;
 assign wire5858 = ( (~ k)  &  (~ m)  &  (~ n)  &  _8619 ) ;
 assign wire5860 = ( n_n1155  &  n_n700  &  n_n1191 ) | ( n_n700  &  n_n820  &  n_n1191 ) ;
 assign wire5864 = ( wire594 ) | ( wire113  &  wire203 ) ;
 assign wire5865 = ( wire587 ) | ( wire588 ) | ( wire5860 ) ;
 assign wire5866 = ( wire593 ) | ( wire598 ) | ( n_n1210  &  wire208 ) ;
 assign wire5867 = ( n_n3060 ) | ( wire585 ) | ( wire586 ) | ( wire590 ) ;
 assign wire5870 = ( wire5864 ) | ( wire5865 ) | ( wire5867 ) ;
 assign wire5871 = ( wire40  &  wire1039 ) | ( wire40  &  wire5270 ) | ( wire1039  &  wire5858 ) | ( wire5270  &  wire5858 ) ;
 assign wire5875 = ( h  &  i  &  (~ j)  &  k ) ;
 assign wire5876 = ( (~ wire104)  &  wire5875 ) ;
 assign wire5877 = ( n_n711  &  wire293 ) | ( wire30  &  wire293 ) ;
 assign wire5888 = ( (~ h)  &  (~ k) ) | ( j  &  (~ k) ) ;
 assign wire5897 = ( n_n2953 ) | ( wire567 ) | ( wire575 ) ;
 assign wire5898 = ( wire568 ) | ( wire576 ) | ( wire5876  &  wire5877 ) ;
 assign wire5899 = ( wire571 ) | ( _217 ) | ( _218 ) ;
 assign wire5901 = ( wire565 ) | ( wire566 ) | ( wire569 ) | ( wire577 ) ;
 assign wire5925 = ( wire540 ) | ( _202 ) | ( _203 ) ;
 assign wire5927 = ( wire536 ) | ( wire539 ) | ( wire541 ) | ( wire542 ) ;
 assign wire5928 = ( wire543 ) | ( wire544 ) | ( wire545 ) | ( wire549 ) ;
 assign wire5929 = ( wire550 ) | ( wire551 ) | ( n_n1264  &  wire209 ) ;
 assign wire5930 = ( wire537 ) | ( wire554 ) | ( n_n1220  &  wire50 ) ;
 assign wire5934 = ( wire548 ) | ( _182 ) | ( _183 ) ;
 assign wire5943 = ( e  &  (~ f)  &  m  &  (~ n) ) ;
 assign wire5944 = ( (~ c)  &  d  &  (~ g)  &  (~ h) ) ;
 assign wire5945 = ( c  &  (~ f)  &  (~ h)  &  i ) ;
 assign wire5951 = ( wire282  &  wire5944 ) | ( wire282  &  wire5945 ) ;
 assign wire5954 = ( wire528 ) | ( wire5951 ) | ( wire373  &  wire5943 ) ;
 assign wire5955 = ( wire532 ) | ( wire533 ) | ( wire534 ) | ( wire535 ) ;
 assign wire5961 = ( b  &  (~ f)  &  (~ h)  &  i ) ;
 assign wire5962 = ( (~ b)  &  (~ e)  &  g  &  (~ h) ) ;
 assign wire5963 = ( b  &  e  &  (~ f)  &  (~ h) ) ;
 assign wire5967 = ( wire227  &  wire5961 ) | ( wire227  &  wire5962 ) ;
 assign wire5969 = ( wire520 ) | ( wire521 ) | ( wire522 ) | ( wire523 ) ;
 assign wire5970 = ( wire527 ) | ( wire5967 ) | ( wire227  &  wire5963 ) ;
 assign wire5981 = ( (~ i)  &  (~ k)  &  m  &  (~ n) ) ;
 assign wire5982 = ( f  &  k  &  m  &  (~ n) ) ;
 assign wire5986 = ( wire22  &  wire283 ) | ( n_n1171  &  wire286 ) ;
 assign wire5990 = ( n_n1187  &  n_n1189  &  wire5981 ) | ( n_n1187  &  n_n1189  &  wire5982 ) ;
 assign wire5998 = ( wire508 ) | ( wire509 ) | ( wire510 ) | ( wire512 ) ;
 assign wire5999 = ( wire499 ) | ( wire513 ) | ( wire516 ) | ( wire5986 ) ;
 assign wire6035 = ( wire481 ) | ( wire483 ) | ( wire487 ) ;
 assign wire6036 = ( wire484 ) | ( wire488 ) | ( wire489 ) | ( wire490 ) ;
 assign wire6037 = ( wire491 ) | ( wire492 ) | ( wire493 ) | ( wire494 ) ;
 assign wire6038 = ( wire480 ) | ( wire482 ) | ( wire495 ) | ( wire496 ) ;
 assign wire6041 = ( wire485 ) | ( wire486 ) | ( wire6035 ) | ( wire6038 ) ;
 assign wire6045 = ( f  &  (~ i)  &  k  &  (~ m) ) ;
 assign wire6057 = ( n_n1095  &  n_n1227 ) | ( n_n1203  &  wire226 ) ;
 assign wire6062 = ( wire70  &  n_n1160 ) | ( n_n1161  &  wire285 ) ;
 assign wire6064 = ( _70 ) | ( n_n1227  &  (~ n_n1091)  &  _8998 ) ;
 assign wire6065 = ( wire463 ) | ( wire465 ) | ( wire466 ) | ( wire467 ) ;
 assign wire6066 = ( wire469 ) | ( _9021 ) | ( wire254  &  wire6054 ) ;
 assign wire6067 = ( wire461 ) | ( wire6057 ) | ( wire6062 ) ;
 assign wire6070 = ( wire6064 ) | ( wire6065 ) | ( wire6066 ) | ( wire6067 ) ;
 assign wire6071 = ( wire5999 ) | ( wire6041 ) | ( _9076 ) | ( _9128 ) ;
 assign wire6100 = ( wire443 ) | ( wire444 ) | ( wire445 ) | ( wire447 ) ;
 assign wire6101 = ( wire448 ) | ( wire449 ) | ( wire450 ) | ( wire451 ) ;
 assign wire6102 = ( wire452 ) | ( wire453 ) | ( wire454 ) | ( wire455 ) ;
 assign wire6103 = ( wire456 ) | ( wire457 ) | ( wire458 ) | ( wire460 ) ;
 assign wire6106 = ( wire446 ) | ( wire459 ) | ( wire6100 ) | ( wire6103 ) ;
 assign wire6123 = ( (~ b)  &  g  &  h ) ;
 assign wire6125 = ( m ) | ( (~ i)  &  k ) | ( (~ i)  &  l ) | ( (~ k)  &  l ) ;
 assign wire6132 = ( wire435 ) | ( _119 ) | ( _120 ) ;
 assign wire6133 = ( wire248  &  wire6125 ) | ( wire37  &  (~ n_n1216)  &  wire248 ) ;
 assign wire6135 = ( wire431 ) | ( wire432 ) | ( wire433 ) | ( wire434 ) ;
 assign wire6138 = ( wire429 ) | ( wire430 ) | ( wire442 ) | ( wire6135 ) ;
 assign wire6139 = ( wire6132 ) | ( wire6133 ) | ( _8890 ) ;
 assign wire6141 = ( (~ h)  &  i  &  (~ k) ) | ( (~ h)  &  (~ j)  &  (~ k) ) ;
 assign wire6142 = ( (~ h)  &  i  &  (~ k) ) ;
 assign wire6143 = ( (~ h)  &  i  &  (~ k) ) ;
 assign wire6144 = ( (~ i)  &  (~ m)  &  n ) ;
 assign wire6145 = ( n_n1190  &  wire6143 ) | ( n_n1160  &  wire6144 ) ;
 assign wire6147 = ( n_n1056  &  wire6141 ) | ( n_n1219  &  wire6142 ) ;
 assign wire6156 = ( c  &  (~ m)  &  n ) | ( d  &  (~ m)  &  n ) ;
 assign wire6158 = ( g  &  (~ m)  &  n ) ;
 assign wire6159 = ( n_n1091  &  wire6156 ) | ( n_n1080  &  wire6158 ) ;
 assign wire6160 = ( wire114  &  wire404 ) | ( n_n1190  &  wire305 ) ;
 assign wire6161 = ( n_n1080  &  (~ wire204) ) | ( wire286  &  wire137 ) ;
 assign wire6165 = ( k  &  n_n1177  &  n_n1028 ) | ( n_n1177  &  n_n1072  &  n_n1028 ) ;
 assign wire6176 = ( (~ n_n671)  &  (~ n_n700)  &  (~ n_n1260) ) ;
 assign wire6183 = ( (~ b)  &  (~ m)  &  n  &  wire286 ) ;
 assign wire6184 = ( _36 ) | ( _37 ) | ( _38 ) ;
 assign wire6194 = ( wire407  &  n_n1191 ) | ( wire226  &  wire249 ) ;
 assign wire6195 = ( wire120  &  n_n1039 ) | ( wire120  &  n_n1072 ) ;
 assign wire6200 = ( n_n1028  &  _9142 ) | ( n_n1028  &  _9143 ) ;
 assign wire6203 = ( wire334 ) | ( wire404  &  (~ n_n1121)  &  wire6176 ) ;
 assign wire6204 = ( wire333 ) | ( wire336 ) | ( wire6183  &  wire6184 ) ;
 assign wire6205 = ( wire337 ) | ( wire338 ) | ( wire339 ) | ( wire340 ) ;
 assign wire6206 = ( wire341 ) | ( wire342 ) | ( wire6200 ) ;
 assign wire6207 = ( wire6194 ) | ( wire6195 ) | ( _9164 ) ;
 assign wire6210 = ( wire6203 ) | ( wire6204 ) | ( wire6207 ) ;
 assign wire6213 = ( c  &  d ) | ( (~ c)  &  f ) | ( d  &  f ) | ( c  &  (~ f) ) | ( (~ c)  &  g ) | ( d  &  g ) | ( (~ f)  &  g ) ;
 assign wire6220 = ( (~ c)  &  (~ f)  &  i ) | ( (~ c)  &  g  &  i ) ;
 assign wire6222 = ( (~ j)  &  k  &  (~ m)  &  (~ n) ) ;
 assign wire6224 = ( (~ n_n857)  &  (~ n_n1260)  &  wire6222 ) ;
 assign wire6238 = ( (~ c)  &  (~ d)  &  (~ e)  &  f ) ;
 assign wire6239 = ( (~ a)  &  (~ e)  &  (~ f) ) ;
 assign wire6240 = ( i  &  (~ k)  &  (~ m)  &  (~ n) ) ;
 assign wire6241 = ( g  &  (~ l)  &  (~ m)  &  (~ n) ) ;
 assign wire6245 = ( wire170  &  wire6238 ) | ( n_n857  &  wire170  &  wire305 ) ;
 assign wire6246 = ( n_n1091  &  wire6240 ) | ( n_n1167  &  wire6241 ) ;
 assign wire6248 = ( n_n1189  &  _8970 ) | ( wire6224  &  _8976 ) ;
 assign wire6249 = ( wire316 ) | ( wire161  &  wire6239 ) ;
 assign wire6250 = ( wire317 ) | ( wire318 ) | ( wire85  &  _8993 ) ;
 assign wire6281 = ( wire253 ) | ( wire271 ) | ( wire272 ) | ( wire274 ) ;
 assign wire6282 = ( wire276 ) | ( wire278 ) | ( _9192 ) ;
 assign wire6283 = ( wire252 ) | ( wire269 ) | ( wire280 ) | ( wire281 ) ;
 assign wire6285 = ( wire6281 ) | ( wire6282 ) | ( wire6283 ) ;
 assign wire6286 = ( wire6205 ) | ( wire6206 ) | ( wire6210 ) | ( wire6285 ) ;
 assign wire6290 = ( (~ c)  &  h  &  (~ j) ) | ( (~ d)  &  h  &  (~ j) ) ;
 assign wire6292 = ( wire178 ) | ( n_n1036  &  wire6290 ) ;
 assign wire6298 = ( wire150 ) | ( wire163 ) | ( wire180 ) | ( wire6292 ) ;
 assign wire6300 = ( wire5954 ) | ( wire5955 ) | ( wire5969 ) | ( wire5970 ) ;
 assign wire6301 = ( wire140 ) | ( wire6298 ) | ( _8786 ) | ( _8801 ) ;
 assign wire6307 = ( g  &  (~ h)  &  (~ i) ) ;
 assign wire6309 = ( m  &  (~ n)  &  n_n997  &  wire6307 ) ;
 assign wire6317 = ( wire63 ) | ( n_n996  &  n_n1072  &  wire6309 ) ;
 assign wire6318 = ( wire42 ) | ( wire61 ) | ( wire66 ) ;
 assign _36 = ( f ) | ( b  &  e ) | ( b  &  (~ g) ) | ( (~ e)  &  (~ g) ) ;
 assign _37 = ( e  &  (~ n) ) | ( f  &  (~ n) ) | ( (~ g)  &  (~ n) ) ;
 assign _38 = ( e  &  m ) | ( f  &  m ) | ( (~ g)  &  m ) ;
 assign _70 = ( wire226  &  (~ wire395)  &  wire6045 ) ;
 assign _119 = ( n_n1261  &  n_n1260  &  (~ n_n1215)  &  _8882 ) ;
 assign _120 = ( n_n1261  &  (~ n_n1217)  &  n_n1260  &  _8882 ) ;
 assign _122 = ( (~ g)  &  n_n1261  &  wire85  &  _8878 ) ;
 assign _126 = ( n_n1217  &  n_n1215  &  wire6123 ) ;
 assign _182 = ( n_n711  &  n_n1210  &  n_n1094 ) | ( wire30  &  n_n1210  &  n_n1094 ) ;
 assign _183 = ( n_n841  &  n_n1210  &  _8711 ) ;
 assign _202 = ( n_n840  &  wire30  &  wire230  &  n_n1210 ) ;
 assign _203 = ( n_n840  &  n_n711  &  wire230  &  n_n1210 ) ;
 assign _217 = ( n_n920  &  n_n1201  &  wire5888  &  _7780 ) ;
 assign _218 = ( n_n918  &  n_n1195  &  wire5888  &  _7783 ) ;
 assign _224 = ( n_n920  &  n_n1201  &  n_n996  &  _7780 ) ;
 assign _225 = ( n_n918  &  n_n996  &  n_n1195  &  _7783 ) ;
 assign _226 = ( n_n840  &  wire221  &  wire5813 ) ;
 assign _227 = ( n_n709  &  wire221  &  _8574 ) ;
 assign _255 = ( n_n709  &  wire70  &  _8574 ) ;
 assign _256 = ( wire70  &  wire5813  &  _8577 ) ;
 assign _274 = ( wire41  &  wire5831 ) | ( wire5831  &  _8553 ) ;
 assign _275 = ( wire41  &  wire81 ) | ( wire81  &  _8553 ) ;
 assign _294 = ( wire113  &  n_n1228  &  wire15 ) ;
 assign _298 = ( n_n1207  &  n_n1228  &  wire15  &  _8533 ) ;
 assign _300 = ( wire22  &  n_n766  &  wire15 ) ;
 assign _313 = ( n_n904  &  wire190  &  n_n940 ) ;
 assign _314 = ( n_n904  &  wire22  &  _8063 ) ;
 assign _331 = ( wire31  &  n_n1187  &  n_n949  &  wire368 ) ;
 assign _333 = ( n_n1220  &  n_n876  &  n_n1082 ) ;
 assign _334 = ( n_n876  &  n_n1219  &  _8344 ) ;
 assign _335 = ( n_n1220  &  n_n949  &  n_n1082  &  _8469 ) ;
 assign _336 = ( n_n949  &  n_n1219  &  _8344  &  _8469 ) ;
 assign _373 = ( wire22  &  n_n857  &  n_n761 ) | ( wire113  &  n_n857  &  n_n761 ) ;
 assign _378 = ( wire69  &  wire5694  &  wire5695 ) | ( wire5694  &  wire5695  &  _8362 ) ;
 assign _379 = ( wire69  &  wire739  &  wire5695 ) | ( wire739  &  wire5695  &  _8362 ) ;
 assign _405 = ( n_n876  &  n_n1219  &  _8344 ) ;
 assign _446 = ( n_n1207  &  n_n893  &  n_n1177  &  _8202 ) ;
 assign _493 = ( b  &  (~ c)  &  d  &  (~ g) ) ;
 assign _494 = ( b  &  (~ c)  &  d  &  (~ f) ) ;
 assign _497 = ( n_n709  &  wire76  &  wire230 ) ;
 assign _507 = ( n_n876  &  wire190  &  n_n940 ) ;
 assign _508 = ( wire22  &  n_n876  &  _8063 ) ;
 assign _513 = ( n_n709  &  n_n1210  &  wire164 ) ;
 assign _559 = ( b  &  (~ d)  &  e  &  i ) ;
 assign _560 = ( b  &  (~ d)  &  e  &  (~ h) ) ;
 assign _561 = ( b  &  (~ d)  &  e  &  g ) ;
 assign _566 = ( wire58  &  wire29  &  n_n765 ) ;
 assign _576 = ( n_n618  &  wire34  &  n_n1204 ) | ( n_n618  &  n_n1204  &  wire35 ) ;
 assign _577 = ( n_n617  &  wire34  &  n_n1204 ) | ( n_n617  &  n_n1204  &  wire35 ) ;
 assign _589 = ( n_n978  &  wire211 ) ;
 assign _594 = ( n_n619  &  n_n623  &  n_n1216 ) ;
 assign _595 = ( wire34  &  n_n619  &  n_n1204 ) | ( n_n619  &  n_n1204  &  wire35 ) ;
 assign _611 = ( n_n840  &  n_n823  &  n_n982 ) ;
 assign _612 = ( n_n709  &  n_n982  &  _7745 ) ;
 assign _621 = ( wire76  &  n_n841  &  wire47 ) ;
 assign _624 = ( n_n711  &  wire76  &  n_n1094 ) | ( wire30  &  wire76  &  n_n1094 ) ;
 assign _665 = ( n_n920  &  n_n1201  &  wire265  &  _7780 ) ;
 assign _666 = ( n_n918  &  wire265  &  n_n1195  &  _7783 ) ;
 assign _670 = ( n_n904  &  wire228  &  _7776 ) | ( n_n904  &  wire265  &  _7776 ) ;
 assign _679 = ( n_n1036  &  n_n823  &  _7743 ) ;
 assign _680 = ( n_n709  &  n_n1036  &  _7745 ) ;
 assign _763 = ( n_n711  &  wire84  &  _7479 ) | ( n_n711  &  wire84  &  _7481 ) ;
 assign _803 = ( (~ e)  &  l  &  m  &  (~ n) ) ;
 assign _804 = ( (~ d)  &  l  &  m  &  (~ n) ) ;
 assign _814 = ( n_n893  &  n_n1177  &  n_n1253  &  _7528 ) ;
 assign _843 = ( n_n1207  &  wire84  &  wire202 ) ;
 assign _860 = ( g  &  wire233  &  n_n918  &  _7433 ) ;
 assign _861 = ( g  &  n_n1261  &  wire233  &  _7437 ) ;
 assign _877 = ( n_n1166  &  n_n1204  &  n_n628 ) ;
 assign _905 = ( n_n709  &  wire22  &  n_n857 ) | ( n_n709  &  wire113  &  n_n857 ) ;
 assign _7270 = ( (~ l)  &  m  &  (~ n) ) ;
 assign _7308 = ( b  &  (~ d)  &  e  &  (~ f) ) ;
 assign _7373 = ( c  &  (~ d)  &  f  &  wire65 ) ;
 assign _7387 = ( (~ f)  &  g  &  h ) ;
 assign _7390 = ( wire1155 ) | ( _877 ) | ( wire162  &  _7373 ) ;
 assign _7433 = ( (~ e)  &  m  &  (~ n) ) ;
 assign _7437 = ( (~ d)  &  e  &  m  &  (~ n) ) ;
 assign _7453 = ( wire1130 ) | ( wire1131 ) | ( _860 ) | ( _861 ) ;
 assign _7462 = ( e  &  (~ f) ) | ( (~ e)  &  g ) | ( (~ f)  &  g ) ;
 assign _7467 = ( (~ d)  &  e  &  (~ g) ) ;
 assign _7479 = ( (~ f)  &  (~ g)  &  (~ h) ) ;
 assign _7481 = ( (~ f)  &  g  &  (~ h) ) ;
 assign _7503 = ( (~ d)  &  e  &  m  &  (~ n) ) ;
 assign _7511 = ( d  &  e  &  m  &  (~ n) ) ;
 assign _7524 = ( d  &  e  &  m  &  (~ n) ) ;
 assign _7528 = ( (~ e)  &  f  &  (~ h) ) ;
 assign _7541 = ( (~ e)  &  g  &  (~ h) ) ;
 assign _7556 = ( d  &  e  &  m  &  (~ n) ) ;
 assign _7569 = ( d  &  e  &  m  &  (~ n) ) ;
 assign _7632 = ( a  &  (~ c)  &  d ) ;
 assign _7649 = ( wire5226 ) | ( wire94  &  _7632 ) ;
 assign _7662 = ( (~ e)  &  g  &  (~ i)  &  (~ n) ) ;
 assign _7671 = ( (~ e)  &  g  &  i ) ;
 assign _7743 = ( b  &  d  &  (~ e) ) ;
 assign _7745 = ( (~ f)  &  h  &  j ) ;
 assign _7751 = ( b  &  (~ d)  &  e  &  j ) ;
 assign _7757 = ( (~ c)  &  d  &  (~ e)  &  j ) ;
 assign _7759 = ( b  &  d  &  (~ e)  &  j ) ;
 assign _7776 = ( (~ e)  &  g  &  (~ i) ) ;
 assign _7780 = ( (~ n)  &  m ) ;
 assign _7783 = ( (~ n)  &  m ) ;
 assign _7794 = ( f  &  g  &  (~ h) ) ;
 assign _7798 = ( k  &  m  &  (~ n) ) ;
 assign _7815 = ( k  &  m  &  (~ n) ) ;
 assign _7833 = ( (~ f)  &  g  &  j ) ;
 assign _7862 = ( l  &  (~ m)  &  n ) ;
 assign _7877 = ( _611 ) | ( _612 ) | ( n_n978  &  wire208 ) ;
 assign _7920 = ( n_n617  &  n_n623  &  _7862 ) | ( n_n618  &  n_n623  &  _7862 ) ;
 assign _7925 = ( a  &  c  &  (~ d) ) ;
 assign _7927 = ( (~ e)  &  g  &  i ) ;
 assign _8063 = ( e  &  f  &  h ) ;
 assign _8076 = ( wire850 ) | ( _497 ) | ( _507 ) | ( _508 ) ;
 assign _8084 = ( (~ b)  &  d  &  f ) ;
 assign _8097 = ( c  &  e  &  wire120 ) ;
 assign _8115 = ( wire849 ) | ( wire5513 ) | ( wire92  &  _8097 ) ;
 assign _8116 = ( n_n1425 ) | ( wire843 ) | ( wire845 ) | ( wire858 ) ;
 assign _8202 = ( b  &  d  &  (~ e) ) ;
 assign _8227 = ( wire789 ) | ( wire791 ) ;
 assign _8242 = ( wire5618 ) | ( wire802 ) ;
 assign _8243 = ( wire5619 ) | ( wire5611 ) | ( wire5615 ) | ( _8227 ) ;
 assign _8290 = ( (~ c)  &  (~ d)  &  (~ f)  &  (~ g) ) ;
 assign _8318 = ( n_n2602 ) | ( wire775 ) | ( wire776 ) | ( n_n2511 ) ;
 assign _8344 = ( e  &  h  &  k ) ;
 assign _8362 = ( wire31  &  wire368 ) ;
 assign _8370 = ( a  &  c  &  e  &  (~ f) ) ;
 assign _8385 = ( k  &  m  &  (~ n) ) ;
 assign _8388 = ( (~ n_n1082)  &  wire5699 ) | ( wire5699  &  (~ _8385) ) ;
 assign _8391 = ( a  &  c  &  (~ d) ) ;
 assign _8394 = ( wire716 ) | ( wire44  &  (~ wire743)  &  _8388 ) ;
 assign _8427 = ( (~ e)  &  g  &  h ) ;
 assign _8439 = ( f  &  (~ g)  &  (~ h)  &  i ) ;
 assign _8469 = ( (~ n)  &  m ) ;
 assign _8474 = ( _333 ) | ( _334 ) | ( _335 ) | ( _336 ) ;
 assign _8487 = ( d  &  (~ e)  &  m  &  (~ n) ) ;
 assign _8504 = ( wire646 ) | ( wire650 ) | ( wire653 ) ;
 assign _8515 = ( _313 ) | ( _314 ) | ( wire200  &  n_n872 ) ;
 assign _8524 = ( wire664 ) | ( wire5795 ) | ( _8504 ) | ( _8515 ) ;
 assign _8533 = ( k  &  m  &  (~ n) ) ;
 assign _8543 = ( n_n2953 ) | ( wire619 ) | ( _294 ) | ( _300 ) ;
 assign _8553 = ( n_n1161  &  n_n904 ) | ( wire16  &  _7794 ) ;
 assign _8574 = ( (~ f)  &  h  &  i ) ;
 assign _8577 = ( b  &  d  &  (~ e) ) ;
 assign _8608 = ( (~ e)  &  g  &  i ) ;
 assign _8619 = ( h  &  i  &  j ) ;
 assign _8636 = ( (~ n)  &  m ) ;
 assign _8639 = ( n_n698  &  wire81  &  _8636 ) | ( n_n698  &  wire583  &  _8636 ) ;
 assign _8646 = ( _224 ) | ( _225 ) | ( _226 ) | ( _227 ) ;
 assign _8668 = ( wire5898 ) | ( wire5899 ) | ( _8639 ) | ( _8646 ) ;
 assign _8701 = ( wire5814 ) | ( wire547 ) | ( _255 ) | ( _256 ) ;
 assign _8711 = ( b  &  e  &  (~ f) ) ;
 assign _8715 = ( wire5938 ) | ( wire5905 ) | ( wire5906 ) | ( _8668 ) ;
 assign _8731 = ( (~ e)  &  f  &  m  &  (~ n) ) ;
 assign _8732 = ( a  &  b  &  c  &  (~ d) ) ;
 assign _8742 = ( (~ j)  &  (~ m)  &  n ) ;
 assign _8746 = ( (~ e)  &  (~ l)  &  m  &  (~ n) ) ;
 assign _8747 = ( a  &  b  &  c  &  (~ d) ) ;
 assign _8748 = ( (~ k)  &  m  &  (~ n) ) ;
 assign _8750 = ( i  &  (~ m)  &  (~ n) ) ;
 assign _8769 = ( n_n1089  &  wire127 ) | ( wire127  &  n_n1160 ) ;
 assign _8771 = ( i  &  m  &  (~ n) ) ;
 assign _8772 = ( (~ g)  &  c ) ;
 assign _8776 = ( n_n1039  &  _8771 ) | ( wire226  &  _8772 ) ;
 assign _8786 = ( wire173 ) | ( wire177 ) | ( n_n1036  &  n_n1022 ) ;
 assign _8794 = ( (~ j)  &  (~ k)  &  (~ l) ) ;
 assign _8801 = ( wire6145 ) | ( wire6147 ) | ( _8769 ) | ( _8776 ) ;
 assign _8819 = ( (~ d)  &  (~ e)  &  (~ f)  &  j ) ;
 assign _8820 = ( (~ d)  &  (~ e)  &  (~ f)  &  i ) ;
 assign _8823 = ( (~ l)  &  (~ m)  &  (~ n) ) ;
 assign _8830 = ( i  &  (~ m)  &  n ) | ( j  &  (~ m)  &  n ) ;
 assign _8835 = ( (~ l)  &  (~ m)  &  n ) ;
 assign _8851 = ( (~ h)  &  i  &  (~ m)  &  n ) ;
 assign _8855 = ( (~ e)  &  (~ f)  &  (~ m)  &  n ) ;
 assign _8868 = ( (~ g)  &  m  &  (~ n) ) | ( (~ h)  &  m  &  (~ n) ) ;
 assign _8878 = ( (~ d)  &  (~ e)  &  m  &  (~ n) ) ;
 assign _8880 = ( h  &  (~ i)  &  (~ m)  &  n ) ;
 assign _8882 = ( (~ n)  &  m ) ;
 assign _8890 = ( wire440 ) | ( wire441 ) | ( _122 ) | ( _126 ) ;
 assign _8939 = ( (~ i)  &  (~ m)  &  (~ n) ) ;
 assign _8940 = ( c  &  (~ d)  &  (~ e)  &  (~ f) ) ;
 assign _8970 = ( (~ l)  &  m  &  (~ n) ) ;
 assign _8976 = ( (~ d)  &  wire6220 ) | ( e  &  wire6220 ) | ( (~ g)  &  wire6220 ) ;
 assign _8993 = ( (~ d)  &  (~ e)  &  (~ f)  &  (~ g) ) ;
 assign _8998 = ( (~ g)  &  (~ h)  &  (~ n) ) ;
 assign _9007 = ( (~ g)  &  l  &  (~ m)  &  (~ n) ) ;
 assign _9018 = ( (~ e)  &  (~ h)  &  i ) ;
 assign _9020 = ( (~ c)  &  d  &  (~ g) ) ;
 assign _9021 = ( wire70  &  _9018 ) | ( wire226  &  _9020 ) ;
 assign _9051 = ( wire504 ) | ( wire505 ) | ( wire5990 ) ;
 assign _9054 = ( (~ a)  &  (~ e)  &  (~ f)  &  (~ g) ) ;
 assign _9055 = ( (~ g)  &  m  &  (~ n) ) ;
 assign _9062 = ( (~ b)  &  f  &  (~ h) ) ;
 assign _9064 = ( (~ h)  &  (~ i)  &  (~ j) ) ;
 assign _9065 = ( wire301  &  _9062 ) | ( wire58  &  _9064 ) ;
 assign _9067 = ( (~ j)  &  (~ m)  &  n ) | ( k  &  (~ m)  &  n ) ;
 assign _9075 = ( wire85  &  _9054 ) | ( n_n1189  &  wire85  &  _9055 ) ;
 assign _9076 = ( wire500 ) | ( wire501 ) | ( _9065 ) | ( _9075 ) ;
 assign _9092 = ( h  &  i  &  (~ m)  &  n ) ;
 assign _9094 = ( h  &  i  &  (~ m)  &  n ) ;
 assign _9128 = ( wire5998 ) | ( wire6036 ) | ( wire6037 ) | ( _9051 ) ;
 assign _9142 = ( b  &  (~ m)  &  n ) | ( j  &  (~ m)  &  n ) ;
 assign _9143 = ( k  &  (~ m)  &  n ) ;
 assign _9161 = ( i  &  (~ m)  &  n ) ;
 assign _9163 = ( (~ d)  &  (~ m)  &  n ) ;
 assign _9164 = ( n_n1028  &  _9161 ) | ( n_n1121  &  _9163 ) ;
 assign _9184 = ( e  &  (~ g)  &  h  &  (~ j) ) ;
 assign _9185 = ( (~ c)  &  (~ d)  &  (~ e)  &  h ) ;
 assign _9186 = ( (~ c)  &  (~ d)  &  (~ e)  &  g ) ;
 assign _9190 = ( (~ c)  &  e  &  (~ f) ) ;
 assign _9192 = ( n_n1036  &  _9184 ) | ( wire6272  &  _9190 ) ;
 assign _9203 = ( (~ g)  &  (~ h)  &  (~ m)  &  (~ n) ) ;
 assign _9209 = ( wire6251 ) | ( wire6252 ) | ( wire6256 ) | ( wire6070 ) ;


endmodule

