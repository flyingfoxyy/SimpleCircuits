module apex2_mapped (
	i_30_, i_20_, i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, 
	i_27_, i_14_, i_3_, i_28_, i_13_, i_4_, i_25_, i_12_, i_1_, i_26_, 
	i_11_, i_2_, i_23_, i_18_, i_24_, i_17_, i_0_, i_21_, i_16_, i_22_, 
	i_15_, i_32_, i_31_, i_34_, i_33_, i_19_, i_36_, i_35_, i_38_, i_29_, 
	i_37_, o_1_, o_2_, o_0_);

input i_30_, i_20_, i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_27_, i_14_, i_3_, i_28_, i_13_, i_4_, i_25_, i_12_, i_1_, i_26_, i_11_, i_2_, i_23_, i_18_, i_24_, i_17_, i_0_, i_21_, i_16_, i_22_, i_15_, i_32_, i_31_, i_34_, i_33_, i_19_, i_36_, i_35_, i_38_, i_29_, i_37_;

output o_1_, o_2_, o_0_;

wire wire7250, wire7257, wire7714, wire7747, n_n1542, wire8096, wire59, n_n1862, wire7370, wire7371, wire7383, n_n1827, n_n1870, wire627, n_n1829, wire7432, wire7433, wire7441, wire990, wire991, wire992, wire993, n_n1866, wire983, wire987, wire7727, wire7728, n_n1865, wire7771, n_n1548, n_n1545, wire7923, wire8079, wire232, n_n1443, wire79, n_n460, wire462, wire227, wire493, wire58, n_n1441, wire43, wire302, n_n1433, n_n1425, wire54, n_n1396, wire10, n_n1404, n_n1390, wire415, n_n1372, n_n1369, n_n1429, n_n1454, n_n1489, n_n1353, n_n1361, n_n1423, n_n1295, n_n1439, wire3, n_n1438, n_n1397, n_n1274, n_n1334, n_n1368, n_n1216, wire290, n_n1391, n_n1478, n_n1307, n_n1374, n_n805, n_n1504, n_n841, n_n853, n_n793, n_n1315, n_n1092, n_n1406, n_n1466, wire224, n_n1278, n_n787, n_n1197, n_n762, n_n1038, n_n1314, n_n1375, wire13, n_n1141, wire7086, n_n544, n_n1486, n_n1408, n_n1318, n_n504, wire404, wire297, n_n416, n_n1305, n_n1118, n_n1279, n_n358, n_n1048, n_n1144, n_n307, n_n1263, n_n1306, n_n620, n_n1288, n_n1018, n_n1400, n_n819, wire7419, wire7425, n_n394, n_n458, wire7426, n_n391, n_n1055, n_n461, wire7411, n_n372, n_n1179, wire7265, wire257, n_n300, n_n1225, wire7412, n_n294, n_n301, n_n880, n_n1100, wire51, wire260, n_n437, n_n571, n_n1258, wire263, n_n825, n_n1437, n_n1340, n_n180, n_n132, n_n152, n_n1300, n_n1472, wire50, wire52, wire85, n_n1303, wire223, wire264, wire61, wire388, wire446, wire262, wire18, wire436, wire529, wire7511, wire7512, n_n1147, n_n1089, wire298, wire244, wire7789, wire410, wire7785, wire516, n_n1322, wire7243, wire530, wire935, wire7793, wire7794, wire7795, n_n1580, n_n1326, wire245, wire277, wire340, n_n1213, wire533, n_n1323, wire532, wire7806, wire7807, wire7808, n_n1579, wire80, wire536, n_n1285, wire535, wire918, wire7812, wire7813, n_n1581, n_n1519, n_n1419, n_n1302, n_n1401, wire283, n_n1192, n_n1257, n_n1133, n_n1128, n_n586, n_n1523, n_n269, wire259, n_n242, n_n1202, wire258, n_n355, n_n1345, wire7413, n_n371, n_n316, n_n735, wire7423, n_n315, n_n984, n_n1458, n_n177, n_n1241, n_n179, n_n245, n_n1431, wire7491, wire7266, wire70, wire7492, wire212, wire239, wire288, wire539, wire7409, wire537, wire7494, wire7495, n_n1881, n_n576, n_n1499, wire47, wire44, wire7749, wire7847, wire307, wire541, n_n329, wire468, wire67, wire367, wire540, n_n195, wire864, wire7874, wire7875, wire86, wire275, wire483, wire500, wire41, wire221, wire495, wire7189, wire543, wire7866, wire7916, wire7917, wire7920, n_n1497, n_n1384, n_n1393, n_n1282, n_n839, n_n1311, n_n263, n_n363, n_n584, n_n1033, wire7420, n_n309, wire7424, n_n317, n_n712, n_n284, n_n1028, n_n178, wire57, wire77, wire83, wire372, wire380, wire71, wire395, wire503, n_n1387, n_n1359, n_n1080, n_n1254, wire196, wire7926, wire7927, n_n1585, n_n1422, wire8, wire38, wire1661, wire7682, wire112, wire7029, wire127, wire546, wire7938, n_n1556, n_n1459, n_n1377, n_n1312, n_n820, n_n706, wire205, n_n1191, wire7051, n_n608, n_n1058, n_n916, n_n629, wire12, n_n338, wire261, n_n129, n_n26, wire463, wire966, wire967, wire338, wire7753, wire547, wire451, wire7952, wire7953, wire7954, n_n1574, wire412, wire7963, wire7964, wire7965, n_n1575, wire7979, wire7981, n_n1578, wire195, wire7989, wire7990, wire7991, n_n1576, wire8003, n_n1577, wire174, wire176, wire8035, wire8036, wire8037, n_n1573, wire8046, wire8047, n_n1572, wire8052, wire8054, n_n1251, n_n998, wire124, wire132, wire550, wire8061, wire8062, n_n1583, n_n1582, wire557, wire555, wire8072, n_n1584, wire214, wire265, wire267, wire559, wire6920, wire312, wire6948, wire6949, wire126, wire7653, wire128, wire1649, wire1650, wire452, wire7761, wire363, wire420, wire7769, wire455, wire956, wire958, wire7776, wire7777, wire568, n_n1511, n_n130, wire475, wire7050, n_n849, n_n1059, wire222, n_n18, n_n21, wire7942, wire299, wire6993, wire342, wire7831, wire478, wire572, wire48, wire385, wire7822, wire418, wire578, wire384, wire576, wire253, wire330, wire405, wire583, wire1281, wire1283, n_n1847, wire585, wire7615, n_n1889, wire361, wire353, wire4, wire7276, wire56, wire226, wire7272, wire1449, wire1450, wire7282, n_n1856, wire81, wire377, wire1457, wire7267, wire7290, n_n1825, wire1428, wire1429, wire1430, wire1431, n_n1854, wire1382, wire1383, wire1384, wire7345, n_n1861, wire319, wire6951, wire6952, wire599, wire6958, wire598, wire6957, wire597, wire6961, wire6962, wire6963, n_n1718, wire317, wire365, wire601, wire273, wire256, wire600, wire6876, wire233, wire246, wire492, wire63, wire268, wire431, wire6899, wire508, wire7053, wire7976, wire301, wire7827, wire7828, wire608, wire360, wire437, wire891, wire610, n_n1149, wire447, wire434, wire7415, wire7466, wire235, wire1264, wire1265, wire1266, wire1267, n_n1846, wire1111, wire616, wire615, wire614, wire1105, wire1106, n_n1892, wire35, wire7631, wire7632, n_n1837, wire7301, wire249, wire311, wire78, wire329, wire344, wire1372, wire1377, wire7357, wire7358, wire218, wire7377, wire310, wire315, wire387, wire408, wire784, wire1337, wire7400, wire271, wire278, wire346, wire1330, wire320, wire416, wire630, wire629, wire1715, wire1717, wire6977, n_n1719, wire248, wire634, wire6937, wire6938, wire632, wire88, wire1565, wire1566, wire1567, wire1697, wire1701, wire6989, wire6990, n_n1720, wire1690, wire7001, n_n1716, wire1683, wire7010, wire7011, n_n1715, wire1659, n_n1723, wire7033, wire7044, wire7045, wire440, wire644, wire643, wire1086, wire1087, wire254, wire381, wire430, wire429, wire1289, n_n1852, wire755, wire1314, wire1316, n_n1843, wire75, wire654, wire276, wire7427, wire423, wire314, wire7136, wire664, wire663, wire29, wire491, wire7062, n_n1690, wire668, wire383, wire669, wire390, wire435, wire1323, wire1324, wire1256, wire1257, wire1258, wire1259, n_n1844, wire270, wire677, wire7477, n_n1821, wire272, wire379, wire482, wire74, wire189, wire687, wire68, wire692, wire7502, wire7503, wire7504, wire524, wire694, wire6960, wire7017, wire693, wire1587, wire7110, n_n1714, wire470, wire698, wire1542, wire7169, wire697, n_n1703, wire8010, wire295, wire7523, wire286, wire1214, wire7006, wire306, wire6984, wire7173, wire7174, wire705, wire7177, wire704, wire1525, wire7183, n_n1704, wire708, wire1511, wire7188, wire712, wire289, wire327, wire335, wire7356, wire456, wire305, wire717, wire716, wire6928, wire1498, wire1499, wire1500, wire1501, n_n1701, wire1490, wire1493, wire7221, wire274, wire7121, wire351, wire724, wire7898, wire8021, wire8022, wire723, wire394, wire6996, wire6997, wire322, wire727, wire1581, wire7116, wire7117, n_n1713, wire731, wire151, wire345, wire735, wire7686, wire734, wire7547, wire502, wire1190, wire1191, wire7548, wire7549, n_n1875, wire1202, wire1203, wire7537, wire7538, n_n1873, wire7570, n_n1831, wire7598, wire740, wire7639, wire739, wire7622, wire7642, n_n1818, wire1043, wire7680, n_n1834, n_n1887, wire7705, n_n1835, wire744, wire745, wire1053, wire1054, wire7661, wire457, wire465, wire510, wire1474, wire7244, n_n1712, wire515, wire1634, wire771, wire7588, wire7591, wire425, wire454, wire1338, wire7399, wire1069, wire792, wire7699, wire7145, wire484, wire7148, wire489, wire7428, wire422, wire349, wire413, wire7342, wire7343, wire37, wire211, wire65, wire1663, wire802, wire95, wire96, wire143, wire7178, wire458, wire7274, wire231, wire7055, wire251, wire334, wire343, wire7890, wire356, wire402, wire1432, wire1433, wire1434, wire406, wire1342, wire1343, wire7576, wire438, wire1340, wire1341, wire498, wire517, wire521, wire522, wire7254, wire526, wire544, wire7259, wire582, wire590, wire593, wire604, wire6892, wire6894, wire603, wire6913, wire606, wire624, wire635, wire1570, wire1572, wire1573, wire638, wire657, wire661, wire666, wire7473, wire679, wire1604, wire683, wire710, wire713, wire7217, wire721, wire741, wire759, wire758, wire767, wire1766, wire22, wire1767, wire1768, wire34, wire105, wire107, wire8090, wire8091, wire8086, wire6947, wire110, wire111, wire117, wire8056, wire8057, wire130, wire133, wire134, wire142, wire150, wire7058, wire8042, wire8043, wire158, wire160, wire161, wire163, wire169, wire164, wire8008, wire166, wire172, wire8007, wire178, wire7802, wire183, wire184, wire7803, wire185, wire187, wire7997, wire7999, wire7984, wire192, wire194, wire200, wire201, wire197, wire198, wire7105, wire7971, wire234, wire304, wire7787, wire336, wire339, wire7784, wire350, wire7961, wire417, wire7949, wire424, wire7940, wire427, wire439, wire7945, wire469, wire471, wire7930, wire494, wire6982, wire7931, wire497, wire507, wire7025, wire512, wire813, wire7900, wire825, wire829, wire7901, wire833, wire7903, wire834, wire7887, wire7892, wire843, wire849, wire857, wire850, wire7868, wire7871, wire7819, wire881, wire7858, wire7859, wire7862, wire875, wire7860, wire7820, wire910, wire911, wire906, wire7791, wire919, wire7798, wire924, wire925, wire926, wire928, wire7782, wire933, wire937, wire939, wire942, wire943, wire948, wire945, wire7778, wire950, wire953, wire7765, wire7766, wire7751, wire7757, wire969, wire981, wire7736, wire977, wire978, wire988, wire7258, wire7723, wire1406, wire7716, wire994, wire996, wire7718, wire7717, wire7701, wire999, wire7702, wire1000, wire7704, wire1008, wire1009, wire7308, wire7690, wire1010, wire7691, wire1011, wire1015, wire1012, wire1014, wire1017, wire1022, wire1023, wire1024, wire7670, wire1029, wire1030, wire1032, wire1033, wire1041, wire1044, wire1045, wire7655, wire1050, wire7657, wire1051, wire1052, wire7644, wire1060, wire7647, wire1062, wire1064, wire1077, wire7638, wire1070, wire1082, wire7636, wire1080, wire1081, wire1089, wire1091, wire1095, wire1100, wire1101, wire7616, wire1112, wire7618, wire1113, wire1121, wire7619, wire1114, wire1123, wire7612, wire7600, wire1131, wire7602, wire1132, wire7603, wire1133, wire1134, wire1137, wire1135, wire1136, wire1147, wire1139, wire1140, wire1150, wire1141, wire1142, wire1143, wire7582, wire1152, wire1156, wire1157, wire7572, wire1159, wire1161, wire1164, wire1162, wire1168, wire7559, wire1173, wire1176, wire1197, wire7541, wire7543, wire1198, wire7532, wire1201, wire7534, wire1211, wire1227, wire7488, wire1230, wire1234, wire1235, wire7479, wire1238, wire1240, wire1242, wire1253, wire7474, wire1247, wire1249, wire1260, wire7469, wire7470, wire7431, wire1263, wire7465, wire7271, wire7459, wire1268, wire1271, wire7456, wire1274, wire7454, wire7446, wire1286, wire1291, wire1303, wire1305, wire7430, wire1308, wire1309, wire1317, wire1319, wire7402, wire1325, wire1347, wire7388, wire1349, wire7390, wire1350, wire1351, wire7375, wire1356, wire1357, wire7364, wire1367, wire1379, wire7352, wire7344, wire7332, wire1392, wire7317, wire1399, wire1404, wire1405, wire1403, wire7324, wire1426, wire1412, wire1408, wire1414, wire1435, wire1436, wire1416, wire1417, wire7297, wire1419, wire7311, wire7296, wire7298, wire7299, wire1443, wire7284, wire7285, wire1437, wire7288, wire1439, wire7275, wire7281, wire1460, wire7261, wire1456, wire1461, wire1463, wire1464, wire7264, wire6906, wire1480, wire6998, wire1476, wire7108, wire7224, wire7214, wire7228, wire1483, wire7229, wire1484, wire1576, wire1577, wire7230, wire1507, wire1508, wire7212, wire7215, wire7216, wire7218, wire7219, wire7195, wire7199, wire1502, wire7205, wire7197, wire1514, wire7185, wire7187, wire1509, wire7191, wire6885, wire7186, wire1539, wire7158, wire7160, wire1534, wire7161, wire7163, wire7159, wire7151, wire1546, wire1548, wire1550, wire1551, wire1552, wire1549, wire1553, wire1554, wire7153, wire1561, wire1559, wire6882, wire7120, wire1574, wire7126, wire7130, wire7123, wire7059, wire1580, wire1583, wire1582, wire1585, wire1586, wire1592, wire1593, wire7009, wire1589, wire1591, wire1600, wire7099, wire1597, wire1603, wire7080, wire1607, wire7084, wire1608, wire1611, wire7083, wire7063, wire7064, wire1618, wire1623, wire1625, wire7072, wire1622, wire7068, wire7069, wire7070, wire7046, wire1628, wire1632, wire7054, wire1635, wire1637, wire1640, wire1651, wire1652, wire1653, wire7031, wire1654, wire1656, wire1657, wire7028, wire7026, wire7027, wire1668, wire1675, wire1676, wire1670, wire6959, wire1672, wire1677, wire1678, wire1684, wire1691, wire1696, wire6979, wire1698, wire1699, wire1700, wire1702, wire1703, wire1704, wire6955, wire1706, wire1709, wire1710, wire6971, wire6973, wire1718, wire1719, wire6967, wire1730, wire1731, wire1726, wire6939, wire1738, wire6908, wire1748, wire1749, wire1750, wire1747, wire1753, wire6910, wire6912, wire6884, wire1756, wire1757, wire1758, wire6889, wire6879, wire6880, wire6891, wire6898, wire6901, wire6903, wire6905, wire6917, wire6919, wire6922, wire6923, wire6924, wire6926, wire6927, wire6930, wire6931, wire6933, wire6934, wire6936, wire6941, wire6942, wire6943, wire6953, wire6994, wire7004, wire7014, wire7022, wire7036, wire7037, wire7040, wire7041, wire7043, wire7075, wire7076, wire7079, wire7085, wire7087, wire7089, wire7090, wire7093, wire7095, wire7096, wire7097, wire7102, wire7103, wire7104, wire7114, wire7119, wire7134, wire7135, wire7137, wire7139, wire7140, wire7141, wire7142, wire7143, wire7152, wire7157, wire7165, wire7166, wire7175, wire7179, wire7190, wire7203, wire7204, wire7208, wire7210, wire7211, wire7234, wire7238, wire7239, wire7240, wire7247, wire7248, wire7256, wire7268, wire7269, wire7277, wire7286, wire7295, wire7306, wire7309, wire7312, wire7319, wire7320, wire7321, wire7322, wire7323, wire7325, wire7327, wire7328, wire7329, wire7330, wire7331, wire7333, wire7334, wire7335, wire7336, wire7337, wire7339, wire7340, wire7341, wire7348, wire7350, wire7351, wire7354, wire7355, wire7361, wire7362, wire7363, wire7365, wire7366, wire7367, wire7368, wire7372, wire7373, wire7374, wire7379, wire7380, wire7385, wire7386, wire7387, wire7394, wire7395, wire7457, wire7458, wire7483, wire7485, wire7510, wire7516, wire7521, wire7525, wire7526, wire7529, wire7531, wire7536, wire7545, wire7552, wire7553, wire7555, wire7567, wire7574, wire7577, wire7580, wire7585, wire7586, wire7592, wire7595, wire7609, wire7621, wire7626, wire7627, wire7651, wire7676, wire7678, wire7689, wire7703, wire7711, wire7721, wire7725, wire7726, wire7731, wire7732, wire7733, wire7734, wire7737, wire7738, wire7740, wire7741, wire7743, wire7744, wire7750, wire7763, wire7772, wire7781, wire7810, wire7811, wire7817, wire7823, wire7825, wire7829, wire7830, wire7832, wire7834, wire7835, wire7836, wire7837, wire7838, wire7840, wire7842, wire7843, wire7844, wire7845, wire7849, wire7852, wire7853, wire7854, wire7855, wire7856, wire7857, wire7863, wire7864, wire7867, wire7869, wire7870, wire7879, wire7881, wire7885, wire7888, wire7889, wire7893, wire7895, wire7896, wire7897, wire7899, wire7902, wire7906, wire7907, wire7909, wire7910, wire7911, wire7912, wire7913, wire7914, wire7915, wire7918, wire7921, wire7932, wire7935, wire7936, wire7941, wire7947, wire7957, wire7958, wire7959, wire7960, wire7969, wire7986, wire7994, wire8014, wire8019, wire8023, wire8026, wire8027, wire8028, wire8029, wire8030, wire8031, wire8039, wire8041, wire8077, wire8082, wire8084, wire8093, wire8094, _3, _4, _31, _32, _41, _42, _43, _62, _63, _64, _67, _75, _77, _78, _79, _80, _81, _82, _90, _96, _97, _107, _180, _188, _189, _221, _231, _232, _240, _278, _279, _282, _283, _292, _293, _294, _303, _322, _335, _336, _338, _342, _343, _363, _364, _365, _390, _400, _401, _402, _406, _407, _410, _411, _415, _418, _419, _439, _442, _451, _460, _490, _495, _510, _526, _530, _531, _539, _543, _585, _588, _589, _595, _606, _609, _612, _613, _614, _615, _617, _624, _626, _627, _635, _637, _655, _656, _657, _658, _662, _664, _665, _668, _674, _676, _677, _678, _679, _683, _684, _685, _686, _702, _733, _744, _746, _747, _749, _750, _756, _757, _758, _761, _763, _767, _781, _782, _788, _789, _791, _795, _796, _797, _799, _800, _803, _816, _817, _818, _820, _821, _822, _823, _832, _833, _834, _835, _844, _860, _881, _899, _927, _928, _929, _963, _975, _983, _993, _995, _996, _1002, _1003, _1005, _1006, _1015, _1016, _1020, _1021, _1027, _1070, _1074, _1076, _1082, _1083, _1084, _1089, _1090, _1098, _1099, _1102, _1103, _1104, _1105, _1106, _1108, _1109, _1110, _1111, _1114, _1115, _1134, _1135, _9202, _9206, _9225, _9227, _9290, _9309, _9314, _9318, _9322, _9325, _9328, _9338, _9344, _9347, _9351, _9354, _9361, _9379, _9399, _9404, _9408, _9409, _9456, _9459, _9463, _9466, _9470, _9480, _9483, _9494, _9495, _9498, _9499, _9511, _9514, _9542, _9551, _9553, _9577, _9583, _9584, _9587, _9598, _9607, _9611, _9613, _9616, _9619, _9621, _9636, _9644, _9652, _9659, _9673, _9674, _9678, _9683, _9684, _9686, _9688, _9724, _9733, _9736, _9737, _9740, _9748, _9751, _9753, _9754, _9755, _9758, _9760, _9781, _9784, _9804, _9821, _9834, _9836, _9847, _9851, _9857, _9868, _9872, _9876, _9880, _9882, _9889, _9890, _9892, _9895, _9896, _9898, _9899, _9901, _9907, _9908, _9913, _9918, _9919, _9922, _9929, _9934, _9950, _9959, _9963, _9992, _9996, _9998, _9999, _10003, _10004, _10022, _10025, _10034, _10038, _10041, _10045, _10051, _10053, _10062, _10073, _10075, _10085, _10108, _10112, _10125, _10130, _10132, _10133, _10137, _10142, _10143, _10151, _10160, _10169, _10171, _10173, _10175, _10176, _10177, _10181, _10184, _10186, _10188, _10190, _10192, _10197, _10205, _10216, _10232, _10281, _10282, _10283, _10286, _10288, _10290, _10292, _10294, _10313, _10317, _10319, _10324, _10326, _10331, _10332, _10341, _10353, _10370, _10372, _10377, _10386, _10408, _10409, _10425, _10426, _10430, _10432, _10445, _10448, _10457, _10458, _10460, _10465, _10469, _10475, _10477, _10478, _10480, _10484, _10485, _10491, _10496, _10498, _10504, _10524, _10526, _10531, _10533, _10534, _10536, _10560, _10575, _10578, _10586, _10606, _10607, _10625, _10626, _10628, _10631, _10632, _10634, _10635, _10646, _10648, _10651, _10658, _10663, _10665, _10667, _10679, _10690, _10693, _10705, _10708, _10715, _10716, _10717, _10721, _10722, _10731, _10746, _10748, _10754, _10759, _10762, _10782, _10785, _10790, _10811, _10814, _10816, _10819, _10822, _10823, _10826, _10827, _10828, _10829, _10830, _10831, _10833, _10846, _10849, _10850, _10870, _10876, _10877, _10879, _10885, _10889, _10917, _10918, _10933, _10937, _10942, _10948, _10950, _10962, _10970, _10972, _10974, _10984, _10985, _10990, _10991, _10994, _10995, _10998, _10999, _11001, _11016, _11020, _11021, _11023, _11024, _11027, _11029, _11033, _11037, _11051, _11052, _11053, _11055, _11056, _11063, _11077, _11087, _11089, _11093, _11094, _11097, _11113, _11117, _11118, _11119, _11120, _11141, _11146, _11170, _11202, _11205, _11215, _11227, _11262, _11294, _11296, _11307, _11309, _11313, _11315, _11325, _11326, _11333, _11334, _11336, _11343, _11350, _11354, _11360, _11361, _11362, _11363, _11365, _11366, _11372, _11388, _11391, _11393, _11395, _11400, _11419, _11422, _11424, _11425, _11428, _11430, _11431, _11443, _11479, _11482, _11489, _11495, _11510, _11519, _11521, _11531, _11532, _11544;

assign o_1_ = ( wire7239 ) | ( wire7240 ) | ( _9901 ) | ( _9963 ) ;
 assign o_2_ = ( wire7747 ) | ( wire7744 ) | ( _10759 ) | ( _10974 ) ;
 assign o_0_ = ( n_n1542 ) | ( wire8096 ) | ( _11544 ) ;
 assign wire7250 = ( wire1597 ) | ( wire7104 ) | ( wire7247 ) | ( wire7248 ) ;
 assign wire7257 = ( wire7256 ) | ( _844 ) | ( wire526  &  _9907 ) ;
 assign wire7714 = ( n_n1818 ) | ( n_n1834 ) | ( n_n1835 ) | ( wire7711 ) ;
 assign wire7747 = ( wire7441 ) | ( wire7350 ) | ( _10833 ) | ( _10972 ) ;
 assign n_n1542 = ( n_n1548 ) | ( n_n1545 ) | ( wire7923 ) | ( wire8079 ) ;
 assign wire8096 = ( wire945 ) | ( wire7781 ) | ( wire8093 ) | ( wire8094 ) ;
 assign wire59 = ( (~ i_33_)  &  i_37_ ) ;
 assign n_n1862 = ( wire1372 ) | ( wire1377 ) | ( wire7357 ) | ( wire7358 ) ;
 assign wire7370 = ( wire7368 ) | ( n_n1454  &  n_n416  &  wire7356 ) ;
 assign wire7371 = ( wire1367 ) | ( wire7366 ) | ( wire7367 ) ;
 assign wire7383 = ( wire1356 ) | ( wire1357 ) | ( wire7379 ) | ( wire7380 ) ;
 assign n_n1827 = ( n_n1862 ) | ( wire7370 ) | ( wire7371 ) | ( wire7383 ) ;
 assign n_n1870 = ( wire1337 ) | ( wire7400 ) | ( n_n1489  &  wire784 ) ;
 assign wire627 = ( wire1330 ) | ( wire52  &  wire223 ) | ( wire52  &  wire261 ) ;
 assign n_n1829 = ( n_n1870 ) | ( wire1347 ) | ( _439 ) | ( _10790 ) ;
 assign wire7432 = ( wire1308 ) | ( n_n284  &  wire75 ) ;
 assign wire7433 = ( wire1309 ) | ( n_n300  &  wire654 ) ;
 assign wire7441 = ( _10830 ) | ( _10831 ) ;
 assign wire990 = ( n_n416  &  n_n1300  &  wire457 ) | ( n_n1300  &  n_n706  &  wire457 ) ;
 assign wire991 = ( (~ i_24_)  &  wire297  &  wire7716 ) | ( (~ i_24_)  &  wire1406  &  wire7716 ) ;
 assign wire992 = ( n_n805  &  wire994 ) | ( n_n805  &  n_n1302  &  n_n849 ) ;
 assign wire993 = ( wire7547  &  wire996  &  _9996 ) | ( wire7547  &  wire7718  &  _9996 ) ;
 assign n_n1866 = ( wire990 ) | ( wire991 ) | ( wire992 ) | ( wire993 ) ;
 assign wire983 = ( n_n1197  &  wire988  &  _10721 ) | ( n_n1197  &  _10721  &  _10722 ) ;
 assign wire987 = ( n_n805  &  n_n1466  &  n_n849 ) ;
 assign wire7727 = ( _510 ) | ( n_n805  &  wire7725  &  _10003 ) ;
 assign wire7728 = ( (~ i_10_)  &  wire310 ) | ( n_n316  &  wire7726 ) ;
 assign n_n1865 = ( wire983 ) | ( wire987 ) | ( wire7727 ) | ( wire7728 ) ;
 assign wire7771 = ( wire953 ) | ( _11016 ) ;
 assign n_n1548 = ( wire7866 ) | ( _282 ) | ( _283 ) | ( _11093 ) ;
 assign n_n1545 = ( wire8052 ) | ( wire8054 ) | ( _11294 ) ;
 assign wire7923 = ( wire7853 ) | ( wire7921 ) | ( _11388 ) ;
 assign wire8079 = ( n_n1556 ) | ( n_n1582 ) | ( n_n1584 ) | ( wire8077 ) ;
 assign wire232 = ( (~ i_9_)  &  (~ i_5_)  &  (~ i_6_)  &  (~ i_4_) ) ;
 assign n_n1443 = ( (~ i_13_)  &  (~ i_17_)  &  (~ i_16_) ) ;
 assign wire79 = ( (~ i_27_)  &  (~ i_26_)  &  (~ i_24_)  &  i_36_ ) ;
 assign n_n460 = ( (~ i_28_)  &  (~ i_32_)  &  i_29_ ) ;
 assign wire462 = ( n_n1443  &  wire79  &  n_n460 ) ;
 assign wire227 = ( (~ i_32_)  &  (~ i_34_)  &  i_36_  &  i_35_ ) ;
 assign wire493 = ( (~ i_27_)  &  (~ i_28_)  &  (~ i_29_)  &  wire227 ) ;
 assign wire58 = ( (~ i_28_)  &  (~ i_26_) ) ;
 assign n_n1441 = ( (~ i_27_)  &  (~ i_28_)  &  (~ i_26_) ) ;
 assign wire43 = ( (~ i_13_)  &  (~ i_16_) ) ;
 assign wire302 = ( (~ i_32_)  &  (~ i_31_) ) ;
 assign n_n1433 = ( (~ i_32_)  &  (~ i_31_)  &  i_34_ ) ;
 assign n_n1425 = ( (~ i_30_)  &  (~ i_28_)  &  (~ i_26_) ) ;
 assign wire54 = ( (~ i_23_)  &  (~ i_24_) ) ;
 assign n_n1396 = ( i_25_  &  (~ i_23_)  &  (~ i_24_) ) ;
 assign wire10 = ( (~ i_14_)  &  (~ i_16_) ) ;
 assign n_n1404 = ( (~ i_14_)  &  (~ i_12_)  &  (~ i_16_) ) ;
 assign n_n1390 = ( (~ i_23_)  &  (~ i_24_)  &  (~ i_16_) ) ;
 assign wire415 = ( (~ i_14_)  &  (~ i_12_) ) ;
 assign n_n1372 = ( i_7_  &  (~ i_14_)  &  (~ i_12_) ) ;
 assign n_n1369 = ( (~ i_27_)  &  (~ i_26_)  &  (~ i_24_) ) ;
 assign n_n1429 = ( (~ i_13_)  &  (~ i_12_)  &  (~ i_16_) ) ;
 assign n_n1454 = ( (~ i_25_)  &  (~ i_26_)  &  (~ i_24_) ) ;
 assign n_n1489 = ( (~ i_30_)  &  (~ i_28_)  &  (~ i_29_) ) ;
 assign n_n1353 = ( i_9_  &  (~ i_10_)  &  (~ i_8_) ) ;
 assign n_n1361 = ( (~ i_35_)  &  i_38_ ) ;
 assign n_n1423 = ( (~ i_28_)  &  (~ i_25_)  &  (~ i_24_) ) ;
 assign n_n1295 = ( i_34_  &  i_37_ ) ;
 assign n_n1439 = ( (~ i_28_)  &  (~ i_24_)  &  (~ i_29_) ) ;
 assign wire3 = ( i_30_ ) | ( i_32_ ) ;
 assign n_n1438 = ( (~ i_30_)  &  (~ i_32_)  &  (~ i_31_) ) ;
 assign n_n1397 = ( (~ i_34_)  &  i_35_ ) ;
 assign n_n1274 = ( (~ i_20_)  &  (~ i_23_)  &  (~ i_17_) ) ;
 assign n_n1334 = ( i_31_  &  i_34_ ) ;
 assign n_n1368 = ( (~ i_28_)  &  i_29_ ) ;
 assign n_n1216 = ( (~ i_27_)  &  (~ i_28_)  &  (~ i_24_) ) ;
 assign wire290 = ( (~ i_13_)  &  (~ i_12_) ) ;
 assign n_n1391 = ( i_7_  &  (~ i_13_)  &  (~ i_12_) ) ;
 assign n_n1478 = ( (~ i_28_)  &  (~ i_25_)  &  (~ i_26_) ) ;
 assign n_n1307 = ( (~ i_5_)  &  (~ i_4_)  &  (~ i_2_) ) ;
 assign n_n1374 = ( i_34_  &  i_33_ ) ;
 assign n_n805 = ( i_34_  &  (~ i_35_)  &  i_38_ ) ;
 assign n_n1504 = ( i_31_  &  (~ i_34_)  &  i_35_ ) ;
 assign n_n841 = ( (~ i_9_)  &  (~ i_8_)  &  (~ i_6_) ) ;
 assign n_n853 = ( (~ i_9_)  &  (~ i_10_)  &  (~ i_6_) ) ;
 assign n_n793 = ( (~ i_27_)  &  (~ i_28_)  &  (~ i_23_) ) ;
 assign n_n1315 = ( (~ i_9_)  &  i_7_  &  (~ i_12_) ) ;
 assign n_n1092 = ( i_20_  &  (~ i_23_)  &  (~ i_21_) ) ;
 assign n_n1406 = ( (~ i_27_)  &  (~ i_28_)  &  i_29_ ) ;
 assign n_n1466 = ( (~ i_28_)  &  (~ i_25_)  &  (~ i_29_) ) ;
 assign wire224 = ( (~ i_5_)  &  (~ i_6_) ) ;
 assign n_n1278 = ( (~ i_7_)  &  (~ i_5_)  &  (~ i_6_) ) ;
 assign n_n787 = ( i_3_  &  (~ i_4_)  &  (~ i_2_) ) ;
 assign n_n1197 = ( (~ i_33_)  &  (~ i_35_)  &  i_38_ ) ;
 assign n_n762 = ( (~ i_30_)  &  (~ i_32_)  &  n_n1197 ) ;
 assign n_n1038 = ( i_9_  &  (~ i_8_)  &  (~ i_3_) ) ;
 assign n_n1314 = ( (~ i_13_)  &  (~ i_23_)  &  (~ i_16_) ) ;
 assign n_n1375 = ( (~ i_27_)  &  (~ i_28_)  &  (~ i_29_) ) ;
 assign wire13 = ( (~ i_7_)  &  (~ i_8_) ) ;
 assign n_n1141 = ( (~ i_7_)  &  (~ i_8_)  &  (~ i_12_) ) ;
 assign wire7086 = ( (~ i_13_)  &  (~ i_23_)  &  (~ i_24_)  &  (~ i_16_) ) ;
 assign n_n544 = ( (~ i_6_)  &  (~ i_12_)  &  n_n1307  &  wire7086 ) ;
 assign n_n1486 = ( (~ i_28_)  &  (~ i_26_)  &  (~ i_29_) ) ;
 assign n_n1408 = ( (~ i_14_)  &  (~ i_17_)  &  (~ i_16_) ) ;
 assign n_n1318 = ( (~ i_35_)  &  i_37_ ) ;
 assign n_n504 = ( (~ i_33_)  &  (~ i_35_)  &  i_37_ ) ;
 assign wire404 = ( (~ i_9_)  &  i_3_  &  (~ i_4_)  &  (~ i_2_) ) ;
 assign wire297 = ( wire404  &  _10475 ) ;
 assign n_n416 = ( (~ i_8_)  &  (~ i_18_)  &  n_n1278  &  wire404 ) ;
 assign n_n1305 = ( (~ i_32_)  &  (~ i_33_)  &  (~ i_29_) ) ;
 assign n_n1118 = ( (~ i_8_)  &  (~ i_5_)  &  (~ i_6_) ) ;
 assign n_n1279 = ( (~ i_4_)  &  (~ i_1_)  &  (~ i_2_) ) ;
 assign n_n358 = ( n_n1278  &  n_n1408  &  n_n1279 ) ;
 assign n_n1048 = ( i_9_  &  (~ i_13_)  &  i_18_ ) ;
 assign n_n1144 = ( (~ i_8_)  &  (~ i_6_)  &  (~ i_12_) ) ;
 assign n_n307 = ( n_n1307  &  n_n1048  &  n_n1144 ) ;
 assign n_n1263 = ( (~ i_14_)  &  (~ i_23_)  &  (~ i_16_) ) ;
 assign n_n1306 = ( (~ i_7_)  &  (~ i_6_)  &  (~ i_12_) ) ;
 assign n_n620 = ( n_n1307  &  n_n1263  &  n_n1306 ) ;
 assign n_n1288 = ( (~ i_28_)  &  (~ i_32_)  &  (~ i_29_) ) ;
 assign n_n1018 = ( (~ i_27_)  &  (~ i_23_)  &  (~ i_24_) ) ;
 assign n_n1400 = ( (~ i_23_)  &  (~ i_24_)  &  (~ i_17_) ) ;
 assign n_n819 = ( i_9_  &  (~ i_5_)  &  (~ i_6_) ) ;
 assign wire7419 = ( (~ i_3_)  &  (~ i_13_)  &  (~ i_12_) ) ;
 assign wire7425 = ( i_9_  &  (~ i_5_)  &  (~ i_6_)  &  i_11_ ) ;
 assign n_n394 = ( (~ i_4_)  &  (~ i_2_)  &  wire7419  &  wire7425 ) ;
 assign n_n458 = ( n_n1443  &  n_n1278  &  n_n1279 ) ;
 assign wire7426 = ( i_9_  &  (~ i_13_)  &  i_11_  &  i_18_ ) ;
 assign n_n391 = ( (~ i_6_)  &  (~ i_12_)  &  n_n1307  &  wire7426 ) ;
 assign n_n1055 = ( i_9_  &  (~ i_13_)  &  i_11_ ) ;
 assign n_n461 = ( (~ i_5_)  &  (~ i_6_)  &  (~ i_4_) ) ;
 assign wire7411 = ( (~ i_3_)  &  (~ i_1_)  &  (~ i_2_) ) ;
 assign n_n372 = ( n_n1055  &  n_n461  &  wire7411 ) ;
 assign n_n1179 = ( (~ i_32_)  &  (~ i_35_)  &  i_38_ ) ;
 assign wire7265 = ( (~ i_28_)  &  (~ i_25_)  &  (~ i_26_) ) ;
 assign wire257 = ( (~ i_24_)  &  (~ i_22_)  &  wire7265 ) ;
 assign n_n300 = ( (~ i_24_)  &  (~ i_22_)  &  n_n1179  &  wire7265 ) ;
 assign n_n1225 = ( (~ i_28_)  &  i_34_  &  (~ i_29_) ) ;
 assign wire7412 = ( i_9_  &  (~ i_13_)  &  i_19_ ) ;
 assign n_n294 = ( n_n461  &  wire7411  &  wire7412 ) ;
 assign n_n301 = ( (~ i_10_)  &  (~ i_13_)  &  (~ i_16_) ) ;
 assign n_n880 = ( i_36_  &  (~ i_35_) ) ;
 assign n_n1100 = ( (~ i_9_)  &  (~ i_7_)  &  (~ i_6_) ) ;
 assign wire51 = ( (~ i_5_)  &  (~ i_6_)  &  n_n1279 ) ;
 assign wire260 = ( (~ i_14_)  &  (~ i_23_)  &  (~ i_17_)  &  (~ i_16_) ) ;
 assign n_n437 = ( (~ i_5_)  &  (~ i_6_)  &  n_n1279  &  wire260 ) ;
 assign n_n571 = ( i_35_  &  i_37_ ) ;
 assign n_n1258 = ( (~ i_27_)  &  (~ i_23_)  &  (~ i_17_) ) ;
 assign wire263 = ( (~ i_17_)  &  (~ i_16_) ) ;
 assign n_n825 = ( (~ i_17_)  &  (~ i_21_)  &  (~ i_16_) ) ;
 assign n_n1437 = ( i_34_  &  (~ i_33_)  &  (~ i_35_) ) ;
 assign n_n1340 = ( (~ i_32_)  &  i_34_  &  (~ i_33_) ) ;
 assign n_n180 = ( (~ i_9_)  &  (~ i_13_)  &  (~ i_16_) ) ;
 assign n_n132 = ( (~ i_18_)  &  (~ i_17_)  &  (~ i_16_) ) ;
 assign n_n152 = ( (~ i_4_)  &  (~ i_1_)  &  (~ i_0_) ) ;
 assign n_n1300 = ( (~ i_33_)  &  i_38_ ) ;
 assign n_n1472 = ( (~ i_30_)  &  (~ i_32_)  &  (~ i_29_) ) ;
 assign wire50 = ( (~ i_4_)  &  (~ i_1_)  &  (~ i_2_)  &  _9992 ) ;
 assign wire52 = ( (~ i_28_)  &  (~ i_22_)  &  n_n1454 ) ;
 assign wire85 = ( (~ i_9_)  &  (~ i_7_)  &  (~ i_6_)  &  _9748 ) ;
 assign n_n1303 = ( (~ i_7_)  &  (~ i_8_)  &  (~ i_6_) ) ;
 assign wire223 = ( (~ i_9_)  &  (~ i_10_)  &  n_n1307  &  n_n1303 ) ;
 assign wire264 = ( (~ i_31_)  &  (~ i_35_)  &  i_38_ ) ;
 assign wire61 = ( (~ i_28_)  &  (~ i_26_)  &  (~ i_24_)  &  (~ i_22_) ) ;
 assign wire388 = ( (~ i_33_)  &  i_38_  &  wire61 ) ;
 assign wire446 = ( (~ i_32_)  &  (~ i_31_)  &  (~ i_35_)  &  i_38_ ) ;
 assign wire262 = ( i_9_  &  (~ i_3_)  &  (~ i_13_)  &  i_11_ ) ;
 assign wire18 = ( i_9_  &  (~ i_3_)  &  (~ i_13_) ) | ( i_9_  &  (~ i_13_)  &  i_18_ ) ;
 assign wire436 = ( i_9_  &  (~ i_13_)  &  i_11_  &  i_18_ ) ;
 assign wire529 = ( wire262 ) | ( wire436 ) | ( i_19_  &  wire18 ) ;
 assign wire7511 = ( _781 ) | ( _782 ) ;
 assign wire7512 = ( wire223  &  wire388 ) | ( wire50  &  wire7510 ) ;
 assign n_n1147 = ( (~ i_7_)  &  (~ i_13_)  &  (~ i_12_) ) ;
 assign n_n1089 = ( (~ i_7_)  &  (~ i_14_)  &  (~ i_12_) ) ;
 assign wire298 = ( (~ i_24_)  &  i_34_ ) ;
 assign wire244 = ( i_34_  &  i_36_ ) ;
 assign wire7789 = ( (~ i_30_)  &  (~ i_7_)  &  (~ i_32_) ) ;
 assign wire410 = ( n_n1375  &  n_n1400  &  wire244  &  wire7789 ) ;
 assign wire7785 = ( (~ i_7_)  &  i_36_ ) ;
 assign wire516 = ( n_n1441  &  n_n1400  &  n_n1472  &  wire7785 ) ;
 assign n_n1322 = ( (~ i_23_)  &  (~ i_17_)  &  (~ i_16_) ) ;
 assign wire7243 = ( (~ i_7_)  &  (~ i_8_)  &  (~ i_13_) ) ;
 assign wire530 = ( n_n1314  &  n_n1141 ) | ( n_n1322  &  wire7243 ) ;
 assign wire935 = ( _62 ) | ( _63 ) ;
 assign wire7793 = ( wire933 ) | ( n_n1216  &  wire530  &  wire7784 ) ;
 assign wire7794 = ( wire937 ) | ( (~ i_14_)  &  (~ i_16_)  &  wire516 ) ;
 assign wire7795 = ( wire939 ) | ( (~ i_13_)  &  (~ i_16_)  &  wire410 ) ;
 assign n_n1580 = ( wire935 ) | ( wire7793 ) | ( wire7794 ) | ( wire7795 ) ;
 assign n_n1326 = ( (~ i_28_)  &  (~ i_34_)  &  i_29_ ) ;
 assign wire245 = ( (~ i_23_)  &  (~ i_24_)  &  i_21_  &  i_34_ ) ;
 assign wire277 = ( (~ i_30_)  &  (~ i_28_) ) ;
 assign wire340 = ( i_14_  &  (~ i_32_)  &  (~ i_31_)  &  i_33_ ) ;
 assign n_n1213 = ( (~ i_26_)  &  (~ i_23_)  &  (~ i_24_) ) ;
 assign wire533 = ( (~ i_13_)  &  (~ i_12_)  &  (~ i_16_) ) | ( (~ i_13_)  &  (~ i_17_)  &  (~ i_16_) ) ;
 assign n_n1323 = ( (~ i_9_)  &  i_7_  &  (~ i_13_) ) ;
 assign wire532 = ( wire43  &  n_n1315 ) | ( wire263  &  n_n1323 ) ;
 assign wire7806 = ( wire926 ) | ( wire532  &  n_n1511  &  wire7802 ) ;
 assign wire7807 = ( wire928 ) | ( (~ i_14_)  &  (~ i_16_)  &  wire410 ) ;
 assign wire7808 = ( wire924 ) | ( wire925 ) | ( _43 ) ;
 assign n_n1579 = ( wire7806 ) | ( wire7807 ) | ( wire7808 ) ;
 assign wire80 = ( (~ i_27_)  &  (~ i_28_)  &  (~ i_24_)  &  (~ i_29_) ) ;
 assign wire536 = ( n_n1314  &  n_n1141 ) | ( n_n1322  &  wire7243 ) ;
 assign n_n1285 = ( (~ i_9_)  &  i_7_  &  (~ i_14_) ) ;
 assign wire535 = ( n_n1315  &  n_n1263 ) | ( n_n1322  &  n_n1285 ) ;
 assign wire918 = ( n_n1406  &  n_n1213  &  _9325  &  _11482 ) ;
 assign wire7812 = ( wire535  &  wire7810 ) | ( wire536  &  wire7811 ) ;
 assign wire7813 = ( wire919 ) | ( (~ i_13_)  &  (~ i_16_)  &  wire516 ) ;
 assign n_n1581 = ( wire7812 ) | ( wire7813 ) | ( _11489 ) ;
 assign n_n1519 = ( i_12_  &  (~ i_24_)  &  i_17_ ) ;
 assign n_n1419 = ( (~ i_34_)  &  i_35_  &  i_38_ ) ;
 assign n_n1302 = ( (~ i_28_)  &  (~ i_33_)  &  (~ i_29_) ) ;
 assign n_n1401 = ( i_7_  &  (~ i_13_)  &  (~ i_16_) ) ;
 assign wire283 = ( (~ i_8_)  &  (~ i_2_) ) ;
 assign n_n1192 = ( i_9_  &  (~ i_8_)  &  (~ i_2_) ) ;
 assign n_n1257 = ( (~ i_28_)  &  i_33_  &  (~ i_29_) ) ;
 assign n_n1133 = ( (~ i_32_)  &  (~ i_31_)  &  (~ i_29_) ) ;
 assign n_n1128 = ( (~ i_28_)  &  (~ i_31_)  &  (~ i_29_) ) ;
 assign n_n586 = ( (~ i_13_)  &  i_12_  &  i_11_ ) ;
 assign n_n1523 = ( (~ i_26_)  &  (~ i_24_)  &  (~ i_22_) ) ;
 assign n_n269 = ( n_n1307  &  n_n1314  &  n_n1306 ) ;
 assign wire259 = ( (~ i_8_)  &  (~ i_13_)  &  (~ i_16_) ) ;
 assign n_n242 = ( n_n1278  &  n_n1279  &  wire259 ) ;
 assign n_n1202 = ( (~ i_32_)  &  (~ i_34_)  &  i_35_ ) ;
 assign wire258 = ( (~ i_8_)  &  (~ i_14_)  &  (~ i_16_) ) ;
 assign n_n355 = ( n_n1278  &  n_n1279  &  wire258 ) ;
 assign n_n1345 = ( (~ i_30_)  &  (~ i_28_)  &  (~ i_31_) ) ;
 assign wire7413 = ( (~ i_13_)  &  i_11_  &  i_18_ ) ;
 assign n_n371 = ( n_n1279  &  n_n819  &  wire7413 ) ;
 assign n_n316 = ( (~ i_28_)  &  (~ i_32_)  &  n_n1197  &  n_n1523 ) ;
 assign n_n735 = ( (~ i_13_)  &  i_18_  &  i_19_ ) ;
 assign wire7423 = ( i_9_  &  (~ i_13_)  &  i_18_  &  i_19_ ) ;
 assign n_n315 = ( (~ i_6_)  &  (~ i_12_)  &  n_n1307  &  wire7423 ) ;
 assign n_n984 = ( (~ i_27_)  &  (~ i_28_)  &  i_31_ ) ;
 assign n_n1458 = ( (~ i_32_)  &  (~ i_33_)  &  (~ i_35_) ) ;
 assign n_n177 = ( (~ i_23_)  &  (~ i_17_)  &  (~ i_19_) ) ;
 assign n_n1241 = ( i_34_  &  (~ i_33_)  &  (~ i_29_) ) ;
 assign n_n179 = ( (~ i_23_)  &  (~ i_18_)  &  (~ i_17_) ) ;
 assign n_n245 = ( (~ i_5_)  &  (~ i_4_)  &  (~ i_0_) ) ;
 assign n_n1431 = ( (~ i_30_)  &  (~ i_28_)  &  (~ i_32_) ) ;
 assign wire7491 = ( i_20_  &  (~ i_21_)  &  (~ i_22_) ) ;
 assign wire7266 = ( (~ i_28_)  &  (~ i_33_)  &  i_38_ ) ;
 assign wire70 = ( (~ i_28_)  &  (~ i_33_)  &  i_38_  &  _10425 ) ;
 assign wire7492 = ( (~ i_8_)  &  (~ i_24_)  &  i_38_ ) ;
 assign wire212 = ( n_n1278  &  n_n1279  &  wire7492 ) ;
 assign wire239 = ( (~ i_25_)  &  (~ i_24_)  &  i_38_ ) ;
 assign wire288 = ( (~ i_28_)  &  i_34_  &  (~ i_33_)  &  (~ i_29_) ) ;
 assign wire539 = ( (~ i_13_)  &  (~ i_12_)  &  (~ i_16_) ) | ( (~ i_13_)  &  (~ i_17_)  &  (~ i_16_) ) ;
 assign wire7409 = ( (~ i_32_)  &  i_34_  &  (~ i_29_) ) ;
 assign wire537 = ( n_n1439  &  n_n1340 ) | ( n_n1423  &  wire7409 ) ;
 assign wire7494 = ( wire1234 ) | ( n_n1279  &  wire537  &  _10176 ) ;
 assign wire7495 = ( wire1235 ) | ( _626 ) | ( _627 ) ;
 assign n_n1881 = ( wire7494 ) | ( wire7495 ) | ( wire1230 ) | ( _635 ) ;
 assign n_n576 = ( (~ i_32_)  &  i_36_  &  (~ i_35_) ) ;
 assign n_n1499 = ( (~ i_28_)  &  i_31_  &  (~ i_29_) ) ;
 assign wire47 = ( (~ i_23_)  &  (~ i_34_)  &  i_35_ ) ;
 assign wire44 = ( (~ i_27_)  &  (~ i_28_)  &  (~ i_26_)  &  i_29_ ) ;
 assign wire7749 = ( (~ i_23_)  &  (~ i_24_)  &  (~ i_21_) ) ;
 assign wire7847 = ( (~ i_5_)  &  (~ i_6_)  &  (~ i_4_)  &  (~ i_31_) ) ;
 assign wire307 = ( n_n576  &  wire44  &  wire7749  &  wire7847 ) ;
 assign wire541 = ( (~ i_13_)  &  (~ i_12_)  &  (~ i_16_) ) | ( (~ i_13_)  &  (~ i_17_)  &  (~ i_16_) ) ;
 assign n_n329 = ( (~ i_5_)  &  (~ i_6_)  &  n_n1279  &  wire6920 ) ;
 assign wire468 = ( (~ i_28_)  &  (~ i_31_)  &  (~ i_29_)  &  _11325 ) ;
 assign wire67 = ( (~ i_26_)  &  (~ i_23_)  &  (~ i_24_)  &  _11027 ) ;
 assign wire367 = ( n_n1443  &  n_n1307  &  n_n853 ) ;
 assign wire540 = ( n_n329  &  wire468 ) | ( wire67  &  wire367 ) ;
 assign n_n195 = ( n_n1408  &  n_n1118  &  n_n1279 ) ;
 assign wire864 = ( i_36_  &  wire7871 ) | ( wire7868  &  _11037 ) ;
 assign wire7874 = ( wire500  &  wire312 ) | ( n_n437  &  wire7867 ) ;
 assign wire7875 = ( n_n1404  &  wire307 ) | ( n_n329  &  wire483 ) ;
 assign wire86 = ( i_34_  &  i_36_  &  (~ i_35_) ) ;
 assign wire275 = ( (~ i_23_)  &  (~ i_34_)  &  i_35_  &  _11077 ) ;
 assign wire483 = ( n_n1216  &  n_n1133  &  wire86 ) ;
 assign wire500 = ( n_n1018  &  n_n1128  &  wire86 ) ;
 assign wire41 = ( (~ i_9_)  &  (~ i_8_)  &  (~ i_6_)  &  _9494 ) ;
 assign wire221 = ( (~ i_27_)  &  (~ i_23_)  &  (~ i_24_)  &  _9480 ) ;
 assign wire495 = ( n_n1307  &  n_n1408  &  n_n839 ) ;
 assign wire7189 = ( n_n1375  &  n_n1400  &  n_n916 ) ;
 assign wire543 = ( wire221  &  wire495 ) | ( wire41  &  wire7189 ) ;
 assign wire7866 = ( wire875 ) | ( wire7864 ) | ( wire559  &  wire7856 ) ;
 assign wire7916 = ( n_n358  &  wire7910 ) | ( n_n263  &  wire7912 ) ;
 assign wire7917 = ( wire493  &  n_n269 ) | ( wire360  &  wire7911 ) ;
 assign wire7920 = ( wire7918 ) | ( n_n880  &  wire829 ) | ( n_n880  &  wire7915 ) ;
 assign n_n1497 = ( (~ i_28_)  &  (~ i_26_)  &  (~ i_24_) ) ;
 assign n_n1384 = ( i_14_  &  (~ i_13_)  &  (~ i_12_) ) ;
 assign n_n1393 = ( (~ i_32_)  &  (~ i_31_)  &  i_33_ ) ;
 assign n_n1282 = ( (~ i_23_)  &  (~ i_17_)  &  (~ i_21_) ) ;
 assign n_n839 = ( (~ i_9_)  &  (~ i_6_)  &  i_13_ ) ;
 assign n_n1311 = ( (~ i_32_)  &  (~ i_34_)  &  (~ i_33_) ) ;
 assign n_n263 = ( n_n1429  &  n_n1307  &  n_n1303 ) ;
 assign n_n363 = ( n_n1404  &  n_n1307  &  n_n1303 ) ;
 assign n_n584 = ( (~ i_13_)  &  i_12_  &  i_18_ ) ;
 assign n_n1033 = ( i_9_  &  (~ i_8_)  &  i_11_ ) ;
 assign wire7420 = ( i_9_  &  (~ i_8_)  &  (~ i_5_)  &  (~ i_6_) ) ;
 assign n_n309 = ( (~ i_4_)  &  (~ i_2_)  &  wire7419  &  wire7420 ) ;
 assign wire7424 = ( i_9_  &  (~ i_5_)  &  (~ i_6_)  &  i_19_ ) ;
 assign n_n317 = ( (~ i_4_)  &  (~ i_2_)  &  wire7419  &  wire7424 ) ;
 assign n_n712 = ( i_10_  &  i_7_  &  (~ i_11_) ) ;
 assign n_n284 = ( n_n1279  &  n_n819  &  n_n735 ) ;
 assign n_n1028 = ( i_9_  &  (~ i_8_)  &  (~ i_13_) ) ;
 assign n_n178 = ( (~ i_13_)  &  (~ i_11_)  &  (~ i_16_) ) ;
 assign wire57 = ( (~ i_30_)  &  (~ i_29_) ) ;
 assign wire77 = ( (~ i_30_)  &  (~ i_7_)  &  (~ i_8_) ) ;
 assign wire83 = ( (~ i_28_)  &  i_22_ ) ;
 assign wire372 = ( (~ i_28_)  &  (~ i_34_)  &  i_35_  &  i_29_ ) ;
 assign wire380 = ( (~ i_33_)  &  i_38_  &  n_n1486 ) ;
 assign wire71 = ( (~ i_28_)  &  (~ i_25_)  &  (~ i_26_)  &  (~ i_29_) ) ;
 assign wire395 = ( (~ i_24_)  &  i_38_  &  wire71 ) ;
 assign wire503 = ( (~ i_26_)  &  (~ i_24_)  &  (~ i_33_)  &  i_38_ ) ;
 assign n_n1387 = ( i_14_  &  (~ i_13_)  &  (~ i_16_) ) ;
 assign n_n1359 = ( i_9_  &  (~ i_10_)  &  (~ i_24_) ) ;
 assign n_n1080 = ( (~ i_27_)  &  (~ i_23_)  &  i_21_ ) ;
 assign n_n1254 = ( (~ i_23_)  &  (~ i_21_)  &  (~ i_16_) ) ;
 assign wire196 = ( n_n1489  &  n_n1393  &  wire1649 ) | ( n_n1489  &  n_n1393  &  wire1650 ) ;
 assign wire7926 = ( n_n1438  &  wire6948  &  wire6949 ) | ( n_n1438  &  wire6948  &  wire7653 ) ;
 assign wire7927 = ( wire813 ) | ( n_n1374  &  n_n1375  &  wire38 ) ;
 assign n_n1585 = ( wire7927 ) | ( _96 ) | ( _97 ) | ( _11400 ) ;
 assign n_n1422 = ( (~ i_32_)  &  i_34_  &  (~ i_35_) ) ;
 assign wire8 = ( (~ i_14_)  &  (~ i_12_)  &  (~ i_16_) ) | ( (~ i_14_)  &  (~ i_17_)  &  (~ i_16_) ) ;
 assign wire38 = ( n_n1390  &  n_n1384 ) | ( n_n1400  &  n_n1387 ) ;
 assign wire1661 = ( n_n1406  &  wire802  &  wire7025 ) ;
 assign wire7682 = ( (~ i_23_)  &  (~ i_24_)  &  i_34_ ) ;
 assign wire112 = ( n_n1489  &  wire340  &  wire7682 ) ;
 assign wire7029 = ( (~ i_30_)  &  i_22_  &  (~ i_32_)  &  (~ i_31_) ) ;
 assign wire127 = ( wire372  &  wire7029 ) ;
 assign wire546 = ( (~ i_14_)  &  (~ i_12_)  &  (~ i_16_) ) | ( (~ i_14_)  &  (~ i_17_)  &  (~ i_16_) ) ;
 assign wire7938 = ( wire494 ) | ( wire497 ) | ( wire7935 ) | ( wire7936 ) ;
 assign n_n1556 = ( n_n1585 ) | ( wire1661 ) | ( wire7938 ) | ( _90 ) ;
 assign n_n1459 = ( (~ i_30_)  &  (~ i_31_)  &  (~ i_29_) ) ;
 assign n_n1377 = ( i_7_  &  (~ i_14_)  &  (~ i_16_) ) ;
 assign n_n1312 = ( (~ i_23_)  &  (~ i_24_)  &  i_21_ ) ;
 assign n_n820 = ( (~ i_30_)  &  (~ i_34_)  &  i_36_  &  i_35_ ) ;
 assign n_n706 = ( n_n1307  &  n_n1303  &  _10469 ) ;
 assign wire205 = ( (~ i_24_)  &  (~ i_22_) ) ;
 assign n_n1191 = ( (~ i_10_)  &  (~ i_24_)  &  (~ i_22_) ) ;
 assign wire7051 = ( (~ i_14_)  &  (~ i_23_)  &  (~ i_24_)  &  (~ i_16_) ) ;
 assign n_n608 = ( (~ i_6_)  &  (~ i_12_)  &  n_n1307  &  wire7051 ) ;
 assign n_n1058 = ( i_9_  &  (~ i_3_)  &  i_11_ ) ;
 assign n_n916 = ( (~ i_14_)  &  i_13_  &  (~ i_16_) ) ;
 assign n_n629 = ( (~ i_20_)  &  (~ i_17_)  &  (~ i_16_) ) ;
 assign wire12 = ( (~ i_24_)  &  (~ i_35_)  &  i_38_ ) ;
 assign n_n338 = ( i_19_  &  wire288  &  wire12 ) ;
 assign wire261 = ( (~ i_9_)  &  i_13_  &  n_n1307  &  n_n1303 ) ;
 assign n_n129 = ( n_n1307  &  n_n1303  &  _9781 ) ;
 assign n_n26 = ( i_3_  &  (~ i_4_)  &  (~ i_0_) ) ;
 assign wire463 = ( n_n1443  &  n_n1369  &  _10985 ) ;
 assign wire966 = ( n_n1375  &  n_n1322  &  _9686  &  _10995 ) ;
 assign wire967 = ( wire273  &  wire1766 ) | ( n_n129  &  n_n130  &  wire273 ) ;
 assign wire338 = ( (~ i_5_)  &  i_3_  &  (~ i_4_)  &  (~ i_18_) ) ;
 assign wire7753 = ( (~ i_8_)  &  (~ i_11_)  &  (~ i_19_) ) ;
 assign wire547 = ( n_n841  &  wire338 ) | ( wire232  &  wire7753 ) ;
 assign wire451 = ( (~ i_14_)  &  wire517 ) | ( (~ i_14_)  &  wire65  &  wire7945 ) ;
 assign wire7952 = ( wire299  &  wire572 ) | ( wire342  &  wire7941 ) ;
 assign wire7953 = ( wire471 ) | ( n_n1429  &  wire478 ) ;
 assign wire7954 = ( wire469 ) | ( wire7947  &  _11227 ) ;
 assign n_n1574 = ( wire451 ) | ( wire7952 ) | ( wire7953 ) | ( wire7954 ) ;
 assign wire412 = ( (~ i_13_)  &  wire517 ) | ( (~ i_13_)  &  wire65  &  wire7961 ) ;
 assign wire7963 = ( wire7957  &  wire7958 ) | ( wire385  &  wire7959 ) ;
 assign wire7964 = ( wire417 ) | ( n_n1375  &  n_n1400  &  wire7960 ) ;
 assign wire7965 = ( wire424 ) | ( n_n1375  &  wire427 ) | ( n_n1375  &  wire439 ) ;
 assign n_n1575 = ( wire412 ) | ( wire7963 ) | ( wire7964 ) | ( wire7965 ) ;
 assign wire7979 = ( wire350 ) | ( n_n1213  &  n_n984  &  wire608 ) ;
 assign wire7981 = ( wire339 ) | ( (~ i_13_)  &  (~ i_16_)  &  wire301 ) ;
 assign n_n1578 = ( wire7979 ) | ( wire7981 ) | ( _11146 ) ;
 assign wire195 = ( n_n880  &  n_n1459  &  wire200 ) | ( n_n880  &  n_n1459  &  wire201 ) ;
 assign wire7989 = ( wire192 ) | ( wire194 ) ;
 assign wire7990 = ( wire197 ) | ( n_n1375  &  n_n1400  &  wire7986 ) ;
 assign wire7991 = ( wire198 ) | ( (~ i_14_)  &  (~ i_16_)  &  wire301 ) ;
 assign n_n1576 = ( wire195 ) | ( wire7989 ) | ( wire7990 ) | ( wire7991 ) ;
 assign wire8003 = ( wire184 ) | ( wire187 ) | ( wire74  &  wire7994 ) ;
 assign n_n1577 = ( wire8003 ) | ( wire183 ) | ( wire185 ) | ( _180 ) ;
 assign wire174 = ( i_36_  &  wire8007 ) | ( n_n363  &  _11094 ) ;
 assign wire176 = ( wire7053  &  wire8008  &  _9404  &  _11097 ) ;
 assign wire8035 = ( wire8029  &  wire8030 ) | ( wire723  &  wire8031 ) ;
 assign wire8036 = ( wire160 ) | ( wire79  &  n_n1288  &  n_n269 ) ;
 assign wire8037 = ( wire158 ) | ( wire161 ) | ( wire724  &  wire8028 ) ;
 assign n_n1573 = ( wire8035 ) | ( wire8036 ) | ( wire8037 ) ;
 assign wire8046 = ( n_n1404  &  wire478 ) | ( n_n263  &  wire8041 ) ;
 assign wire8047 = ( wire142 ) | ( wire150 ) | ( wire731  &  wire8039 ) ;
 assign n_n1572 = ( wire8046 ) | ( wire8047 ) | ( _221 ) ;
 assign wire8052 = ( n_n1572 ) | ( wire164 ) | ( wire8023 ) | ( wire8026 ) ;
 assign wire8054 = ( n_n1574 ) | ( n_n1575 ) | ( n_n1577 ) | ( n_n1573 ) ;
 assign n_n1251 = ( (~ i_27_)  &  (~ i_23_)  &  (~ i_16_) ) ;
 assign n_n998 = ( (~ i_25_)  &  (~ i_24_)  &  i_19_ ) ;
 assign wire124 = ( n_n1397  &  n_n1258  &  n_n1257  &  n_n1387 ) ;
 assign wire132 = ( n_n1397  &  n_n1257  &  n_n1384  &  n_n1251 ) ;
 assign wire550 = ( wire10  &  n_n1282 ) | ( wire290  &  n_n1254 ) ;
 assign wire8061 = ( wire133 ) | ( n_n1369  &  wire550  &  _11428 ) ;
 assign wire8062 = ( wire124 ) | ( wire132 ) | ( wire130 ) | ( wire134 ) ;
 assign n_n1583 = ( wire8061 ) | ( wire8062 ) | ( _31 ) | ( _32 ) ;
 assign n_n1582 = ( _11430 ) | ( _11431 ) ;
 assign wire557 = ( (~ i_9_)  &  i_7_  &  (~ i_14_) ) | ( (~ i_9_)  &  i_7_  &  (~ i_13_) ) ;
 assign wire555 = ( n_n1315  &  n_n1314 ) | ( n_n1322  &  wire557 ) ;
 assign wire8072 = ( wire111 ) | ( wire1651 ) | ( wire1652 ) ;
 assign n_n1584 = ( wire8072 ) | ( wire110 ) | ( _64 ) | ( _67 ) ;
 assign wire214 = ( (~ i_28_)  &  (~ i_34_)  &  i_35_  &  (~ i_29_) ) ;
 assign wire265 = ( (~ i_31_)  &  i_36_  &  (~ i_35_) ) ;
 assign wire267 = ( (~ i_27_)  &  (~ i_28_)  &  (~ i_23_)  &  (~ i_29_) ) ;
 assign wire559 = ( n_n1443  &  n_n1118  &  n_n1279 ) | ( n_n1408  &  n_n1118  &  n_n1279 ) ;
 assign wire6920 = ( (~ i_13_)  &  (~ i_23_)  &  (~ i_17_)  &  (~ i_16_) ) ;
 assign wire312 = ( n_n1443  &  n_n1118  &  n_n1279 ) ;
 assign wire6948 = ( (~ i_34_)  &  i_33_  &  i_35_ ) ;
 assign wire6949 = ( (~ i_28_)  &  i_25_  &  (~ i_29_) ) ;
 assign wire126 = ( n_n1438  &  wire6948  &  wire6949 ) ;
 assign wire7653 = ( i_14_  &  (~ i_28_)  &  (~ i_29_) ) ;
 assign wire128 = ( n_n1438  &  wire6948  &  wire7653 ) ;
 assign wire1649 = ( i_25_  &  (~ i_26_)  &  (~ i_24_)  &  (~ i_34_) ) ;
 assign wire1650 = ( i_25_  &  (~ i_23_)  &  (~ i_24_)  &  i_34_ ) ;
 assign wire452 = ( (~ i_26_)  &  (~ i_24_)  &  (~ i_34_) ) ;
 assign wire7761 = ( (~ i_7_)  &  (~ i_8_)  &  i_36_ ) ;
 assign wire363 = ( n_n1369  &  n_n1368  &  n_n1282  &  wire7761 ) ;
 assign wire420 = ( (~ i_14_)  &  i_13_  &  (~ i_17_)  &  (~ i_16_) ) ;
 assign wire7769 = ( (~ i_7_)  &  (~ i_32_)  &  i_36_ ) ;
 assign wire455 = ( wire232  &  wire44  &  wire7749  &  wire7769 ) ;
 assign wire956 = ( wire484  &  wire7765 ) | ( wire489  &  wire7765 ) ;
 assign wire958 = ( n_n1375  &  n_n1322  &  _9686  &  _11021 ) ;
 assign wire7776 = ( (~ i_14_)  &  i_13_  &  n_n825 ) ;
 assign wire7777 = ( n_n1406  &  n_n1213  &  n_n576 ) ;
 assign wire568 = ( n_n301  &  wire363 ) | ( wire7776  &  wire7777 ) ;
 assign n_n1511 = ( (~ i_28_)  &  i_31_  &  i_34_ ) ;
 assign n_n130 = ( (~ i_17_)  &  (~ i_16_)  &  (~ i_19_) ) ;
 assign wire475 = ( (~ i_6_)  &  (~ i_12_)  &  n_n1353  &  n_n1307 ) ;
 assign wire7050 = ( (~ i_6_)  &  (~ i_12_) ) ;
 assign n_n849 = ( n_n1353  &  n_n1307  &  _10708 ) ;
 assign n_n1059 = ( (~ i_34_)  &  (~ i_33_)  &  i_35_  &  i_38_ ) ;
 assign wire222 = ( (~ i_26_)  &  (~ i_23_)  &  (~ i_24_)  &  _9659 ) ;
 assign n_n18 = ( n_n1406  &  n_n1213  &  _9908 ) ;
 assign n_n21 = ( n_n1406  &  n_n1213  &  _9919 ) ;
 assign wire7942 = ( i_21_  &  i_31_  &  (~ i_34_)  &  i_35_ ) ;
 assign wire299 = ( (~ i_27_)  &  (~ i_28_)  &  (~ i_23_)  &  wire7942 ) ;
 assign wire6993 = ( (~ i_8_)  &  (~ i_14_)  &  (~ i_12_) ) ;
 assign wire342 = ( (~ i_8_)  &  (~ i_14_)  &  (~ i_12_)  &  _11215 ) ;
 assign wire7831 = ( (~ i_23_)  &  (~ i_24_)  &  (~ i_21_) ) ;
 assign wire478 = ( n_n1441  &  n_n1438  &  n_n880  &  wire7831 ) ;
 assign wire572 = ( wire43  &  n_n1315 ) | ( wire263  &  n_n1323 ) ;
 assign wire48 = ( (~ i_23_)  &  (~ i_24_)  &  (~ i_17_)  &  _9483 ) ;
 assign wire385 = ( i_36_  &  (~ i_35_)  &  n_n1459 ) ;
 assign wire7822 = ( (~ i_28_)  &  (~ i_23_)  &  (~ i_17_)  &  (~ i_21_) ) ;
 assign wire418 = ( wire79  &  wire7822 ) ;
 assign wire578 = ( i_3_  &  (~ i_18_) ) | ( (~ i_11_)  &  (~ i_19_) ) ;
 assign wire384 = ( n_n1375  &  n_n1400  &  n_n301 ) ;
 assign wire576 = ( wire367  &  wire221 ) | ( wire41  &  wire384 ) ;
 assign wire253 = ( (~ i_35_)  &  i_38_  &  n_n1439  &  n_n1340 ) ;
 assign wire330 = ( (~ i_24_)  &  (~ i_35_)  &  i_38_  &  wire71 ) ;
 assign wire405 = ( i_10_  &  i_12_ ) ;
 assign wire583 = ( n_n394 ) | ( n_n391 ) | ( n_n315 ) | ( n_n317 ) ;
 assign wire1281 = ( wire349  &  wire7454 ) | ( wire7259  &  wire7258  &  wire7454 ) ;
 assign wire1283 = ( wire71  &  wire12  &  wire423 ) | ( wire71  &  wire12  &  wire435 ) ;
 assign n_n1847 = ( wire1281 ) | ( wire1283 ) | ( wire253  &  wire583 ) ;
 assign wire585 = ( i_14_  &  i_13_ ) | ( i_12_  &  i_17_ ) ;
 assign wire7615 = ( wire1123 ) | ( _749 ) | ( _750 ) ;
 assign n_n1889 = ( wire7615 ) | ( _756 ) | ( _757 ) | ( _758 ) ;
 assign wire361 = ( (~ i_9_)  &  (~ i_6_)  &  (~ i_11_)  &  (~ i_19_) ) ;
 assign wire353 = ( (~ i_9_)  &  (~ i_5_)  &  (~ i_6_)  &  (~ i_18_) ) ;
 assign wire4 = ( n_n1307  &  wire361 ) | ( n_n787  &  wire353 ) ;
 assign wire7276 = ( (~ i_25_)  &  (~ i_24_)  &  (~ i_22_) ) ;
 assign wire56 = ( (~ i_35_)  &  i_38_  &  n_n1425  &  wire7276 ) ;
 assign wire226 = ( (~ i_31_)  &  (~ i_33_)  &  (~ i_35_)  &  i_38_ ) ;
 assign wire7272 = ( (~ i_7_)  &  (~ i_26_)  &  (~ i_24_)  &  (~ i_22_) ) ;
 assign wire1449 = ( (~ i_24_)  &  wire231  &  wire7275 ) | ( (~ i_24_)  &  wire521  &  wire7275 ) ;
 assign wire1450 = ( wire56  &  wire7281 ) | ( n_n1038  &  wire56  &  wire590 ) ;
 assign wire7282 = ( _390 ) | ( wire4  &  wire7269 ) ;
 assign n_n1856 = ( wire1449 ) | ( wire1450 ) | ( wire7282 ) ;
 assign wire81 = ( (~ i_35_)  &  i_38_  &  n_n1454 ) ;
 assign wire377 = ( (~ i_30_)  &  (~ i_28_)  &  n_n1197  &  n_n1523 ) ;
 assign wire1457 = ( i_38_  &  wire1461 ) | ( n_n416  &  _10849 ) ;
 assign wire7267 = ( wire1456 ) | ( n_n416  &  wire70 ) | ( wire70  &  n_n706 ) ;
 assign wire7290 = ( wire1437 ) | ( wire1439 ) | ( n_n706  &  wire7286 ) ;
 assign n_n1825 = ( n_n1856 ) | ( wire1457 ) | ( wire7267 ) | ( wire7290 ) ;
 assign wire1428 = ( i_10_  &  i_18_  &  n_n586  &  wire329 ) ;
 assign wire1429 = ( (~ i_24_)  &  wire231  &  wire7296 ) | ( (~ i_24_)  &  wire521  &  wire7296 ) ;
 assign wire1430 = ( (~ i_30_)  &  wire311  &  wire1435 ) | ( (~ i_30_)  &  wire311  &  wire1436 ) ;
 assign wire1431 = ( wire249  &  wire406 ) | ( n_n586  &  wire249  &  wire7271 ) ;
 assign n_n1854 = ( wire1428 ) | ( wire1429 ) | ( wire1430 ) | ( wire1431 ) ;
 assign wire1382 = ( n_n1466  &  wire223  &  n_n1419 ) | ( n_n1466  &  n_n1419  &  wire346 ) ;
 assign wire1383 = ( wire56  &  wire7344 ) | ( (~ i_13_)  &  wire56  &  wire37 ) ;
 assign wire1384 = ( n_n805  &  n_n1466  &  wire394 ) ;
 assign wire7345 = ( wire475  &  wire7340 ) | ( n_n300  &  wire7341 ) ;
 assign n_n1861 = ( wire1382 ) | ( wire1383 ) | ( wire1384 ) | ( wire7345 ) ;
 assign wire319 = ( (~ i_28_)  &  i_29_  &  n_n1369  &  n_n1274 ) ;
 assign wire6951 = ( (~ i_24_)  &  (~ i_34_) ) ;
 assign wire6952 = ( (~ i_23_)  &  (~ i_24_)  &  i_34_ ) ;
 assign wire599 = ( n_n1425  &  wire6951 ) | ( wire277  &  wire6952 ) ;
 assign wire6958 = ( (~ i_27_)  &  (~ i_28_)  &  (~ i_26_)  &  i_33_ ) ;
 assign wire598 = ( n_n1406  &  wire245 ) | ( n_n1396  &  wire6958 ) ;
 assign wire6957 = ( (~ i_7_)  &  (~ i_34_)  &  i_35_  &  i_37_ ) ;
 assign wire597 = ( i_21_  &  wire372 ) | ( n_n1302  &  wire6957 ) ;
 assign wire6961 = ( wire1710 ) | ( n_n1393  &  wire599  &  wire6953 ) ;
 assign wire6962 = ( wire1706 ) | ( n_n1438  &  wire597 ) ;
 assign wire6963 = ( wire1709 ) | ( n_n1429  &  wire598 ) ;
 assign n_n1718 = ( wire6961 ) | ( wire6962 ) | ( wire6963 ) ;
 assign wire317 = ( i_34_  &  i_37_  &  n_n1018  &  n_n1302 ) ;
 assign wire365 = ( (~ i_27_)  &  (~ i_28_)  &  (~ i_29_)  &  i_37_ ) ;
 assign wire601 = ( n_n358  &  wire221 ) | ( n_n355  &  wire48 ) ;
 assign wire273 = ( (~ i_28_)  &  i_34_  &  (~ i_29_)  &  _9459 ) ;
 assign wire256 = ( (~ i_32_)  &  i_34_  &  (~ i_29_)  &  _9456 ) ;
 assign wire600 = ( n_n195  &  wire273 ) | ( n_n437  &  wire256 ) ;
 assign wire6876 = ( (~ i_9_)  &  (~ i_7_)  &  (~ i_8_)  &  (~ i_6_) ) ;
 assign wire233 = ( n_n1406  &  n_n1213  &  n_n629  &  wire6876 ) ;
 assign wire246 = ( (~ i_34_)  &  (~ i_33_)  &  i_35_  &  i_37_ ) ;
 assign wire492 = ( i_35_  &  i_37_  &  n_n1375  &  n_n1311 ) ;
 assign wire63 = ( (~ i_20_)  &  (~ i_23_)  &  n_n460  &  n_n1369 ) ;
 assign wire268 = ( (~ i_14_)  &  (~ i_16_)  &  i_37_ ) ;
 assign wire431 = ( (~ i_11_)  &  (~ i_17_)  &  (~ i_16_)  &  (~ i_19_) ) ;
 assign wire6899 = ( (~ i_20_)  &  (~ i_23_)  &  (~ i_24_) ) ;
 assign wire508 = ( n_n1303  &  n_n245  &  wire44  &  wire6899 ) ;
 assign wire7053 = ( (~ i_30_)  &  (~ i_27_)  &  (~ i_28_) ) ;
 assign wire7976 = ( (~ i_21_)  &  i_36_ ) ;
 assign wire301 = ( n_n1141  &  n_n1213  &  wire7053  &  wire7976 ) ;
 assign wire7827 = ( i_10_  &  i_7_  &  i_13_ ) ;
 assign wire7828 = ( i_10_  &  i_7_  &  (~ i_12_) ) ;
 assign wire608 = ( n_n1408  &  wire7827 ) | ( n_n916  &  wire7828 ) ;
 assign wire360 = ( (~ i_8_)  &  (~ i_6_)  &  (~ i_12_)  &  _9999 ) ;
 assign wire437 = ( i_10_  &  i_7_  &  i_3_  &  (~ i_18_) ) ;
 assign wire891 = ( i_10_  &  i_7_  &  (~ i_11_)  &  (~ i_19_) ) ;
 assign wire610 = ( n_n1443  &  wire437 ) | ( n_n1429  &  wire437 ) | ( n_n1443  &  wire891 ) ;
 assign n_n1149 = ( (~ i_32_)  &  wire226 ) ;
 assign wire447 = ( (~ i_28_)  &  (~ i_24_)  &  i_34_  &  (~ i_29_) ) ;
 assign wire434 = ( n_n1307  &  n_n1033  &  _10498 ) ;
 assign wire7415 = ( (~ i_13_)  &  (~ i_4_)  &  (~ i_12_)  &  (~ i_2_) ) ;
 assign wire7466 = ( (~ i_30_)  &  (~ i_8_)  &  (~ i_28_)  &  (~ i_31_) ) ;
 assign wire235 = ( n_n1197  &  n_n1523  &  wire7466 ) ;
 assign wire1264 = ( wire1323  &  wire7465 ) | ( wire1324  &  wire7465 ) ;
 assign wire1265 = ( wire235  &  wire406 ) | ( n_n586  &  wire235  &  wire7271 ) ;
 assign wire1266 = ( wire288  &  wire12  &  wire434 ) | ( wire288  &  wire12  &  wire422 ) ;
 assign wire1267 = ( i_19_  &  wire288  &  n_n309  &  wire12 ) ;
 assign n_n1846 = ( wire1264 ) | ( wire1265 ) | ( wire1266 ) | ( wire1267 ) ;
 assign wire1111 = ( (~ i_28_)  &  i_31_  &  i_34_  &  (~ i_29_) ) ;
 assign wire616 = ( wire1111 ) | ( _746 ) | ( _747 ) ;
 assign wire615 = ( i_14_  &  i_13_ ) | ( i_12_  &  i_17_ ) ;
 assign wire614 = ( _744 ) | ( i_14_  &  i_13_  &  (~ i_24_) ) ;
 assign wire1105 = ( i_29_  &  wire61  &  wire615 ) ;
 assign wire1106 = ( i_21_  &  (~ i_22_)  &  wire372 ) ;
 assign n_n1892 = ( wire1105 ) | ( wire1106 ) | ( wire616  &  wire614 ) ;
 assign wire35 = ( i_30_  &  i_27_ ) | ( i_27_  &  i_32_ ) | ( i_16_  &  i_32_ ) ;
 assign wire7631 = ( wire35  &  wire7626 ) | ( n_n1519  &  wire7627 ) ;
 assign wire7632 = ( wire1095 ) | ( wire214  &  wire95 ) | ( wire214  &  wire96 ) ;
 assign n_n1837 = ( n_n1892 ) | ( wire7632 ) | ( _10232 ) ;
 assign wire7301 = ( (~ i_7_)  &  (~ i_32_)  &  i_38_ ) ;
 assign wire249 = ( n_n1425  &  wire7276  &  wire7301 ) ;
 assign wire311 = ( (~ i_28_)  &  (~ i_25_)  &  (~ i_26_)  &  i_38_ ) ;
 assign wire78 = ( (~ i_28_)  &  (~ i_25_)  &  (~ i_26_)  &  (~ i_22_) ) ;
 assign wire329 = ( (~ i_24_)  &  i_38_  &  wire77  &  wire78 ) ;
 assign wire344 = ( (~ i_28_)  &  (~ i_32_)  &  (~ i_33_)  &  (~ i_29_) ) ;
 assign wire1372 = ( wire1379  &  wire7352 ) | ( (~ i_22_)  &  wire343  &  wire7352 ) ;
 assign wire1377 = ( n_n1523  &  wire289  &  _10646 ) ;
 assign wire7357 = ( _490 ) | ( n_n819  &  wire7354  &  _10648 ) ;
 assign wire7358 = ( n_n706  &  wire456 ) | ( wire327  &  wire7355 ) ;
 assign wire218 = ( (~ i_9_)  &  (~ i_6_)  &  i_13_  &  _10782 ) ;
 assign wire7377 = ( (~ i_28_)  &  i_35_  &  i_38_  &  (~ i_29_) ) ;
 assign wire310 = ( n_n1307  &  n_n1100  &  n_n1311  &  wire7377 ) ;
 assign wire315 = ( i_34_  &  (~ i_35_)  &  i_38_  &  _10003 ) ;
 assign wire387 = ( (~ i_28_)  &  (~ i_33_)  &  (~ i_29_)  &  _10665 ) ;
 assign wire408 = ( (~ i_9_)  &  (~ i_8_)  &  (~ i_6_)  &  _10690 ) ;
 assign wire784 = ( wire1338 ) | ( wire425  &  wire7399 ) | ( wire454  &  wire7399 ) ;
 assign wire1337 = ( n_n1523  &  wire7266  &  wire346 ) ;
 assign wire7400 = ( _460 ) | ( wire61  &  wire261  &  _10142 ) ;
 assign wire271 = ( (~ i_28_)  &  (~ i_25_)  &  (~ i_29_)  &  _10480 ) ;
 assign wire278 = ( (~ i_30_)  &  (~ i_24_) ) ;
 assign wire346 = ( i_13_  &  (~ i_32_)  &  n_n1307  &  n_n1100 ) ;
 assign wire1330 = ( n_n1489  &  wire18  &  n_n1422  &  n_n998 ) ;
 assign wire320 = ( i_31_  &  i_34_  &  n_n1375 ) ;
 assign wire416 = ( (~ i_14_)  &  (~ i_35_)  &  i_37_ ) ;
 assign wire630 = ( n_n1406  &  wire245 ) | ( n_n1396  &  wire6958 ) ;
 assign wire629 = ( (~ i_14_)  &  (~ i_12_)  &  (~ i_16_) ) | ( (~ i_14_)  &  (~ i_17_)  &  (~ i_16_) ) ;
 assign wire1715 = ( wire302  &  n_n1489  &  wire452  &  wire416 ) ;
 assign wire1717 = ( n_n1390  &  n_n1372  &  n_n1334  &  n_n1375 ) ;
 assign wire6977 = ( wire1718 ) | ( wire1719 ) | ( n_n1443  &  wire630 ) ;
 assign n_n1719 = ( wire6977 ) | ( _9225 ) ;
 assign wire248 = ( i_34_  &  (~ i_35_)  &  i_37_ ) ;
 assign wire634 = ( (~ i_10_)  &  (~ i_14_)  &  (~ i_16_) ) | ( (~ i_14_)  &  i_13_  &  (~ i_16_) ) ;
 assign wire6937 = ( (~ i_27_)  &  (~ i_23_)  &  (~ i_24_)  &  _9514 ) ;
 assign wire6938 = ( (~ i_27_)  &  (~ i_28_)  &  (~ i_24_)  &  _9511 ) ;
 assign wire632 = ( wire312  &  wire6937 ) | ( n_n329  &  wire6938 ) ;
 assign wire88 = ( n_n245  &  wire44  &  wire6899 ) ;
 assign wire1565 = ( n_n1375  &  n_n1202  &  wire351 ) | ( n_n1375  &  n_n1202  &  wire1574 ) ;
 assign wire1566 = ( wire1576  &  wire7126 ) | ( wire1577  &  wire7126 ) ;
 assign wire1567 = ( _899 ) | ( n_n1274  &  n_n245  &  wire638 ) ;
 assign wire1697 = ( n_n1425  &  wire6979  &  _9227 ) ;
 assign wire1701 = ( n_n1433  &  wire54  &  n_n1489  &  wire416 ) ;
 assign wire6989 = ( wire1696 ) | ( wire1698 ) | ( wire1703 ) ;
 assign wire6990 = ( wire1699 ) | ( wire1700 ) | ( wire1702 ) | ( wire1704 ) ;
 assign n_n1720 = ( wire1697 ) | ( wire1701 ) | ( wire6989 ) | ( wire6990 ) ;
 assign wire1690 = ( n_n1406  &  n_n1213  &  _9325  &  _9328 ) ;
 assign wire7001 = ( wire1691 ) | ( _1105 ) | ( _1106 ) ;
 assign n_n1716 = ( wire7001 ) | ( _1108 ) | ( _1109 ) | ( _9338 ) ;
 assign wire1683 = ( n_n1406  &  n_n1213  &  _9325  &  _9347 ) ;
 assign wire7010 = ( _1102 ) | ( i_37_  &  wire8  &  wire306 ) ;
 assign wire7011 = ( wire1684 ) | ( _1098 ) | ( _1099 ) ;
 assign n_n1715 = ( wire7010 ) | ( wire7011 ) | ( _9361 ) ;
 assign wire1659 = ( n_n1441  &  n_n1400  &  wire7028 ) ;
 assign n_n1723 = ( wire1661 ) | ( wire1659 ) | ( _1084 ) ;
 assign wire7033 = ( (~ i_23_)  &  i_21_  &  (~ i_22_) ) ;
 assign wire7044 = ( n_n1718 ) | ( n_n1719 ) | ( n_n1720 ) | ( wire7043 ) ;
 assign wire7045 = ( n_n1716 ) | ( n_n1715 ) | ( n_n1723 ) | ( wire7022 ) ;
 assign wire440 = ( i_21_  &  (~ i_19_)  &  n_n712 ) ;
 assign wire644 = ( n_n1408  &  wire7827 ) | ( n_n916  &  wire7828 ) ;
 assign wire643 = ( n_n358  &  wire221 ) | ( n_n355  &  wire48 ) ;
 assign wire1086 = ( n_n1439  &  wire143 ) | ( n_n1439  &  wire1089 ) ;
 assign wire1087 = ( i_23_  &  wire1091 ) | ( i_23_  &  wire3  &  n_n1497 ) ;
 assign wire254 = ( (~ i_35_)  &  i_38_  &  n_n1305  &  n_n1497 ) ;
 assign wire381 = ( (~ i_35_)  &  i_38_  &  n_n1454  &  n_n1288 ) ;
 assign wire430 = ( (~ i_28_)  &  (~ i_26_)  &  (~ i_33_)  &  (~ i_29_) ) ;
 assign wire429 = ( (~ i_25_)  &  (~ i_34_)  &  i_35_  &  i_38_ ) ;
 assign wire1289 = ( (~ i_24_)  &  wire271  &  wire231 ) | ( (~ i_24_)  &  wire271  &  wire521 ) ;
 assign n_n1852 = ( wire1286 ) | ( _10478 ) | ( _10485 ) ;
 assign wire755 = ( n_n394 ) | ( n_n391 ) | ( n_n315 ) | ( n_n317 ) ;
 assign wire1314 = ( n_n294  &  wire253 ) | ( n_n371  &  wire253 ) | ( n_n284  &  wire253 ) ;
 assign wire1316 = ( wire288  &  wire12  &  wire423 ) | ( wire288  &  wire12  &  wire435 ) ;
 assign n_n1843 = ( wire1314 ) | ( wire1316 ) | ( n_n316  &  wire755 ) ;
 assign wire75 = ( (~ i_35_)  &  i_38_  &  n_n1423  &  wire7409 ) ;
 assign wire654 = ( n_n394 ) | ( n_n391 ) | ( n_n315 ) | ( n_n317 ) ;
 assign wire276 = ( (~ i_24_)  &  (~ i_35_)  &  i_38_  &  wire78 ) ;
 assign wire7427 = ( i_9_  &  (~ i_8_)  &  (~ i_13_)  &  i_11_ ) ;
 assign wire423 = ( n_n461  &  wire7411  &  wire7427 ) ;
 assign wire314 = ( n_n460  &  n_n1369  &  n_n1100 ) ;
 assign wire7136 = ( (~ i_14_)  &  (~ i_16_)  &  n_n1274 ) ;
 assign wire664 = ( (~ i_14_)  &  wire233 ) | ( wire314  &  wire7136 ) ;
 assign wire663 = ( (~ i_10_)  &  (~ i_14_)  &  (~ i_16_) ) | ( (~ i_14_)  &  i_13_  &  (~ i_16_) ) ;
 assign wire29 = ( (~ i_13_)  &  (~ i_12_)  &  (~ i_16_) ) | ( (~ i_13_)  &  (~ i_17_)  &  (~ i_16_) ) ;
 assign wire491 = ( n_n1307  &  n_n1314  &  n_n1144 ) ;
 assign wire7062 = ( wire1628 ) | ( _9584 ) | ( wire515  &  _9577 ) ;
 assign n_n1690 = ( wire7062 ) | ( wire7093 ) | ( _975 ) | ( _9636 ) ;
 assign wire668 = ( (~ i_14_)  &  (~ i_12_)  &  (~ i_16_) ) | ( (~ i_14_)  &  (~ i_17_)  &  (~ i_16_) ) ;
 assign wire383 = ( wire79  &  n_n460  &  n_n461  &  n_n1254 ) ;
 assign wire669 = ( n_n1408  &  wire7827 ) | ( n_n916  &  wire7828 ) ;
 assign wire390 = ( (~ i_33_)  &  (~ i_35_)  &  i_38_  &  wire61 ) ;
 assign wire435 = ( n_n1118  &  n_n1279  &  wire7428 ) ;
 assign wire1323 = ( n_n461  &  wire7411  &  n_n1028 ) ;
 assign wire1324 = ( n_n1118  &  n_n1279  &  n_n1048 ) ;
 assign wire1256 = ( wire1260  &  wire7469 ) | ( n_n735  &  wire405  &  wire7469 ) ;
 assign wire1257 = ( n_n307  &  wire7470 ) | ( n_n309  &  wire7470 ) ;
 assign wire1258 = ( wire12  &  wire434  &  wire7431 ) | ( wire12  &  wire422  &  wire7431 ) ;
 assign wire1259 = ( n_n1439  &  n_n1340  &  _10575  &  _10578 ) ;
 assign n_n1844 = ( wire1256 ) | ( wire1257 ) | ( wire1258 ) | ( wire1259 ) ;
 assign wire270 = ( (~ i_32_)  &  (~ i_35_)  &  i_38_  &  _10748 ) ;
 assign wire677 = ( n_n394 ) | ( n_n391 ) | ( n_n315 ) | ( n_n317 ) ;
 assign wire7477 = ( wire1247 ) | ( wire1249 ) | ( wire75  &  wire677 ) ;
 assign n_n1821 = ( n_n1846 ) | ( n_n1844 ) | ( wire7477 ) ;
 assign wire272 = ( n_n1307  &  n_n1288  &  n_n1100 ) ;
 assign wire379 = ( (~ i_34_)  &  i_35_  &  i_38_  &  _10889 ) ;
 assign wire482 = ( (~ i_35_)  &  i_37_  &  n_n1216  &  n_n1241 ) ;
 assign wire74 = ( (~ i_23_)  &  (~ i_24_)  &  (~ i_17_)  &  _11262 ) ;
 assign wire189 = ( i_14_  &  (~ i_28_)  &  n_n1438  &  wire6948 ) ;
 assign wire687 = ( (~ i_14_)  &  (~ i_12_)  &  (~ i_16_) ) | ( (~ i_14_)  &  (~ i_17_)  &  (~ i_16_) ) ;
 assign wire68 = ( i_9_  &  i_12_ ) ;
 assign wire692 = ( n_n1439  &  n_n1340 ) | ( n_n1423  &  wire7409 ) ;
 assign wire7502 = ( _624 ) | ( wire212  &  wire71 ) | ( wire212  &  wire430 ) ;
 assign wire7503 = ( wire1227 ) | ( n_n1306  &  wire692  &  _10038 ) ;
 assign wire7504 = ( wire124 ) | ( wire132 ) | ( _617 ) ;
 assign wire524 = ( (~ i_27_)  &  (~ i_28_)  &  (~ i_24_)  &  _9351 ) ;
 assign wire694 = ( (~ i_14_)  &  (~ i_12_)  &  (~ i_16_) ) | ( (~ i_14_)  &  (~ i_17_)  &  (~ i_16_) ) ;
 assign wire6960 = ( i_20_  &  (~ i_17_) ) ;
 assign wire7017 = ( i_20_  &  (~ i_16_) ) ;
 assign wire693 = ( n_n1401  &  wire6960 ) | ( n_n1391  &  wire7017 ) ;
 assign wire1587 = ( n_n504  &  wire57  &  wire1592 ) | ( n_n504  &  wire57  &  wire1593 ) ;
 assign wire7110 = ( wire1589 ) | ( n_n984  &  wire47  &  wire693 ) ;
 assign n_n1714 = ( wire1587 ) | ( wire7110 ) | ( wire1591 ) | ( _1027 ) ;
 assign wire470 = ( (~ i_33_)  &  i_37_  &  n_n1429 ) ;
 assign wire698 = ( wire367  &  wire221 ) | ( wire41  &  wire384 ) ;
 assign wire1542 = ( n_n1258  &  n_n1302  &  _9737  &  _9740 ) ;
 assign wire7169 = ( n_n458  &  wire7165 ) | ( wire384  &  wire7166 ) ;
 assign wire697 = ( wire1542 ) | ( wire7169 ) | ( n_n1437  &  wire698 ) ;
 assign n_n1703 = ( wire1534 ) | ( _9736 ) | ( i_37_  &  wire697 ) ;
 assign wire8010 = ( (~ i_27_)  &  (~ i_26_)  &  (~ i_2_)  &  (~ i_24_) ) ;
 assign wire295 = ( n_n1345  &  n_n576  &  n_n1282  &  wire8010 ) ;
 assign wire7523 = ( (~ i_24_)  &  i_34_  &  i_38_ ) ;
 assign wire286 = ( n_n1307  &  n_n1100  &  wire344  &  wire7523 ) ;
 assign wire1214 = ( n_n1279  &  n_n1202  &  _10169 ) ;
 assign wire7006 = ( (~ i_30_)  &  (~ i_32_)  &  i_31_ ) ;
 assign wire306 = ( n_n1375  &  n_n1213  &  wire7006 ) ;
 assign wire6984 = ( (~ i_30_)  &  (~ i_28_)  &  i_29_ ) ;
 assign wire7173 = ( (~ i_32_)  &  (~ i_29_)  &  n_n793 ) ;
 assign wire7174 = ( (~ i_28_)  &  (~ i_29_)  &  n_n1258 ) ;
 assign wire705 = ( n_n358  &  wire7173 ) | ( n_n355  &  wire7174 ) ;
 assign wire7177 = ( n_n1375  &  n_n1213  &  n_n1458 ) ;
 assign wire704 = ( n_n1404  &  wire508 ) | ( wire367  &  wire7177 ) ;
 assign wire1525 = ( _927 ) | ( _928 ) | ( _929 ) ;
 assign wire7183 = ( wire705  &  wire7175 ) | ( wire458  &  _9760 ) ;
 assign n_n1704 = ( wire1525 ) | ( wire7183 ) | ( i_37_  &  wire704 ) ;
 assign wire708 = ( n_n458  &  wire221 ) | ( n_n242  &  wire48 ) ;
 assign wire1511 = ( wire248  &  wire7191 ) | ( wire710  &  _9652 ) ;
 assign wire7188 = ( i_34_  &  (~ i_33_)  &  i_37_ ) ;
 assign wire712 = ( n_n363  &  wire273 ) | ( n_n620  &  wire256 ) ;
 assign wire289 = ( i_13_  &  (~ i_31_)  &  n_n1307  &  n_n841 ) ;
 assign wire327 = ( (~ i_6_)  &  (~ i_12_)  &  n_n1307  &  n_n1359 ) ;
 assign wire335 = ( i_9_  &  (~ i_5_)  &  (~ i_6_)  &  _10648 ) ;
 assign wire7356 = ( (~ i_28_)  &  i_38_  &  (~ i_29_) ) ;
 assign wire456 = ( (~ i_28_)  &  i_38_  &  (~ i_29_)  &  _10658 ) ;
 assign wire305 = ( (~ i_27_)  &  (~ i_28_)  &  (~ i_26_)  &  i_31_ ) ;
 assign wire717 = ( i_7_  &  (~ i_14_)  &  (~ i_12_) ) | ( i_7_  &  (~ i_13_)  &  (~ i_12_) ) ;
 assign wire716 = ( (~ i_14_)  &  (~ i_12_)  &  (~ i_16_) ) | ( (~ i_14_)  &  (~ i_17_)  &  (~ i_16_) ) ;
 assign wire6928 = ( (~ i_32_)  &  i_34_  &  (~ i_29_) ) ;
 assign wire1498 = ( n_n1278  &  wire404  &  wire7195 ) ;
 assign wire1499 = ( wire1507  &  wire7199 ) | ( wire1508  &  wire7199 ) ;
 assign wire1500 = ( wire365  &  wire1502 ) | ( wire261  &  wire365  &  _9847 ) ;
 assign wire1501 = ( i_37_  &  wire7205 ) | ( i_37_  &  wire272  &  _9857 ) ;
 assign n_n1701 = ( wire1498 ) | ( wire1499 ) | ( wire1500 ) | ( wire1501 ) ;
 assign wire1490 = ( wire1507  &  wire7212 ) | ( wire1508  &  wire7212 ) ;
 assign wire1493 = ( _881 ) | ( n_n1408  &  wire721  &  wire7218 ) ;
 assign wire7221 = ( wire272  &  _9876 ) | ( wire7210  &  _9880 ) ;
 assign wire274 = ( (~ i_20_)  &  (~ i_23_)  &  (~ i_24_)  &  wire44 ) ;
 assign wire7121 = ( (~ i_11_)  &  (~ i_23_)  &  (~ i_17_)  &  (~ i_19_) ) ;
 assign wire351 = ( n_n1307  &  n_n1100  &  wire268  &  wire7121 ) ;
 assign wire724 = ( n_n1408  &  wire7827 ) | ( n_n916  &  wire7828 ) ;
 assign wire7898 = ( (~ i_23_)  &  (~ i_24_)  &  (~ i_19_) ) ;
 assign wire8021 = ( i_3_  &  (~ i_18_) ) ;
 assign wire8022 = ( i_10_  &  i_7_  &  (~ i_23_)  &  (~ i_24_) ) ;
 assign wire723 = ( n_n712  &  wire7898 ) | ( wire8021  &  wire8022 ) ;
 assign wire394 = ( n_n1118  &  n_n1279  &  n_n1359 ) ;
 assign wire6996 = ( (~ i_27_)  &  (~ i_28_)  &  i_25_ ) ;
 assign wire6997 = ( i_20_  &  (~ i_23_)  &  (~ i_24_) ) ;
 assign wire322 = ( i_34_  &  i_33_  &  wire6996  &  wire6997 ) ;
 assign wire727 = ( (~ i_14_)  &  (~ i_12_)  &  (~ i_16_) ) | ( (~ i_14_)  &  (~ i_17_)  &  (~ i_16_) ) ;
 assign wire1581 = ( n_n1443  &  wire322 ) | ( n_n1443  &  wire1583 ) ;
 assign wire7116 = ( wire1580 ) | ( _1020 ) | ( _1021 ) ;
 assign wire7117 = ( wire1582 ) | ( wire1585  &  wire7114 ) | ( wire1586  &  wire7114 ) ;
 assign n_n1713 = ( wire1581 ) | ( wire7116 ) | ( wire7117 ) ;
 assign wire731 = ( n_n712  &  wire7898 ) | ( wire8021  &  wire8022 ) ;
 assign wire151 = ( wire47  &  wire7058  &  wire8042 ) ;
 assign wire345 = ( i_14_  &  (~ i_28_)  &  i_13_  &  i_22_ ) ;
 assign wire735 = ( i_30_ ) | ( i_32_ ) ;
 assign wire7686 = ( i_30_  &  i_12_  &  i_17_ ) | ( i_12_  &  i_17_  &  i_32_ ) ;
 assign wire734 = ( wire345  &  wire735 ) | ( wire83  &  wire7686 ) ;
 assign wire7547 = ( (~ i_28_)  &  (~ i_24_)  &  (~ i_33_)  &  (~ i_29_) ) ;
 assign wire502 = ( n_n1340  &  n_n1128  &  wire12 ) ;
 assign wire1190 = ( wire1197  &  wire7543 ) | ( n_n1028  &  wire7541  &  wire7543 ) ;
 assign wire1191 = ( (~ i_24_)  &  (~ i_29_)  &  wire261  &  wire311 ) ;
 assign wire7548 = ( wire51  &  wire502 ) | ( n_n1149  &  wire7545 ) ;
 assign wire7549 = ( _834 ) | ( _835 ) ;
 assign n_n1875 = ( wire1190 ) | ( wire1191 ) | ( wire7548 ) | ( wire7549 ) ;
 assign wire1202 = ( wire425  &  wire7534 ) | ( wire454  &  wire7534 ) ;
 assign wire1203 = ( wire223  &  n_n1302  &  _10151 ) ;
 assign wire7537 = ( wire1201 ) | ( n_n1423  &  n_n805  &  wire7531 ) ;
 assign wire7538 = ( (~ i_10_)  &  wire286 ) | ( wire257  &  wire7536 ) ;
 assign n_n1873 = ( wire1202 ) | ( wire1203 ) | ( wire7537 ) | ( wire7538 ) ;
 assign wire7570 = ( wire7567 ) | ( _816 ) | ( _817 ) | ( _10051 ) ;
 assign n_n1831 = ( n_n1875 ) | ( wire7570 ) | ( _10053 ) ;
 assign wire7598 = ( n_n1873 ) | ( wire7529 ) | ( _10186 ) ;
 assign wire740 = ( i_20_ ) | ( i_21_ ) ;
 assign wire7639 = ( (~ i_24_)  &  (~ i_22_)  &  i_34_ ) ;
 assign wire739 = ( n_n1523  &  (~ n_n1251) ) | ( wire740  &  wire7639 ) ;
 assign wire7622 = ( wire1132 ) | ( wire1135 ) | ( wire7609 ) | ( wire7621 ) ;
 assign wire7642 = ( _10282 ) | ( _10283 ) ;
 assign n_n1818 = ( n_n1889 ) | ( n_n1837 ) | ( wire7622 ) | ( wire7642 ) ;
 assign wire1043 = ( wire249  &  _10319 ) | ( _678  &  _10319 ) | ( _679  &  _10319 ) ;
 assign wire7680 = ( wire1029 ) | ( wire7676 ) | ( wire7678 ) | ( _668 ) ;
 assign n_n1834 = ( wire7680 ) | ( _10331 ) | ( _10332 ) | ( _10353 ) ;
 assign n_n1887 = ( wire7699 ) | ( _657 ) | ( _658 ) ;
 assign wire7705 = ( wire1000 ) | ( wire214  &  wire1008 ) | ( wire214  &  wire1009 ) ;
 assign n_n1835 = ( n_n1887 ) | ( wire7689 ) | ( _10408 ) | ( _10409 ) ;
 assign wire744 = ( wire262 ) | ( wire436 ) | ( i_19_  &  wire18 ) ;
 assign wire745 = ( (~ i_14_)  &  (~ i_12_)  &  (~ i_16_) ) | ( (~ i_14_)  &  (~ i_17_)  &  (~ i_16_) ) ;
 assign wire1053 = ( _686 ) | ( n_n1353  &  wire7547  &  _10288 ) ;
 assign wire1054 = ( _683 ) | ( _684 ) | ( _685 ) ;
 assign wire7661 = ( wire1050 ) | ( wire1051 ) | ( wire1052 ) ;
 assign wire457 = ( (~ i_28_)  &  (~ i_26_)  &  (~ i_24_)  &  (~ i_29_) ) ;
 assign wire465 = ( n_n1433  &  n_n1466  &  wire12 ) ;
 assign wire510 = ( (~ i_32_)  &  (~ i_35_)  &  i_38_  &  wire71 ) ;
 assign wire1474 = ( (~ i_33_)  &  wire1480 ) | ( (~ i_33_)  &  wire524  &  wire758 ) ;
 assign wire7244 = ( wire1476 ) | ( wire59  &  n_n1429  &  wire306 ) ;
 assign n_n1712 = ( wire1474 ) | ( wire7244 ) | ( _1015 ) | ( _1016 ) ;
 assign wire515 = ( n_n1307  &  n_n1144  &  n_n1263 ) ;
 assign wire1634 = ( n_n1216  &  n_n620  &  wire6928 ) ;
 assign wire771 = ( (~ i_14_)  &  (~ i_12_)  &  (~ i_16_) ) | ( (~ i_14_)  &  (~ i_17_)  &  (~ i_16_) ) ;
 assign wire7588 = ( wire395  &  wire7585 ) | ( wire81  &  wire7586 ) ;
 assign wire7591 = ( wire1156 ) | ( wire1157 ) | ( _803 ) ;
 assign wire425 = ( (~ i_13_)  &  wire1342 ) | ( (~ i_13_)  &  wire1343 ) ;
 assign wire454 = ( i_19_  &  wire1340 ) | ( i_19_  &  wire1341 ) ;
 assign wire1338 = ( wire262  &  wire239  &  n_n1422 ) | ( wire436  &  wire239  &  n_n1422 ) ;
 assign wire7399 = ( (~ i_24_)  &  i_38_  &  n_n1437 ) ;
 assign wire1069 = ( n_n1278  &  n_n1279  &  n_n1523  &  wire7266 ) ;
 assign wire792 = ( (~ i_13_)  &  (~ i_12_)  &  (~ i_16_) ) | ( (~ i_13_)  &  (~ i_17_)  &  (~ i_16_) ) ;
 assign wire7699 = ( wire1010 ) | ( wire1011 ) | ( wire1012 ) | ( wire1014 ) ;
 assign wire7145 = ( (~ i_9_)  &  (~ i_6_)  &  (~ i_23_)  &  (~ i_24_) ) ;
 assign wire484 = ( (~ i_11_)  &  (~ i_19_)  &  n_n1307  &  wire7145 ) ;
 assign wire7148 = ( (~ i_5_)  &  (~ i_6_)  &  (~ i_23_)  &  (~ i_24_) ) ;
 assign wire489 = ( (~ i_9_)  &  (~ i_18_)  &  n_n787  &  wire7148 ) ;
 assign wire7428 = ( i_9_  &  (~ i_13_)  &  i_11_  &  i_18_ ) ;
 assign wire422 = ( n_n1118  &  n_n1058  &  wire7415 ) ;
 assign wire349 = ( (~ i_13_)  &  i_11_  &  i_18_  &  (~ i_22_) ) ;
 assign wire413 = ( (~ i_8_)  &  (~ i_18_)  &  (~ i_17_)  &  (~ i_16_) ) ;
 assign wire7342 = ( i_11_  &  i_18_ ) ;
 assign wire7343 = ( (~ i_2_)  &  i_19_ ) ;
 assign wire37 = ( n_n1192  &  wire7342 ) | ( n_n1038  &  wire7343 ) ;
 assign wire211 = ( (~ i_7_)  &  (~ i_32_) ) ;
 assign wire65 = ( (~ i_7_)  &  (~ i_32_)  &  n_n1213  &  wire7053 ) ;
 assign wire1663 = ( (~ i_24_)  &  (~ i_34_)  &  n_n1425  &  wire7026 ) ;
 assign wire802 = ( (~ i_13_)  &  (~ i_12_)  &  (~ i_16_) ) | ( (~ i_13_)  &  (~ i_17_)  &  (~ i_16_) ) ;
 assign wire95 = ( i_30_  &  i_23_ ) | ( i_27_  &  i_32_ ) | ( i_23_  &  i_32_ ) ;
 assign wire96 = ( i_30_  &  i_27_ ) | ( i_30_  &  i_16_ ) | ( i_16_  &  i_32_ ) ;
 assign wire143 = ( i_30_  &  i_16_  &  i_34_ ) ;
 assign wire7178 = ( n_n1375  &  n_n1400  &  n_n916 ) ;
 assign wire458 = ( (~ i_23_)  &  (~ i_24_)  &  (~ i_17_)  &  _9495 ) ;
 assign wire7274 = ( (~ i_8_)  &  (~ i_5_)  &  (~ i_6_)  &  (~ i_18_) ) ;
 assign wire231 = ( wire404  &  wire7274 ) ;
 assign wire7055 = ( (~ i_20_)  &  (~ i_23_)  &  (~ i_24_) ) ;
 assign wire251 = ( n_n1441  &  wire77  &  wire7055 ) ;
 assign wire334 = ( (~ i_10_)  &  (~ i_14_)  &  (~ i_16_) ) ;
 assign wire343 = ( i_9_  &  (~ i_3_)  &  (~ i_13_)  &  i_11_ ) ;
 assign wire7890 = ( (~ i_7_)  &  (~ i_8_)  &  (~ i_12_)  &  (~ i_21_) ) ;
 assign wire356 = ( n_n1406  &  n_n461  &  n_n1213  &  wire7890 ) ;
 assign wire402 = ( (~ i_20_)  &  (~ i_13_)  &  (~ i_12_)  &  (~ i_16_) ) ;
 assign wire1432 = ( (~ i_13_)  &  i_12_  &  i_18_  &  i_19_ ) ;
 assign wire1433 = ( (~ i_13_)  &  i_12_  &  i_11_  &  i_18_ ) ;
 assign wire1434 = ( (~ i_3_)  &  (~ i_13_)  &  i_12_  &  i_19_ ) ;
 assign wire406 = ( i_10_  &  wire1432 ) | ( i_10_  &  wire1433 ) | ( i_10_  &  wire1434 ) ;
 assign wire1342 = ( i_9_  &  (~ i_8_)  &  i_11_  &  i_18_ ) ;
 assign wire1343 = ( i_9_  &  (~ i_8_)  &  (~ i_3_)  &  i_11_ ) ;
 assign wire7576 = ( (~ i_28_)  &  (~ i_26_)  &  (~ i_24_)  &  (~ i_29_) ) ;
 assign wire438 = ( (~ i_32_)  &  wire226  &  wire7576 ) ;
 assign wire1340 = ( i_9_  &  (~ i_8_)  &  (~ i_13_)  &  i_18_ ) ;
 assign wire1341 = ( i_9_  &  (~ i_8_)  &  (~ i_3_)  &  (~ i_13_) ) ;
 assign wire498 = ( n_n787  &  n_n1118  &  n_n180  &  n_n179 ) ;
 assign wire517 = ( n_n1375  &  wire13  &  n_n1322  &  n_n820 ) ;
 assign wire521 = ( (~ i_11_)  &  (~ i_19_)  &  n_n1307  &  n_n841 ) ;
 assign wire522 = ( n_n1307  &  n_n841  &  n_n177  &  n_n178 ) ;
 assign wire7254 = ( n_n1278  &  n_n26  &  wire413 ) ;
 assign wire526 = ( wire431  &  wire508 ) | ( wire274  &  wire7254 ) ;
 assign wire544 = ( n_n1443  &  wire437 ) | ( n_n1429  &  wire437 ) | ( n_n1429  &  wire891 ) ;
 assign wire7259 = ( (~ i_3_)  &  i_19_ ) | ( i_18_  &  i_19_ ) ;
 assign wire582 = ( wire349 ) | ( (~ i_13_)  &  (~ i_22_)  &  wire7259 ) ;
 assign wire590 = ( (~ i_13_)  &  i_12_  &  i_11_ ) | ( (~ i_13_)  &  i_12_  &  i_19_ ) ;
 assign wire593 = ( (~ i_13_)  &  i_12_  &  i_11_ ) | ( (~ i_13_)  &  i_12_  &  i_19_ ) ;
 assign wire604 = ( n_n245  &  wire361 ) | ( n_n26  &  wire353 ) ;
 assign wire6892 = ( i_3_  &  (~ i_4_)  &  (~ i_0_)  &  wire6891 ) ;
 assign wire6894 = ( (~ i_5_)  &  (~ i_4_)  &  (~ i_0_)  &  _9929 ) ;
 assign wire603 = ( n_n21  &  wire6892 ) | ( n_n18  &  wire6894 ) ;
 assign wire6913 = ( (~ i_32_)  &  (~ i_33_)  &  i_37_ ) ;
 assign wire606 = ( n_n504  &  n_n1118 ) | ( n_n1278  &  wire6913 ) ;
 assign wire624 = ( n_n1307  &  wire361 ) | ( n_n787  &  wire353 ) ;
 assign wire635 = ( (~ i_9_)  &  (~ i_10_)  &  (~ i_6_) ) | ( (~ i_9_)  &  (~ i_6_)  &  i_13_ ) ;
 assign wire1570 = ( n_n460  &  n_n1369  &  n_n1100  &  wire7130 ) ;
 assign wire1572 = ( n_n1369  &  n_n1368  &  n_n841  &  n_n504 ) ;
 assign wire1573 = ( wire59  &  n_n460  &  n_n1369  &  n_n1100 ) ;
 assign wire638 = ( wire1570 ) | ( n_n301  &  wire1572 ) | ( n_n301  &  wire1573 ) ;
 assign wire657 = ( n_n307 ) | ( n_n309 ) | ( wire1323 ) | ( wire1324 ) ;
 assign wire661 = ( i_7_  &  (~ i_14_)  &  (~ i_12_) ) | ( i_7_  &  (~ i_13_)  &  (~ i_12_) ) ;
 assign wire666 = ( wire43  &  n_n1274 ) | ( (~ i_23_)  &  wire402 ) ;
 assign wire7473 = ( (~ i_3_)  &  (~ i_22_) ) ;
 assign wire679 = ( i_12_  &  wire349 ) | ( n_n586  &  wire7473 ) ;
 assign wire1604 = ( (~ i_20_)  &  (~ i_13_)  &  (~ i_17_)  &  (~ i_16_) ) ;
 assign wire683 = ( wire402 ) | ( wire1604 ) ;
 assign wire710 = ( n_n1307  &  n_n853  &  n_n1408 ) | ( n_n1307  &  n_n1408  &  n_n839 ) ;
 assign wire713 = ( n_n712  &  wire7898 ) | ( wire8021  &  wire8022 ) ;
 assign wire7217 = ( (~ i_32_)  &  i_37_ ) ;
 assign wire721 = ( n_n1318  &  n_n1118 ) | ( n_n1278  &  wire7217 ) ;
 assign wire741 = ( i_30_ ) | ( i_32_ ) | ( i_31_ ) ;
 assign wire759 = ( (~ i_13_)  &  (~ i_12_)  &  (~ i_16_) ) | ( (~ i_13_)  &  (~ i_17_)  &  (~ i_16_) ) ;
 assign wire758 = ( n_n1314  &  n_n1141 ) | ( n_n1322  &  wire7243 ) ;
 assign wire767 = ( (~ i_13_)  &  i_12_  &  i_11_ ) | ( (~ i_13_)  &  i_12_  &  i_19_ ) ;
 assign wire1766 = ( n_n1278  &  wire404  &  n_n132  &  wire6882 ) ;
 assign wire22 = ( wire1766  &  wire6923  &  _11531 ) | ( wire6923  &  _11531  &  _11532 ) ;
 assign wire1767 = ( n_n1307  &  n_n1100  &  n_n177  &  n_n178 ) ;
 assign wire1768 = ( n_n1278  &  n_n787  &  n_n180  &  n_n179 ) ;
 assign wire34 = ( wire227  &  n_n1375  &  wire1767 ) | ( wire227  &  n_n1375  &  wire1768 ) ;
 assign wire105 = ( wire232  &  n_n178  &  wire8086 ) ;
 assign wire107 = ( n_n180  &  n_n1303  &  wire338 ) ;
 assign wire8090 = ( (~ i_17_)  &  i_36_  &  n_n1406  &  n_n1213 ) ;
 assign wire8091 = ( (~ i_9_)  &  (~ i_7_)  &  (~ i_6_)  &  (~ i_23_) ) ;
 assign wire8086 = ( (~ i_7_)  &  (~ i_8_)  &  (~ i_19_) ) ;
 assign wire6947 = ( (~ i_27_)  &  (~ i_23_)  &  i_22_  &  i_35_ ) ;
 assign wire110 = ( n_n1429  &  n_n1326  &  wire6947 ) | ( n_n1408  &  n_n1326  &  wire6947 ) ;
 assign wire111 = ( n_n1396  &  n_n1404  &  n_n1374  &  n_n1375 ) ;
 assign wire117 = ( n_n1438  &  wire6948  &  _11425 ) ;
 assign wire8056 = ( i_25_  &  (~ i_32_)  &  (~ i_31_)  &  i_33_ ) ;
 assign wire8057 = ( (~ i_28_)  &  i_31_ ) ;
 assign wire130 = ( n_n1369  &  n_n1315  &  n_n1263  &  wire8057 ) ;
 assign wire133 = ( n_n1443  &  n_n1406  &  n_n1213  &  wire7491 ) ;
 assign wire134 = ( n_n1404  &  n_n1326  &  wire6947 ) ;
 assign wire142 = ( wire10  &  n_n793  &  n_n1315  &  wire7942 ) ;
 assign wire150 = ( n_n1397  &  n_n1092  &  n_n1406  &  n_n1408 ) ;
 assign wire7058 = ( (~ i_27_)  &  (~ i_28_)  &  i_33_ ) ;
 assign wire8042 = ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  (~ i_16_) ) ;
 assign wire8043 = ( (~ i_16_)  &  i_31_  &  (~ i_34_)  &  i_35_ ) ;
 assign wire158 = ( n_n1375  &  n_n1141  &  n_n1263  &  n_n820 ) ;
 assign wire160 = ( wire227  &  n_n1489  &  n_n1089  &  n_n1251 ) ;
 assign wire161 = ( n_n1429  &  n_n1397  &  n_n1092  &  n_n1406 ) ;
 assign wire163 = ( wire245  &  n_n984  &  n_n916  &  wire7828 ) ;
 assign wire169 = ( i_3_  &  (~ i_18_)  &  n_n1429  &  wire8022 ) ;
 assign wire164 = ( wire320  &  wire169 ) | ( n_n1443  &  wire320  &  wire713 ) ;
 assign wire8008 = ( (~ i_2_)  &  (~ i_17_)  &  (~ i_21_)  &  (~ i_16_) ) ;
 assign wire166 = ( wire7053  &  wire8008  &  _9404  &  _11202 ) ;
 assign wire172 = ( n_n1408  &  wire245  &  n_n984  &  wire7827 ) ;
 assign wire8007 = ( n_n263  &  wire273 ) | ( n_n269  &  wire256 ) ;
 assign wire178 = ( n_n1404  &  n_n1397  &  n_n1092  &  n_n1406 ) ;
 assign wire7802 = ( (~ i_27_)  &  (~ i_23_)  &  (~ i_24_)  &  i_21_ ) ;
 assign wire183 = ( wire10  &  n_n1315  &  n_n1511  &  wire7802 ) ;
 assign wire184 = ( n_n1504  &  n_n1375  &  n_n1322  &  n_n1323 ) ;
 assign wire7803 = ( i_34_  &  i_29_ ) ;
 assign wire185 = ( n_n1216  &  n_n1092  &  wire687  &  wire7803 ) ;
 assign wire187 = ( n_n1504  &  n_n1315  &  n_n1314  &  n_n1375 ) ;
 assign wire7997 = ( (~ i_27_)  &  (~ i_23_)  &  (~ i_24_)  &  (~ i_17_) ) ;
 assign wire7999 = ( (~ i_23_)  &  i_34_  &  i_33_ ) ;
 assign wire7984 = ( i_25_  &  i_21_ ) ;
 assign wire192 = ( wire47  &  wire668  &  wire7058  &  wire7984 ) ;
 assign wire194 = ( n_n1504  &  n_n1375  &  n_n1322  &  n_n1285 ) ;
 assign wire200 = ( n_n1441  &  n_n1390  &  wire7105 ) ;
 assign wire201 = ( n_n1441  &  n_n1400  &  wire258 ) ;
 assign wire197 = ( wire79  &  n_n1089  &  n_n1431  &  n_n1254 ) ;
 assign wire198 = ( n_n1504  &  n_n1315  &  n_n1375  &  n_n1263 ) ;
 assign wire7105 = ( (~ i_8_)  &  (~ i_13_)  &  (~ i_12_) ) ;
 assign wire7971 = ( (~ i_23_)  &  (~ i_17_)  &  i_21_ ) ;
 assign wire234 = ( n_n1216  &  n_n1374  &  n_n1387  &  wire7971 ) ;
 assign wire304 = ( wire79  &  n_n1147  &  n_n1431  &  n_n1254 ) ;
 assign wire7787 = ( (~ i_30_)  &  (~ i_32_)  &  i_34_  &  i_36_ ) ;
 assign wire336 = ( n_n1390  &  n_n1375  &  n_n1089  &  wire7787 ) ;
 assign wire339 = ( n_n1425  &  wire340  &  _11141 ) ;
 assign wire7784 = ( (~ i_30_)  &  i_34_  &  i_36_  &  (~ i_29_) ) ;
 assign wire350 = ( n_n1216  &  n_n1141  &  n_n1263  &  wire7784 ) ;
 assign wire7961 = ( (~ i_2_)  &  i_36_  &  n_n825 ) ;
 assign wire417 = ( wire227  &  n_n1489  &  n_n1147  &  n_n1251 ) ;
 assign wire7949 = ( (~ i_30_)  &  (~ i_7_)  &  (~ i_28_)  &  (~ i_29_) ) ;
 assign wire424 = ( wire227  &  wire43  &  n_n1258  &  wire7949 ) ;
 assign wire7940 = ( (~ i_30_)  &  (~ i_31_) ) ;
 assign wire427 = ( n_n1390  &  wire86  &  wire7105  &  wire7940 ) ;
 assign wire439 = ( n_n1314  &  n_n1141  &  n_n820 ) ;
 assign wire7945 = ( (~ i_2_)  &  i_36_  &  n_n825 ) ;
 assign wire469 = ( wire227  &  wire10  &  n_n1258  &  wire7949 ) ;
 assign wire471 = ( n_n1443  &  n_n1397  &  n_n1092  &  n_n1406 ) ;
 assign wire7930 = ( (~ i_32_)  &  (~ i_34_)  &  i_36_  &  (~ i_35_) ) ;
 assign wire494 = ( n_n1497  &  n_n1459  &  wire7930 ) ;
 assign wire6982 = ( (~ i_28_)  &  (~ i_23_)  &  (~ i_24_) ) ;
 assign wire7931 = ( (~ i_32_)  &  i_34_  &  i_36_  &  (~ i_35_) ) ;
 assign wire497 = ( n_n1459  &  wire6982  &  wire7931 ) ;
 assign wire507 = ( n_n1396  &  wire546  &  wire6958 ) ;
 assign wire7025 = ( (~ i_23_)  &  (~ i_24_)  &  i_22_  &  i_34_ ) ;
 assign wire512 = ( n_n1406  &  wire8  &  wire7025 ) ;
 assign wire813 = ( n_n1489  &  wire340  &  wire452 ) ;
 assign wire7900 = ( (~ i_9_)  &  i_2_ ) ;
 assign wire825 = ( wire44  &  wire7749  &  wire420  &  wire7900 ) ;
 assign wire829 = ( n_n1369  &  n_n1128  &  wire515 ) ;
 assign wire7901 = ( (~ i_10_)  &  (~ i_13_)  &  (~ i_17_)  &  (~ i_16_) ) ;
 assign wire833 = ( wire44  &  wire7749  &  wire7900  &  wire7901 ) ;
 assign wire7903 = ( n_n242  &  wire458 ) | ( n_n458  &  wire7902 ) ;
 assign wire834 = ( i_36_  &  wire7903 ) | ( wire356  &  _11360 ) ;
 assign wire7887 = ( n_n1263  &  wire80  &  wire86 ) ;
 assign wire7892 = ( n_n355  &  wire458 ) | ( n_n458  &  wire7889 ) ;
 assign wire843 = ( i_36_  &  wire7892 ) | ( wire356  &  _11362 ) ;
 assign wire849 = ( n_n1322  &  wire80  &  _11087  &  _11089 ) ;
 assign wire857 = ( i_21_  &  (~ i_19_)  &  n_n1443  &  n_n712 ) ;
 assign wire850 = ( wire275  &  wire857 ) | ( i_21_  &  wire275  &  wire544 ) ;
 assign wire7868 = ( (~ i_32_)  &  i_34_  &  n_n1307  &  n_n1100 ) ;
 assign wire7871 = ( n_n458  &  wire7869 ) | ( n_n242  &  wire7870 ) ;
 assign wire7819 = ( (~ i_28_)  &  i_29_  &  n_n1369  &  n_n1254 ) ;
 assign wire881 = ( wire232  &  n_n1406  &  n_n1213  &  wire7860 ) ;
 assign wire7858 = ( _278 ) | ( _279 ) ;
 assign wire7859 = ( (~ i_5_)  &  (~ i_6_)  &  n_n1279  &  wire7857 ) ;
 assign wire7862 = ( (~ i_17_)  &  (~ i_21_)  &  (~ i_16_)  &  _11063 ) ;
 assign wire875 = ( wire881  &  wire7862 ) | ( wire7858  &  wire7859  &  wire7862 ) ;
 assign wire7860 = ( (~ i_10_)  &  (~ i_13_) ) ;
 assign wire7820 = ( (~ i_13_)  &  (~ i_31_)  &  i_36_  &  (~ i_35_) ) ;
 assign wire910 = ( n_n1307  &  n_n1408  &  n_n576  &  n_n839 ) ;
 assign wire911 = ( n_n1443  &  n_n1118  &  n_n1279  &  wire265 ) ;
 assign wire906 = ( n_n1375  &  n_n1213  &  wire910 ) | ( n_n1375  &  n_n1213  &  wire911 ) ;
 assign wire7791 = ( (~ i_27_)  &  (~ i_28_)  &  (~ i_26_)  &  i_36_ ) ;
 assign wire919 = ( n_n1390  &  n_n1472  &  n_n1147  &  wire7791 ) ;
 assign wire7798 = ( i_20_  &  (~ i_26_)  &  (~ i_24_)  &  (~ i_21_) ) ;
 assign wire924 = ( n_n1438  &  n_n1326  &  wire7798 ) ;
 assign wire925 = ( n_n1216  &  wire13  &  wire260  &  wire7784 ) ;
 assign wire926 = ( (~ i_30_)  &  (~ i_28_)  &  wire245  &  wire340 ) ;
 assign wire928 = ( n_n1216  &  n_n1092  &  wire533  &  wire7803 ) ;
 assign wire7782 = ( (~ i_28_)  &  (~ i_24_)  &  i_34_  &  i_29_ ) ;
 assign wire933 = ( n_n1438  &  n_n1092  &  wire7782 ) ;
 assign wire937 = ( n_n1390  &  n_n1375  &  n_n1147  &  wire7787 ) ;
 assign wire939 = ( n_n1390  &  n_n1472  &  n_n1089  &  wire7791 ) ;
 assign wire942 = ( wire420  &  wire7772  &  _11519 ) | ( wire950  &  wire7772  &  _11519 ) ;
 assign wire943 = ( n_n1369  &  wire498  &  _11521 ) | ( n_n1369  &  wire522  &  _11521 ) ;
 assign wire948 = ( n_n576  &  wire484  &  wire7778 ) | ( n_n576  &  wire489  &  wire7778 ) ;
 assign wire945 = ( n_n1443  &  wire948 ) | ( wire455  &  _11510 ) ;
 assign wire7778 = ( (~ i_27_)  &  (~ i_28_)  &  (~ i_26_)  &  (~ i_29_) ) ;
 assign wire950 = ( (~ i_10_)  &  (~ i_13_)  &  (~ i_17_)  &  (~ i_16_) ) ;
 assign wire953 = ( wire80  &  wire86  &  wire498 ) | ( wire80  &  wire86  &  wire522 ) ;
 assign wire7765 = ( n_n1443  &  n_n1375  &  n_n1422 ) ;
 assign wire7766 = ( n_n1216  &  n_n1278  &  wire6928 ) ;
 assign wire7751 = ( wire431  &  wire7750 ) | ( wire969  &  wire7750 ) ;
 assign wire7757 = ( n_n1216  &  n_n1307  &  n_n1100  &  wire6928 ) ;
 assign wire969 = ( i_3_  &  (~ i_18_)  &  (~ i_17_)  &  (~ i_16_) ) ;
 assign wire981 = ( n_n1486  &  n_n1118  &  n_n1279  &  n_n1359 ) ;
 assign wire7736 = ( (~ i_26_)  &  (~ i_24_)  &  n_n1288 ) ;
 assign wire977 = ( n_n1197  &  wire981 ) | ( n_n1197  &  wire335  &  wire7736 ) ;
 assign wire978 = ( (~ i_10_)  &  (~ i_31_)  &  n_n1307  &  n_n841 ) ;
 assign wire988 = ( wire349  &  wire7723 ) | ( wire7259  &  wire7258  &  wire7723 ) ;
 assign wire7258 = ( (~ i_13_)  &  (~ i_22_) ) ;
 assign wire7723 = ( i_9_  &  (~ i_28_)  &  (~ i_26_)  &  (~ i_24_) ) ;
 assign wire1406 = ( (~ i_11_)  &  (~ i_19_)  &  n_n1307  &  n_n1100 ) ;
 assign wire7716 = ( (~ i_28_)  &  (~ i_26_)  &  (~ i_29_)  &  _10705 ) ;
 assign wire994 = ( n_n1307  &  n_n1359  &  wire7050  &  wire7717 ) ;
 assign wire996 = ( (~ i_9_)  &  (~ i_6_)  &  i_13_  &  _10717 ) ;
 assign wire7718 = ( n_n841  &  _10715 ) | ( n_n841  &  _10716 ) ;
 assign wire7717 = ( (~ i_28_)  &  (~ i_25_)  &  (~ i_32_)  &  (~ i_29_) ) ;
 assign wire7701 = ( (~ i_30_)  &  (~ i_7_)  &  (~ i_2_)  &  (~ i_32_) ) ;
 assign wire999 = ( (~ i_33_)  &  i_38_  &  wire61  &  wire7701 ) ;
 assign wire7702 = ( (~ i_32_)  &  (~ i_33_)  &  (~ i_35_)  &  i_38_ ) ;
 assign wire1000 = ( n_n1497  &  n_n1459  &  wire7702 ) ;
 assign wire7704 = ( (~ i_8_)  &  (~ i_26_)  &  (~ i_24_) ) ;
 assign wire1008 = ( i_30_  &  i_12_  &  i_17_ ) | ( i_12_  &  i_17_  &  i_32_ ) ;
 assign wire1009 = ( i_30_  &  i_14_  &  i_13_ ) | ( i_14_  &  i_13_  &  i_32_ ) ;
 assign wire7308 = ( (~ i_28_)  &  (~ i_24_)  &  i_38_ ) ;
 assign wire7690 = ( (~ i_30_)  &  (~ i_8_)  &  (~ i_31_)  &  (~ i_29_) ) ;
 assign wire1010 = ( n_n1437  &  wire7308  &  wire7690 ) ;
 assign wire7691 = ( (~ i_30_)  &  (~ i_7_)  &  (~ i_8_)  &  (~ i_2_) ) ;
 assign wire1011 = ( n_n1523  &  wire7266  &  wire7691 ) ;
 assign wire1015 = ( (~ i_28_)  &  i_12_  &  i_17_  &  i_22_ ) ;
 assign wire1012 = ( n_n1504  &  wire345 ) | ( n_n1504  &  wire1015 ) ;
 assign wire1014 = ( (~ i_7_)  &  (~ i_32_)  &  n_n1489  &  n_n1059 ) ;
 assign wire1017 = ( n_n1423  &  n_n1422  &  n_n1459 ) ;
 assign wire1022 = ( (~ i_7_)  &  (~ i_28_)  &  n_n1472  &  wire429 ) ;
 assign wire1023 = ( n_n1489  &  n_n805  &  _10386 ) ;
 assign wire1024 = ( n_n1489  &  wire13  &  n_n1059 ) | ( n_n1489  &  wire13  &  wire429 ) ;
 assign wire7670 = ( (~ i_30_)  &  (~ i_8_)  &  (~ i_2_) ) ;
 assign wire1029 = ( wire61  &  wire226  &  wire7670 ) ;
 assign wire1030 = ( n_n1353  &  n_n1197  &  n_n1497  &  wire57 ) ;
 assign wire1032 = ( (~ wire3)  &  n_n1197  &  n_n1486  &  n_n1359 ) ;
 assign wire1033 = ( n_n1369  &  n_n1368  &  wire7033  &  wire792 ) ;
 assign wire1041 = ( n_n1353  &  n_n1423  &  n_n805  &  wire57 ) ;
 assign wire1044 = ( n_n1307  &  n_n1303  &  wire430  &  _10324 ) ;
 assign wire1045 = ( n_n1303  &  wire71  &  _10034  &  _10326 ) ;
 assign wire7655 = ( (~ i_8_)  &  (~ i_2_)  &  (~ i_22_) ) ;
 assign wire1050 = ( n_n1454  &  n_n1361  &  n_n1345  &  wire7655 ) ;
 assign wire7657 = ( (~ i_30_)  &  (~ i_2_)  &  (~ i_32_)  &  (~ i_31_) ) ;
 assign wire1051 = ( wire12  &  wire78  &  wire7657 ) ;
 assign wire1052 = ( n_n1369  &  n_n1368  &  wire7033  &  wire745 ) ;
 assign wire7644 = ( i_9_  &  (~ i_10_)  &  (~ i_2_) ) ;
 assign wire1060 = ( n_n1425  &  n_n1179  &  wire7276  &  wire7644 ) ;
 assign wire7647 = ( (~ i_28_)  &  (~ i_25_)  &  i_34_  &  (~ i_29_) ) ;
 assign wire1062 = ( n_n1278  &  n_n1279  &  wire7492  &  wire7647 ) ;
 assign wire1064 = ( (~ i_32_)  &  wire1069 ) | ( (~ i_32_)  &  _614 ) | ( (~ i_32_)  &  _615 ) ;
 assign wire1077 = ( i_12_  &  (~ i_24_)  &  i_17_  &  i_31_ ) ;
 assign wire7638 = ( i_14_  &  i_13_  &  (~ i_24_) ) ;
 assign wire1070 = ( wire58  &  wire1077 ) | ( wire58  &  wire741  &  wire7638 ) ;
 assign wire1082 = ( i_27_  &  i_31_ ) | ( i_23_  &  i_31_ ) | ( i_16_  &  i_31_ ) ;
 assign wire7636 = ( i_30_  &  i_16_ ) | ( i_14_  &  i_33_ ) ;
 assign wire1080 = ( n_n1497  &  wire35 ) | ( n_n1497  &  wire1082 ) | ( n_n1497  &  wire7636 ) ;
 assign wire1081 = ( i_23_  &  wire447 ) ;
 assign wire1089 = ( i_27_  &  i_31_  &  i_34_ ) | ( i_16_  &  i_31_  &  i_34_ ) ;
 assign wire1091 = ( (~ i_28_)  &  (~ i_24_)  &  i_22_  &  i_34_ ) ;
 assign wire1095 = ( (~ i_28_)  &  (~ i_29_)  &  n_n1504  &  (~ n_n1251) ) ;
 assign wire1100 = ( (~ i_28_)  &  i_22_  &  wire143 ) | ( (~ i_28_)  &  i_22_  &  wire1101 ) ;
 assign wire1101 = ( i_14_  &  i_34_  &  i_33_ ) ;
 assign wire7616 = ( (~ i_24_)  &  i_34_  &  (~ i_33_)  &  i_38_ ) ;
 assign wire1112 = ( (~ i_7_)  &  (~ i_28_)  &  n_n1472  &  wire7616 ) ;
 assign wire7618 = ( (~ i_28_)  &  i_22_  &  (~ i_34_)  &  i_35_ ) ;
 assign wire1113 = ( wire95  &  wire7618 ) | ( wire96  &  wire7618 ) ;
 assign wire1121 = ( i_14_  &  i_13_  &  (~ i_24_) ) ;
 assign wire7619 = ( (~ i_28_)  &  i_22_  &  i_31_  &  i_34_ ) ;
 assign wire1114 = ( n_n1519  &  wire7619 ) | ( wire1121  &  wire7619 ) ;
 assign wire1123 = ( (~ i_28_)  &  (~ i_29_)  &  n_n1504  &  wire585 ) ;
 assign wire7612 = ( i_30_  &  (~ i_28_)  &  i_22_ ) | ( (~ i_28_)  &  i_22_  &  i_32_ ) ;
 assign wire7600 = ( (~ i_7_)  &  (~ i_8_)  &  (~ i_24_)  &  i_38_ ) ;
 assign wire1131 = ( (~ i_30_)  &  (~ i_29_)  &  n_n1478  &  wire7600 ) ;
 assign wire7602 = ( (~ i_30_)  &  (~ i_7_)  &  (~ i_32_) ) ;
 assign wire1132 = ( (~ i_24_)  &  i_38_  &  wire71  &  wire7602 ) ;
 assign wire7603 = ( (~ i_30_)  &  (~ i_7_)  &  (~ i_8_)  &  (~ i_24_) ) ;
 assign wire1133 = ( (~ i_33_)  &  i_38_  &  n_n1486  &  wire7603 ) ;
 assign wire1134 = ( i_20_  &  (~ i_22_)  &  wire372 ) ;
 assign wire1137 = ( i_14_  &  (~ i_34_)  &  i_33_  &  i_35_ ) ;
 assign wire1135 = ( wire83  &  wire1137 ) | ( n_n1504  &  wire83  &  (~ n_n1251) ) ;
 assign wire1136 = ( (~ i_7_)  &  (~ i_32_)  &  n_n1489  &  wire503 ) ;
 assign wire1147 = ( (~ i_35_)  &  i_38_  &  n_n1454  &  n_n1128 ) ;
 assign wire1139 = ( _791 ) | ( n_n1307  &  n_n1144  &  wire1147 ) ;
 assign wire1140 = ( _788 ) | ( _789 ) ;
 assign wire1150 = ( n_n1478  &  n_n1133  &  wire12 ) ;
 assign wire1141 = ( n_n1307  &  wire7050  &  wire438 ) | ( n_n1307  &  wire7050  &  wire1150 ) ;
 assign wire1142 = ( n_n1278  &  n_n1279  &  wire7492  &  wire78 ) ;
 assign wire1143 = ( n_n1406  &  n_n1213  &  wire7491  &  wire8 ) ;
 assign wire7582 = ( (~ i_30_)  &  i_12_ ) ;
 assign wire1152 = ( n_n1353  &  wire12  &  wire78  &  wire7582 ) ;
 assign wire1156 = ( (~ i_24_)  &  wire223  &  wire380 ) | ( (~ i_24_)  &  wire380  &  wire261 ) ;
 assign wire1157 = ( n_n1307  &  wire7050  &  wire502 ) | ( n_n1307  &  wire7050  &  wire465 ) ;
 assign wire7572 = ( i_9_  &  (~ i_10_)  &  (~ i_8_)  &  i_12_ ) ;
 assign wire1159 = ( n_n1425  &  n_n1197  &  wire205  &  wire7572 ) ;
 assign wire1161 = ( n_n1118  &  n_n1279  &  wire226  &  wire457 ) ;
 assign wire1164 = ( n_n1478  &  n_n1133  &  wire12 ) ;
 assign wire1162 = ( wire224  &  n_n1279  &  wire438 ) | ( wire224  &  n_n1279  &  wire1164 ) ;
 assign wire1168 = ( n_n1425  &  wire7276  &  _10085 ) ;
 assign wire7559 = ( (~ i_30_)  &  (~ i_32_)  &  (~ i_35_)  &  i_38_ ) ;
 assign wire1173 = ( n_n1179  &  wire262  &  wire71  &  wire278 ) ;
 assign wire1176 = ( n_n1278  &  n_n1279  &  n_n1288  &  n_n1059 ) ;
 assign wire1197 = ( (~ i_13_)  &  wire1342 ) | ( (~ i_13_)  &  wire1343 ) | ( (~ i_13_)  &  wire1198 ) ;
 assign wire7541 = ( i_18_  &  i_19_ ) ;
 assign wire7543 = ( (~ i_30_)  &  (~ i_24_)  &  n_n1197  &  n_n1486 ) ;
 assign wire1198 = ( i_9_  &  (~ i_8_)  &  (~ i_3_)  &  i_19_ ) ;
 assign wire7532 = ( (~ i_8_)  &  (~ i_28_)  &  (~ i_29_) ) ;
 assign wire1201 = ( n_n1278  &  n_n1279  &  n_n1059  &  wire7532 ) ;
 assign wire7534 = ( (~ i_30_)  &  (~ i_29_)  &  n_n1478  &  wire12 ) ;
 assign wire1211 = ( wire1214  &  _10173 ) | ( _767  &  _10173 ) ;
 assign wire1227 = ( wire77  &  wire78  &  _10432 ) ;
 assign wire7488 = ( i_9_  &  (~ i_10_)  &  (~ i_2_) ) ;
 assign wire1230 = ( n_n1197  &  n_n1523  &  n_n1431  &  wire7488 ) ;
 assign wire1234 = ( n_n1406  &  n_n1213  &  wire7491  &  wire539 ) ;
 assign wire1235 = ( n_n1278  &  n_n1279  &  wire7492  &  wire288 ) ;
 assign wire7479 = ( (~ i_28_)  &  (~ i_22_)  &  n_n1454  &  wire264 ) ;
 assign wire1238 = ( wire521  &  wire7479 ) | ( wire404  &  wire7274  &  wire7479 ) ;
 assign wire1240 = ( n_n1466  &  n_n416  &  n_n1419 ) | ( n_n1466  &  n_n1419  &  n_n706 ) ;
 assign wire1242 = ( n_n394  &  wire254 ) | ( n_n391  &  wire254 ) ;
 assign wire1253 = ( (~ i_3_)  &  i_19_  &  _10586 ) | ( i_18_  &  i_19_  &  _10586 ) ;
 assign wire7474 = ( n_n1454  &  n_n1179  &  n_n1345 ) ;
 assign wire1247 = ( wire1253  &  wire7474 ) | ( i_10_  &  wire679  &  wire7474 ) ;
 assign wire1249 = ( i_19_  &  n_n307  &  wire288  &  wire12 ) ;
 assign wire1260 = ( i_10_  &  wire1263 ) | ( i_10_  &  (~ i_3_)  &  wire767 ) ;
 assign wire7469 = ( n_n1425  &  wire7276  &  _10560 ) ;
 assign wire7470 = ( (~ i_35_)  &  i_38_  &  n_n1225  &  n_n998 ) ;
 assign wire7431 = ( (~ i_28_)  &  (~ i_25_)  &  i_34_  &  (~ i_29_) ) ;
 assign wire1263 = ( (~ i_13_)  &  i_12_  &  i_11_  &  i_18_ ) ;
 assign wire7465 = ( (~ i_35_)  &  i_38_  &  n_n1486  &  n_n998 ) ;
 assign wire7271 = ( i_10_  &  (~ i_3_) ) ;
 assign wire7459 = ( (~ i_35_)  &  i_38_  &  n_n1486  &  n_n998 ) ;
 assign wire1268 = ( n_n307  &  wire7459 ) | ( n_n309  &  wire7459 ) ;
 assign wire1271 = ( wire71  &  wire12  &  wire434 ) | ( wire71  &  wire12  &  wire422 ) ;
 assign wire7456 = ( (~ i_24_)  &  (~ i_35_)  &  i_38_  &  wire430 ) ;
 assign wire1274 = ( _10626 ) | ( wire7456  &  _530 ) | ( wire7456  &  _531 ) ;
 assign wire7454 = ( n_n1438  &  n_n1197  &  n_n1497  &  wire405 ) ;
 assign wire7446 = ( wire61  &  wire226 ) ;
 assign wire1286 = ( n_n416  &  n_n1419  &  n_n1302 ) | ( n_n1419  &  n_n1302  &  n_n706 ) ;
 assign wire1291 = ( n_n394  &  wire381 ) | ( n_n391  &  wire381 ) | ( n_n317  &  wire381 ) ;
 assign wire1303 = ( wire435  &  _10823 ) | ( _406  &  _10823 ) | ( _407  &  _10823 ) ;
 assign wire1305 = ( wire12  &  wire78  &  wire423 ) | ( wire12  &  wire78  &  wire435 ) ;
 assign wire7430 = ( (~ i_35_)  &  i_38_  &  n_n1225  &  n_n998 ) ;
 assign wire1308 = ( wire1323  &  wire7430 ) | ( wire1324  &  wire7430 ) ;
 assign wire1309 = ( wire12  &  wire423  &  wire7431 ) | ( wire12  &  wire435  &  wire7431 ) ;
 assign wire1317 = ( n_n372  &  wire75 ) | ( n_n294  &  wire75 ) | ( n_n371  &  wire75 ) ;
 assign wire1319 = ( n_n338  &  wire1323 ) | ( n_n338  &  wire1324 ) ;
 assign wire7402 = ( (~ i_30_)  &  (~ i_24_)  &  n_n805  &  n_n1466 ) ;
 assign wire1325 = ( wire425  &  wire7402 ) | ( wire454  &  wire7402 ) ;
 assign wire1347 = ( _451 ) | ( n_n1197  &  n_n1486  &  n_n849 ) ;
 assign wire7388 = ( (~ i_10_)  &  (~ i_26_)  &  (~ i_24_) ) | ( i_13_  &  (~ i_26_)  &  (~ i_24_) ) ;
 assign wire1349 = ( n_n1307  &  n_n841  &  n_n1128  &  wire7388 ) ;
 assign wire7390 = ( (~ i_28_)  &  (~ i_26_)  &  (~ i_32_)  &  (~ i_29_) ) ;
 assign wire1350 = ( n_n1307  &  n_n1359  &  wire7050  &  wire7390 ) ;
 assign wire1351 = ( n_n1307  &  n_n853  &  n_n1133  &  n_n1497 ) ;
 assign wire7375 = ( wire283  &  wire343 ) | ( i_9_  &  wire283  &  n_n735 ) ;
 assign wire1356 = ( wire377  &  wire7375 ) | ( (~ i_13_)  &  wire377  &  wire37 ) ;
 assign wire1357 = ( wire223  &  n_n1419  &  n_n1302 ) ;
 assign wire7364 = ( (~ i_32_)  &  (~ i_29_)  &  wire311 ) ;
 assign wire1367 = ( (~ i_24_)  &  wire297  &  wire7364 ) | ( (~ i_24_)  &  wire1406  &  wire7364 ) ;
 assign wire1379 = ( i_9_  &  wire349 ) | ( i_9_  &  wire7259  &  wire7258 ) ;
 assign wire7352 = ( (~ i_35_)  &  i_38_  &  n_n1454  &  wire7351 ) ;
 assign wire7344 = ( wire283  &  wire343 ) | ( i_9_  &  wire283  &  n_n735 ) ;
 assign wire7332 = ( i_34_  &  (~ i_33_)  &  i_38_ ) ;
 assign wire1392 = ( _363 ) | ( n_n1439  &  n_n416  &  wire7332 ) ;
 assign wire7317 = ( i_34_  &  i_38_  &  (~ i_29_) ) ;
 assign wire1399 = ( n_n1423  &  n_n416  &  wire7317 ) | ( n_n1423  &  n_n706  &  wire7317 ) ;
 assign wire1404 = ( (~ i_24_)  &  wire297  &  wire7324 ) | ( (~ i_24_)  &  wire1406  &  wire7324 ) ;
 assign wire1405 = ( _322 ) | ( n_n1300  &  wire61  &  wire1426 ) ;
 assign wire1403 = ( (~ i_32_)  &  wire1404 ) | ( (~ i_32_)  &  wire1405 ) ;
 assign wire7324 = ( i_34_  &  i_38_  &  n_n1466 ) ;
 assign wire1426 = ( (~ i_11_)  &  (~ i_19_)  &  n_n1307  &  n_n1100 ) ;
 assign wire1412 = ( n_n1425  &  wire1414 ) | ( n_n1425  &  wire1435 ) | ( n_n1425  &  wire1436 ) ;
 assign wire1408 = ( _343 ) | ( (~ i_33_)  &  i_38_  &  wire1412 ) ;
 assign wire1414 = ( wire205  &  wire1416  &  wire7297 ) | ( wire205  &  wire1417  &  wire7297 ) ;
 assign wire1435 = ( (~ i_24_)  &  (~ i_22_)  &  wire7297  &  wire7298 ) ;
 assign wire1436 = ( i_10_  &  (~ i_3_)  &  n_n586  &  wire7299 ) ;
 assign wire1416 = ( (~ i_13_)  &  i_12_  &  i_18_  &  i_19_ ) ;
 assign wire1417 = ( (~ i_13_)  &  i_12_  &  i_11_  &  i_18_ ) ;
 assign wire7297 = ( i_10_  &  (~ i_7_)  &  (~ i_8_) ) ;
 assign wire1419 = ( _342 ) | ( n_n1419  &  wire344  &  wire1426 ) ;
 assign wire7311 = ( i_34_  &  (~ i_33_)  &  (~ i_35_)  &  i_38_ ) ;
 assign wire7296 = ( (~ i_31_)  &  (~ i_35_)  &  i_38_  &  wire7295 ) ;
 assign wire7298 = ( (~ i_3_)  &  (~ i_13_)  &  i_12_  &  i_19_ ) ;
 assign wire7299 = ( (~ i_7_)  &  (~ i_8_)  &  (~ i_24_)  &  (~ i_22_) ) ;
 assign wire1443 = ( wire68  &  wire349 ) | ( wire68  &  wire7259  &  wire7258 ) ;
 assign wire7284 = ( i_12_  &  (~ i_22_) ) ;
 assign wire7285 = ( (~ i_35_)  &  i_38_  &  n_n1454  &  n_n1431 ) ;
 assign wire1437 = ( wire1443  &  wire7285 ) | ( wire262  &  wire7284  &  wire7285 ) ;
 assign wire7288 = ( n_n584  &  n_n1033 ) | ( n_n735  &  wire7277 ) ;
 assign wire1439 = ( wire377  &  wire7288 ) | ( n_n1038  &  wire377  &  wire593 ) ;
 assign wire7275 = ( (~ i_28_)  &  (~ i_26_)  &  (~ i_29_)  &  wire226 ) ;
 assign wire7281 = ( n_n584  &  n_n1033 ) | ( n_n735  &  wire7277 ) ;
 assign wire1460 = ( i_12_  &  wire61  &  wire262 ) ;
 assign wire7261 = ( i_9_  &  i_12_  &  n_n1497 ) ;
 assign wire1456 = ( n_n762  &  wire1460 ) | ( n_n762  &  wire582  &  wire7261 ) ;
 assign wire1461 = ( n_n1454  &  wire1463  &  wire7264 ) | ( n_n1454  &  wire1464  &  wire7264 ) ;
 assign wire1463 = ( (~ i_18_)  &  (~ i_32_)  &  n_n1278  &  wire404 ) ;
 assign wire1464 = ( n_n1307  &  n_n1100  &  _10850 ) ;
 assign wire7264 = ( (~ i_28_)  &  (~ i_22_) ) ;
 assign wire6906 = ( (~ i_9_)  &  (~ i_7_)  &  (~ i_6_)  &  (~ i_32_) ) ;
 assign wire1480 = ( n_n1489  &  n_n1018  &  wire759  &  wire7108 ) ;
 assign wire6998 = ( (~ i_27_)  &  i_25_ ) ;
 assign wire1476 = ( n_n1257  &  wire47  &  wire29  &  wire6998 ) ;
 assign wire7108 = ( (~ i_32_)  &  i_31_  &  i_34_  &  i_37_ ) ;
 assign wire7224 = ( n_n1443  &  n_n504  &  n_n1118  &  n_n152 ) ;
 assign wire7214 = ( n_n1406  &  n_n1213  &  n_n629 ) ;
 assign wire7228 = ( n_n1443  &  n_n1441  &  n_n1318  &  n_n1305 ) ;
 assign wire1483 = ( wire484  &  wire7228 ) | ( wire489  &  wire7228 ) ;
 assign wire7229 = ( (~ i_35_)  &  i_37_  &  n_n1369  &  n_n1302 ) ;
 assign wire1484 = ( wire498  &  wire7229 ) | ( wire522  &  wire7229 ) ;
 assign wire1576 = ( n_n1303  &  wire431  &  _9821 ) ;
 assign wire1577 = ( n_n1278  &  wire404  &  wire413 ) ;
 assign wire7230 = ( (~ i_14_)  &  i_37_  &  n_n1018  &  n_n1225 ) ;
 assign wire1507 = ( wire404  &  n_n1118  &  n_n179 ) ;
 assign wire1508 = ( n_n1307  &  n_n841  &  wire7197 ) ;
 assign wire7212 = ( (~ i_35_)  &  i_37_  &  n_n1369  &  wire7211 ) ;
 assign wire7215 = ( (~ i_14_)  &  (~ i_32_)  &  (~ i_35_)  &  i_37_ ) ;
 assign wire7216 = ( (~ i_10_)  &  (~ i_14_)  &  (~ i_16_)  &  i_37_ ) ;
 assign wire7218 = ( n_n152  &  wire44  &  wire6899 ) ;
 assign wire7219 = ( (~ i_27_)  &  (~ i_28_)  &  (~ i_26_)  &  _9872 ) ;
 assign wire7195 = ( n_n1216  &  n_n179  &  wire268  &  wire6928 ) ;
 assign wire7199 = ( (~ i_14_)  &  (~ i_16_)  &  wire80  &  wire248 ) ;
 assign wire1502 = ( n_n1408  &  n_n1422  &  wire484 ) | ( n_n1408  &  n_n1422  &  wire489 ) ;
 assign wire7205 = ( wire319  &  wire7203 ) | ( wire223  &  wire7204 ) ;
 assign wire7197 = ( (~ i_11_)  &  (~ i_23_)  &  (~ i_17_)  &  (~ i_19_) ) ;
 assign wire1514 = ( n_n460  &  n_n1369  &  wire6885  &  wire7186 ) ;
 assign wire7185 = ( (~ i_14_)  &  (~ i_16_)  &  n_n1144 ) ;
 assign wire7187 = ( (~ i_35_)  &  i_37_  &  n_n245 ) ;
 assign wire1509 = ( wire1514  &  wire7187 ) | ( wire222  &  wire7185  &  wire7187 ) ;
 assign wire7191 = ( n_n1307  &  n_n841  &  wire7189 ) | ( n_n1307  &  n_n841  &  wire7190 ) ;
 assign wire6885 = ( (~ i_20_)  &  (~ i_23_) ) ;
 assign wire7186 = ( (~ i_6_)  &  (~ i_14_)  &  (~ i_12_)  &  (~ i_16_) ) ;
 assign wire1539 = ( n_n460  &  n_n1369  &  wire6885  &  wire7159 ) ;
 assign wire7158 = ( (~ i_13_)  &  (~ i_16_)  &  n_n1144 ) ;
 assign wire7160 = ( (~ i_33_)  &  (~ i_35_)  &  i_37_  &  _9724 ) ;
 assign wire1534 = ( wire1539  &  wire7160 ) | ( wire222  &  wire7158  &  wire7160 ) ;
 assign wire7161 = ( (~ i_5_)  &  (~ i_4_)  &  (~ i_0_)  &  (~ i_32_) ) ;
 assign wire7163 = ( (~ i_13_)  &  (~ i_16_)  &  (~ i_33_)  &  i_37_ ) ;
 assign wire7159 = ( (~ i_6_)  &  (~ i_13_)  &  (~ i_12_)  &  (~ i_16_) ) ;
 assign wire7151 = ( n_n1443  &  n_n1375  &  n_n1318  &  n_n1340 ) ;
 assign wire1546 = ( wire484  &  wire7151 ) | ( wire489  &  wire7151 ) ;
 assign wire1548 = ( wire482  &  wire498 ) | ( wire482  &  wire522 ) ;
 assign wire1550 = ( n_n1278  &  n_n152  &  wire1553 ) | ( n_n1278  &  n_n152  &  wire1554 ) ;
 assign wire1551 = ( n_n1375  &  n_n1322  &  _9686  &  _9688 ) ;
 assign wire1552 = ( n_n1307  &  n_n1288  &  n_n1100  &  _9683 ) ;
 assign wire1549 = ( wire59  &  wire1550 ) | ( wire59  &  wire1551 ) | ( wire59  &  wire1552 ) ;
 assign wire1553 = ( wire44  &  wire6899  &  wire7153 ) ;
 assign wire1554 = ( n_n1369  &  n_n1274  &  n_n1368  &  wire259 ) ;
 assign wire7153 = ( (~ i_13_)  &  (~ i_17_)  &  (~ i_16_)  &  (~ i_32_) ) ;
 assign wire1561 = ( n_n1278  &  wire404  &  n_n132  &  wire6882 ) ;
 assign wire1559 = ( wire317  &  wire1561 ) | ( wire317  &  _9784 ) ;
 assign wire6882 = ( (~ i_8_)  &  (~ i_13_) ) ;
 assign wire7120 = ( n_n1443  &  n_n504  &  wire7119 ) ;
 assign wire1574 = ( n_n1278  &  wire404  &  n_n179  &  wire7123 ) ;
 assign wire7126 = ( (~ i_14_)  &  i_37_  &  n_n793  &  wire6923 ) ;
 assign wire7130 = ( (~ i_14_)  &  i_13_  &  (~ i_16_)  &  i_37_ ) ;
 assign wire7123 = ( (~ i_14_)  &  (~ i_16_)  &  i_37_ ) ;
 assign wire7059 = ( i_20_  &  i_25_ ) ;
 assign wire1580 = ( wire47  &  wire727  &  wire7058  &  wire7059 ) ;
 assign wire1583 = ( wire59  &  n_n1375  &  n_n1213  &  wire7006 ) ;
 assign wire1582 = ( n_n1429  &  n_n1374  &  wire6996  &  wire6997 ) ;
 assign wire1585 = ( n_n1390  &  n_n1375  &  wire7105 ) ;
 assign wire1586 = ( n_n1375  &  n_n1400  &  wire259 ) ;
 assign wire1592 = ( n_n1441  &  n_n1390  &  wire7105 ) ;
 assign wire1593 = ( n_n1441  &  n_n1400  &  wire259 ) ;
 assign wire7009 = ( (~ i_28_)  &  (~ i_34_)  &  i_35_  &  i_29_ ) ;
 assign wire1589 = ( n_n1080  &  wire694  &  wire7009 ) ;
 assign wire1591 = ( n_n1489  &  n_n1018  &  wire8  &  wire7108 ) ;
 assign wire1600 = ( wire59  &  wire1603 ) | ( wire59  &  wire65  &  wire683 ) ;
 assign wire7099 = ( _1070 ) | ( n_n1429  &  wire251  &  _9409 ) ;
 assign wire1597 = ( (~ i_0_)  &  wire1600 ) | ( (~ i_0_)  &  wire7099 ) ;
 assign wire1603 = ( n_n1443  &  n_n1441  &  wire77  &  wire7055 ) ;
 assign wire7080 = ( (~ i_30_)  &  (~ i_27_)  &  (~ i_28_)  &  (~ i_29_) ) ;
 assign wire1607 = ( n_n1314  &  n_n1141  &  wire246  &  wire7080 ) ;
 assign wire7084 = ( (~ i_0_)  &  (~ i_33_)  &  (~ i_35_)  &  i_37_ ) ;
 assign wire1608 = ( _983 ) | ( wire666  &  _9616 ) ;
 assign wire1611 = ( n_n1225  &  n_n363  &  _9621 ) ;
 assign wire7083 = ( (~ i_20_)  &  (~ i_13_)  &  (~ i_17_)  &  (~ i_16_) ) ;
 assign wire7063 = ( (~ i_30_)  &  i_31_  &  (~ i_29_) ) ;
 assign wire7064 = ( (~ i_32_)  &  (~ i_34_)  &  i_35_  &  i_37_ ) ;
 assign wire1618 = ( n_n793  &  wire771  &  wire7063  &  wire7064 ) ;
 assign wire1623 = ( wire10  &  n_n1369  &  n_n1274  &  n_n1431 ) ;
 assign wire1625 = ( wire7053  &  wire7070  &  _9587 ) ;
 assign wire7072 = ( (~ i_0_)  &  (~ i_35_)  &  i_37_ ) ;
 assign wire1622 = ( n_n1443  &  wire47  &  wire7058  &  wire7059 ) ;
 assign wire7068 = ( (~ i_27_)  &  (~ i_26_)  &  (~ i_23_)  &  (~ i_24_) ) ;
 assign wire7069 = ( (~ i_20_)  &  (~ i_14_)  &  (~ i_12_)  &  (~ i_16_) ) ;
 assign wire7070 = ( (~ i_20_)  &  (~ i_14_)  &  (~ i_17_)  &  (~ i_16_) ) ;
 assign wire7046 = ( (~ i_30_)  &  (~ i_7_)  &  (~ i_8_)  &  (~ i_13_) ) ;
 assign wire1628 = ( n_n1375  &  n_n1322  &  wire246  &  wire7046 ) ;
 assign wire1632 = ( n_n1429  &  wire47  &  wire7058  &  wire7059 ) ;
 assign wire7054 = ( (~ i_20_)  &  (~ i_14_)  &  (~ i_17_)  &  (~ i_16_) ) ;
 assign wire1635 = ( n_n1213  &  wire7053  &  wire211  &  wire7054 ) ;
 assign wire1637 = ( n_n1441  &  n_n1408  &  wire77  &  wire7055 ) ;
 assign wire1640 = ( n_n1334  &  n_n1375  &  n_n1400  &  n_n1401 ) ;
 assign wire1651 = ( n_n1396  &  n_n1374  &  n_n1375  &  n_n1408 ) ;
 assign wire1652 = ( n_n1443  &  n_n1326  &  wire6947 ) ;
 assign wire1653 = ( n_n1390  &  wire305  &  wire717 ) ;
 assign wire7031 = ( i_7_  &  (~ i_14_)  &  (~ i_16_)  &  i_31_ ) ;
 assign wire1654 = ( n_n1441  &  n_n1400  &  wire7031 ) ;
 assign wire1656 = ( n_n1406  &  wire8  &  wire7025 ) ;
 assign wire1657 = ( n_n1443  &  n_n1369  &  n_n1368  &  wire7033 ) ;
 assign wire7028 = ( i_7_  &  (~ i_13_)  &  (~ i_16_)  &  i_31_ ) ;
 assign wire7026 = ( (~ i_32_)  &  (~ i_31_)  &  i_29_ ) ;
 assign wire7027 = ( (~ i_14_)  &  (~ i_12_)  &  (~ i_16_) ) | ( (~ i_14_)  &  (~ i_17_)  &  (~ i_16_) ) ;
 assign wire1668 = ( n_n1397  &  n_n1258  &  n_n1401  &  n_n1499 ) ;
 assign wire1675 = ( (~ i_28_)  &  i_25_  &  n_n1438  &  wire6948 ) ;
 assign wire1676 = ( n_n1216  &  wire6959  &  wire1677 ) | ( n_n1216  &  wire6959  &  wire1678 ) ;
 assign wire1670 = ( i_20_  &  wire1675 ) | ( i_20_  &  wire1676 ) ;
 assign wire6959 = ( (~ i_23_)  &  i_31_  &  i_34_ ) ;
 assign wire1672 = ( n_n1216  &  n_n1391  &  wire7017  &  wire6959 ) ;
 assign wire1677 = ( i_7_  &  (~ i_14_)  &  (~ i_17_)  &  (~ i_16_) ) ;
 assign wire1678 = ( i_7_  &  (~ i_14_)  &  (~ i_12_)  &  (~ i_16_) ) ;
 assign wire1684 = ( n_n1443  &  n_n1080  &  wire7009 ) ;
 assign wire1691 = ( n_n1443  &  n_n1396  &  n_n1374  &  n_n1375 ) ;
 assign wire1696 = ( n_n1318  &  n_n1497  &  n_n1311  &  n_n1459 ) ;
 assign wire6979 = ( (~ i_32_)  &  (~ i_31_)  &  i_29_ ) ;
 assign wire1698 = ( n_n1390  &  n_n1334  &  n_n1391  &  n_n1375 ) ;
 assign wire1699 = ( n_n1334  &  n_n1375  &  n_n1400  &  n_n1377 ) ;
 assign wire1700 = ( n_n1318  &  n_n1340  &  n_n1459  &  wire6982 ) ;
 assign wire1702 = ( n_n1433  &  n_n1312  &  wire6984 ) ;
 assign wire1703 = ( n_n1396  &  n_n1404  &  n_n1374  &  n_n1375 ) ;
 assign wire1704 = ( n_n1429  &  n_n1326  &  wire6947 ) ;
 assign wire6955 = ( (~ i_14_)  &  i_2_  &  (~ i_16_) ) ;
 assign wire1706 = ( n_n1369  &  n_n1274  &  n_n1368  &  wire6955 ) ;
 assign wire1709 = ( n_n1406  &  n_n1408  &  wire245 ) ;
 assign wire1710 = ( n_n1216  &  n_n1401  &  wire6960  &  wire6959 ) ;
 assign wire6971 = ( (~ i_7_)  &  i_34_  &  i_37_ ) ;
 assign wire6973 = ( (~ i_13_)  &  i_2_  &  (~ i_16_) ) ;
 assign wire1718 = ( n_n1369  &  n_n1274  &  n_n1368  &  wire6973 ) ;
 assign wire1719 = ( n_n1326  &  wire629  &  wire6947 ) ;
 assign wire6967 = ( (~ i_32_)  &  (~ i_31_)  &  (~ i_33_) ) ;
 assign wire1730 = ( n_n1307  &  n_n1408  &  wire635  &  wire6939 ) ;
 assign wire1731 = ( n_n1443  &  n_n504  &  n_n1118  &  n_n1279 ) ;
 assign wire1726 = ( n_n1375  &  n_n1213  &  wire1730 ) | ( n_n1375  &  n_n1213  &  wire1731 ) ;
 assign wire6939 = ( (~ i_32_)  &  (~ i_35_)  &  i_37_ ) ;
 assign wire1738 = ( n_n1018  &  n_n1302  &  _9463  &  _9466 ) ;
 assign wire6908 = ( (~ i_14_)  &  (~ i_11_)  &  (~ i_16_)  &  i_37_ ) ;
 assign wire1748 = ( wire1753  &  wire6912 ) | ( n_n21  &  wire6910  &  wire6912 ) ;
 assign wire1749 = ( wire606  &  _9922 ) ;
 assign wire1750 = ( n_n1443  &  n_n504  &  wire353  &  _9918 ) ;
 assign wire1747 = ( n_n26  &  wire1748 ) | ( n_n26  &  wire1749 ) | ( n_n26  &  wire1750 ) ;
 assign wire1753 = ( (~ i_14_)  &  wire44  &  wire6899  &  wire413 ) ;
 assign wire6910 = ( (~ i_14_)  &  (~ i_16_)  &  (~ i_32_) ) ;
 assign wire6912 = ( (~ i_9_)  &  i_37_  &  n_n1278 ) ;
 assign wire6884 = ( wire267  &  wire246 ) ;
 assign wire1756 = ( wire1766  &  wire6884 ) | ( n_n129  &  n_n130  &  wire6884 ) ;
 assign wire1757 = ( _860 ) | ( wire603  &  _9934 ) ;
 assign wire1758 = ( wire492  &  wire1767 ) | ( wire492  &  wire1768 ) ;
 assign wire6889 = ( n_n460  &  n_n1369  &  n_n1408  &  wire6885 ) ;
 assign wire6879 = ( (~ i_10_)  &  (~ i_13_)  &  (~ i_33_)  &  i_37_ ) ;
 assign wire6880 = ( (~ i_5_)  &  (~ i_4_)  &  (~ i_0_)  &  wire6879 ) ;
 assign wire6891 = ( (~ i_9_)  &  (~ i_8_)  &  (~ i_5_)  &  (~ i_6_) ) ;
 assign wire6898 = ( wire1756 ) | ( wire1758 ) | ( wire233  &  wire6880 ) ;
 assign wire6901 = ( (~ i_9_)  &  (~ i_14_)  &  i_37_  &  wire431 ) ;
 assign wire6903 = ( n_n841  &  n_n504  &  n_n245  &  n_n178 ) ;
 assign wire6905 = ( n_n1443  &  n_n504  &  n_n245  &  wire361 ) ;
 assign wire6917 = ( n_n18  &  wire6903 ) | ( wire63  &  wire6905 ) ;
 assign wire6919 = ( wire6917 ) | ( _9959 ) ;
 assign wire6922 = ( n_n1369  &  n_n504  &  n_n1288 ) ;
 assign wire6923 = ( (~ i_34_)  &  i_35_  &  (~ i_29_) ) ;
 assign wire6924 = ( (~ i_34_)  &  i_35_  &  (~ i_29_)  &  _9470 ) ;
 assign wire6926 = ( (~ i_32_)  &  (~ i_34_)  &  i_35_  &  wire365 ) ;
 assign wire6927 = ( i_34_  &  i_37_  &  n_n1216  &  n_n1305 ) ;
 assign wire6930 = ( n_n329  &  wire6922 ) | ( n_n363  &  wire6924 ) ;
 assign wire6931 = ( n_n620  &  wire6926 ) | ( n_n269  &  wire6927 ) ;
 assign wire6933 = ( wire6931 ) | ( (~ i_35_)  &  i_37_  &  wire600 ) ;
 assign wire6934 = ( wire1738 ) | ( wire6930 ) | ( n_n1295  &  wire601 ) ;
 assign wire6936 = ( wire267  &  wire246 ) ;
 assign wire6941 = ( n_n269  &  wire492 ) | ( n_n263  &  wire6936 ) ;
 assign wire6942 = ( wire6941 ) | ( wire634  &  _9498  &  _9499 ) ;
 assign wire6943 = ( wire1726 ) | ( wire248  &  wire632 ) ;
 assign wire6953 = ( i_20_  &  i_25_ ) ;
 assign wire6994 = ( (~ i_30_)  &  (~ i_35_)  &  (~ i_29_)  &  i_37_ ) ;
 assign wire7004 = ( (~ i_30_)  &  i_34_  &  (~ i_35_)  &  i_37_ ) ;
 assign wire7014 = ( (~ i_7_)  &  (~ i_14_)  &  (~ i_28_)  &  i_37_ ) ;
 assign wire7022 = ( wire1670 ) | ( _1082 ) | ( _1083 ) | ( _9399 ) ;
 assign wire7036 = ( wire1657 ) | ( n_n1396  &  wire6958  &  wire716 ) ;
 assign wire7037 = ( wire127 ) | ( wire1653 ) | ( wire1654 ) | ( wire1656 ) ;
 assign wire7040 = ( wire196 ) | ( _1114 ) | ( _1115 ) ;
 assign wire7041 = ( wire126 ) | ( wire1640 ) | ( wire1651 ) | ( wire1652 ) ;
 assign wire7043 = ( wire7036 ) | ( wire7037 ) | ( wire7040 ) | ( wire7041 ) ;
 assign wire7075 = ( wire1618 ) | ( n_n1369  &  wire515  &  _9607 ) ;
 assign wire7076 = ( wire1622 ) | ( n_n1441  &  n_n608  &  _9611 ) ;
 assign wire7079 = ( n_n793  &  wire29  &  wire7063 ) ;
 assign wire7085 = ( (~ i_35_)  &  i_37_  &  n_n1369  &  n_n1302 ) ;
 assign wire7087 = ( (~ i_35_)  &  i_37_  &  n_n1441  &  n_n1305 ) ;
 assign wire7089 = ( wire1607 ) | ( n_n571  &  n_n1311  &  wire7079 ) ;
 assign wire7090 = ( wire491  &  wire7085 ) | ( n_n544  &  wire7087 ) ;
 assign wire7093 = ( wire1608 ) | ( wire1611 ) | ( wire7089 ) | ( wire7090 ) ;
 assign wire7095 = ( (~ i_35_)  &  i_37_  &  n_n1375  &  n_n1340 ) ;
 assign wire7096 = ( (~ i_35_)  &  i_37_  &  n_n1369  &  n_n1288 ) ;
 assign wire7097 = ( (~ i_35_)  &  i_37_  &  n_n1375  &  n_n1213 ) ;
 assign wire7102 = ( n_n544  &  wire7095 ) | ( n_n437  &  wire7096 ) ;
 assign wire7103 = ( wire491  &  wire482 ) | ( n_n195  &  wire7097 ) ;
 assign wire7104 = ( wire7102 ) | ( wire7103 ) ;
 assign wire7114 = ( (~ i_30_)  &  i_34_  &  n_n504 ) ;
 assign wire7119 = ( (~ i_9_)  &  (~ i_10_)  &  (~ i_6_)  &  (~ i_32_) ) ;
 assign wire7134 = ( (~ i_35_)  &  i_37_  &  n_n841  &  n_n245 ) ;
 assign wire7135 = ( n_n1369  &  n_n1274  &  n_n1368  &  wire663 ) ;
 assign wire7137 = ( (~ i_10_)  &  i_37_ ) ;
 assign wire7139 = ( i_34_  &  i_37_  &  n_n1216  &  n_n1305 ) ;
 assign wire7140 = ( n_n1408  &  n_n839  &  wire6939 ) ;
 assign wire7141 = ( wire7134  &  wire7135 ) | ( wire88  &  wire7140 ) ;
 assign wire7142 = ( wire7141 ) | ( wire1767  &  wire7139 ) | ( wire1768  &  wire7139 ) ;
 assign wire7143 = ( wire1559 ) | ( n_n245  &  wire664  &  wire7137 ) ;
 assign wire7152 = ( n_n853  &  n_n1408  &  wire6939 ) ;
 assign wire7157 = ( wire1546 ) | ( wire1548 ) | ( wire88  &  wire7152 ) ;
 assign wire7165 = ( (~ i_34_)  &  i_35_  &  n_n793  &  n_n1305 ) ;
 assign wire7166 = ( n_n1307  &  n_n1100  &  n_n1340 ) ;
 assign wire7175 = ( (~ i_34_)  &  i_35_  &  i_37_ ) ;
 assign wire7179 = ( n_n1375  &  n_n1400  &  wire334 ) ;
 assign wire7190 = ( n_n1375  &  n_n1400  &  wire334 ) ;
 assign wire7203 = ( n_n1278  &  n_n152  &  wire258 ) ;
 assign wire7204 = ( n_n1375  &  n_n1322  &  _9851 ) ;
 assign wire7208 = ( (~ i_27_)  &  (~ i_28_)  &  (~ i_24_)  &  i_37_ ) ;
 assign wire7210 = ( n_n1322  &  n_n1241  &  wire7208 ) ;
 assign wire7211 = ( (~ i_14_)  &  (~ i_28_)  &  (~ i_16_)  &  (~ i_29_) ) ;
 assign wire7234 = ( wire1483 ) | ( _9896 ) | ( wire351  &  _9895 ) ;
 assign wire7238 = ( wire1511 ) | ( wire1549 ) | ( wire7157 ) | ( _9678 ) ;
 assign wire7239 = ( n_n1703 ) | ( n_n1704 ) | ( wire7142 ) | ( wire7143 ) ;
 assign wire7240 = ( wire1567 ) | ( n_n1701 ) | ( _9836 ) | ( _9899 ) ;
 assign wire7247 = ( wire6933 ) | ( wire6934 ) | ( wire6942 ) | ( wire6943 ) ;
 assign wire7248 = ( n_n1714 ) | ( n_n1713 ) | ( n_n1712 ) ;
 assign wire7256 = ( wire1747 ) | ( wire1757 ) | ( wire6898 ) | ( wire6919 ) ;
 assign wire7268 = ( (~ i_26_)  &  (~ i_24_)  &  i_38_ ) ;
 assign wire7269 = ( n_n1128  &  n_n1458  &  wire7268 ) ;
 assign wire7277 = ( i_9_  &  (~ i_8_)  &  i_12_ ) ;
 assign wire7286 = ( (~ i_28_)  &  (~ i_25_)  &  (~ i_26_)  &  _10870 ) ;
 assign wire7295 = ( (~ i_28_)  &  (~ i_25_)  &  (~ i_26_)  &  (~ i_29_) ) ;
 assign wire7306 = ( i_10_  &  i_19_  &  n_n584 ) ;
 assign wire7309 = ( n_n1437  &  n_n1133  &  wire7308 ) ;
 assign wire7312 = ( wire329  &  wire7306 ) | ( wire4  &  wire7309 ) ;
 assign wire7319 = ( i_9_  &  (~ i_10_)  &  (~ i_35_)  &  i_38_ ) ;
 assign wire7320 = ( n_n1118  &  n_n1279  &  wire7319 ) ;
 assign wire7321 = ( (~ i_28_)  &  (~ i_25_)  &  (~ i_26_)  &  _10962 ) ;
 assign wire7322 = ( n_n1279  &  n_n819  &  n_n1191 ) ;
 assign wire7323 = ( (~ i_33_)  &  i_38_  &  wire447 ) ;
 assign wire7325 = ( wire52  &  wire7320 ) | ( wire7321  &  wire7322 ) ;
 assign wire7327 = ( wire1399 ) | ( wire7325 ) | ( n_n706  &  wire7323 ) ;
 assign wire7328 = ( (~ i_32_)  &  (~ i_33_)  &  (~ i_35_)  &  i_38_ ) ;
 assign wire7329 = ( wire58  &  n_n1279  &  n_n819  &  n_n1191 ) ;
 assign wire7330 = ( (~ i_28_)  &  (~ i_25_)  &  (~ i_26_)  &  _10879 ) ;
 assign wire7331 = ( n_n1307  &  n_n841  &  n_n1191 ) ;
 assign wire7333 = ( i_9_  &  (~ i_10_)  &  n_n1118  &  n_n1279 ) ;
 assign wire7334 = ( (~ i_9_)  &  (~ i_6_)  &  i_13_  &  _10885 ) ;
 assign wire7335 = ( wire7328  &  wire7329 ) | ( wire7330  &  wire7331 ) ;
 assign wire7336 = ( wire390  &  wire7333 ) | ( n_n300  &  wire7334 ) ;
 assign wire7337 = ( wire261  &  wire379 ) | ( wire276  &  wire289 ) ;
 assign wire7339 = ( wire7335 ) | ( wire7336 ) | ( wire7337 ) ;
 assign wire7340 = ( (~ i_25_)  &  (~ i_26_)  &  (~ i_24_)  &  _10950 ) ;
 assign wire7341 = ( (~ i_9_)  &  (~ i_10_)  &  (~ i_6_)  &  _10948 ) ;
 assign wire7348 = ( n_n1861 ) | ( wire1403 ) | ( wire7327 ) ;
 assign wire7350 = ( wire1408 ) | ( wire7348 ) | ( _10942 ) | ( _10970 ) ;
 assign wire7351 = ( (~ i_30_)  &  (~ i_28_)  &  (~ i_2_)  &  (~ i_32_) ) ;
 assign wire7354 = ( (~ i_25_)  &  (~ i_24_)  &  n_n805  &  n_n1288 ) ;
 assign wire7355 = ( (~ i_32_)  &  (~ i_35_)  &  i_38_  &  wire78 ) ;
 assign wire7361 = ( (~ i_28_)  &  (~ i_26_)  &  n_n1191  &  wire226 ) ;
 assign wire7362 = ( (~ i_25_)  &  (~ i_24_)  &  n_n805  &  n_n1128 ) ;
 assign wire7363 = ( i_34_  &  (~ i_35_)  &  i_38_  &  _10679 ) ;
 assign wire7365 = ( (~ i_9_)  &  (~ i_6_)  &  i_13_  &  _10663 ) ;
 assign wire7366 = ( wire41  &  wire7361 ) | ( i_13_  &  wire41  &  wire7362 ) ;
 assign wire7367 = ( wire475  &  wire390 ) | ( wire394  &  wire7363 ) ;
 assign wire7368 = ( wire261  &  wire387 ) | ( n_n316  &  wire7365 ) ;
 assign wire7372 = ( (~ i_25_)  &  (~ i_24_)  &  n_n805  &  n_n1128 ) ;
 assign wire7373 = ( n_n1307  &  n_n1133  &  n_n839 ) ;
 assign wire7374 = ( (~ i_9_)  &  (~ i_10_)  &  (~ i_6_)  &  _10693 ) ;
 assign wire7379 = ( wire408  &  wire7372 ) | ( wire315  &  wire7373 ) ;
 assign wire7380 = ( i_13_  &  wire310 ) | ( n_n316  &  wire7374 ) ;
 assign wire7385 = ( n_n1197  &  n_n1133  &  n_n1497 ) ;
 assign wire7386 = ( (~ i_28_)  &  (~ i_25_)  &  (~ i_26_)  &  _10785 ) ;
 assign wire7387 = ( n_n1307  &  n_n853  &  n_n1128 ) ;
 assign wire7394 = ( wire218  &  wire7385 ) | ( wire270  &  wire7387 ) ;
 assign wire7395 = ( wire327  &  wire510 ) | ( n_n849  &  wire7386 ) ;
 assign wire7457 = ( i_10_  &  (~ i_3_)  &  n_n1438  &  n_n586 ) ;
 assign wire7458 = ( _526 ) | ( wire61  &  wire7457  &  _10628 ) ;
 assign wire7483 = ( wire1238 ) | ( wire1242 ) | ( _10534 ) ;
 assign wire7485 = ( wire1291 ) | ( wire7483 ) | ( _10526 ) | ( _10536 ) ;
 assign wire7510 = ( (~ i_24_)  &  (~ i_22_)  &  wire7265  &  wire264 ) ;
 assign wire7516 = ( (~ i_10_)  &  i_34_  &  wire239 ) | ( i_13_  &  i_34_  &  wire239 ) ;
 assign wire7521 = ( (~ i_5_)  &  (~ i_6_)  &  n_n1279  &  wire61 ) ;
 assign wire7525 = ( _763 ) | ( wire272  &  wire7516 ) ;
 assign wire7526 = ( _761 ) | ( (~ i_32_)  &  wire226  &  wire7521 ) ;
 assign wire7529 = ( wire7525 ) | ( wire7526 ) | ( _10184 ) ;
 assign wire7531 = ( (~ i_31_)  &  (~ i_29_)  &  n_n1118  &  n_n1279 ) ;
 assign wire7536 = ( n_n1307  &  n_n1144  &  wire264 ) ;
 assign wire7545 = ( (~ i_6_)  &  (~ i_12_)  &  n_n1307  &  wire61 ) ;
 assign wire7552 = ( n_n1489  &  n_n1458  &  wire7268 ) ;
 assign wire7553 = ( wire395  &  wire346 ) | ( wire744  &  wire7552 ) ;
 assign wire7555 = ( (~ i_25_)  &  i_38_ ) ;
 assign wire7567 = ( wire1176 ) | ( wire224  &  n_n1279  &  wire465 ) ;
 assign wire7574 = ( (~ i_10_)  &  wire503 ) ;
 assign wire7577 = ( (~ i_30_)  &  (~ i_28_)  &  (~ i_22_)  &  (~ i_31_) ) ;
 assign wire7580 = ( wire1159 ) | ( wire1161 ) | ( wire272  &  wire7574 ) ;
 assign wire7585 = ( (~ i_10_)  &  (~ i_32_)  &  n_n1307  &  n_n1100 ) ;
 assign wire7586 = ( n_n1118  &  n_n1279  &  n_n1128 ) ;
 assign wire7592 = ( wire1142 ) | ( wire1143 ) ;
 assign wire7595 = ( wire1139 ) | ( wire1140 ) | ( wire1141 ) | ( wire7592 ) ;
 assign wire7609 = ( wire1131 ) | ( wire1133 ) | ( wire1134 ) | ( wire1136 ) ;
 assign wire7621 = ( wire1112 ) | ( wire1113 ) | ( wire1114 ) ;
 assign wire7626 = ( (~ i_28_)  &  (~ i_24_)  &  i_22_  &  i_34_ ) ;
 assign wire7627 = ( i_30_  &  (~ i_28_)  &  (~ i_26_) ) | ( (~ i_28_)  &  (~ i_26_)  &  i_32_ ) ;
 assign wire7651 = ( wire1060 ) | ( wire1062 ) | ( _609 ) ;
 assign wire7676 = ( wire1032 ) | ( n_n1374  &  n_n1375  &  wire38 ) ;
 assign wire7678 = ( wire128 ) | ( wire1030 ) | ( wire1033 ) ;
 assign wire7689 = ( wire112 ) | ( wire1022 ) | ( n_n1397  &  wire734 ) ;
 assign wire7703 = ( (~ i_30_)  &  (~ i_8_)  &  (~ i_31_) ) ;
 assign wire7711 = ( n_n1881 ) | ( wire7651 ) | ( _10458 ) | ( _10460 ) ;
 assign wire7721 = ( (~ i_24_)  &  i_34_  &  (~ i_35_)  &  i_38_ ) ;
 assign wire7725 = ( n_n1307  &  n_n853  &  n_n1133 ) ;
 assign wire7726 = ( (~ i_5_)  &  (~ i_4_)  &  (~ i_2_)  &  _10731 ) ;
 assign wire7731 = ( (~ i_10_)  &  (~ i_24_)  &  n_n1279  &  n_n819 ) ;
 assign wire7732 = ( (~ i_28_)  &  (~ i_25_)  &  (~ i_26_)  &  _10746 ) ;
 assign wire7733 = ( i_34_  &  (~ i_35_)  &  i_38_  &  wire344 ) ;
 assign wire7734 = ( n_n1307  &  n_n1128  &  n_n839 ) ;
 assign wire7737 = ( wire394  &  wire7732 ) | ( wire327  &  wire7733 ) ;
 assign wire7738 = ( wire510  &  wire7731 ) | ( wire270  &  wire7734 ) ;
 assign wire7740 = ( wire977 ) | ( wire330  &  wire289 ) | ( wire330  &  wire978 ) ;
 assign wire7741 = ( wire7737 ) | ( wire7738 ) | ( _495 ) ;
 assign wire7743 = ( n_n1866 ) | ( n_n1865 ) | ( wire7740 ) | ( wire7741 ) ;
 assign wire7744 = ( n_n1827 ) | ( wire7743 ) ;
 assign wire7750 = ( (~ i_13_)  &  (~ i_32_)  &  i_36_  &  (~ i_35_) ) ;
 assign wire7763 = ( (~ i_14_)  &  i_13_  &  (~ i_16_)  &  wire232 ) ;
 assign wire7772 = ( (~ i_8_)  &  i_36_  &  (~ i_35_) ) ;
 assign wire7781 = ( wire942 ) | ( wire943 ) | ( wire232  &  wire568 ) ;
 assign wire7810 = ( i_31_  &  i_34_  &  wire80 ) ;
 assign wire7811 = ( (~ i_30_)  &  (~ i_28_)  &  (~ i_29_)  &  wire79 ) ;
 assign wire7817 = ( (~ i_9_)  &  i_2_  &  wire578 ) ;
 assign wire7823 = ( n_n355  &  wire418 ) | ( wire463  &  wire7817 ) ;
 assign wire7825 = ( wire7823 ) | ( wire86  &  wire576 ) ;
 assign wire7829 = ( (~ i_28_)  &  i_31_  &  (~ i_34_)  &  i_35_ ) ;
 assign wire7830 = ( (~ i_27_)  &  (~ i_23_)  &  i_21_  &  wire7829 ) ;
 assign wire7832 = ( (~ i_32_)  &  i_36_  &  n_n1441  &  wire7831 ) ;
 assign wire7834 = ( n_n1429  &  n_n1216  &  wire6959 ) ;
 assign wire7835 = ( (~ i_34_)  &  i_35_  &  (~ i_29_)  &  _11350 ) ;
 assign wire7836 = ( wire644  &  wire7830 ) | ( n_n458  &  wire7832 ) ;
 assign wire7837 = ( wire440  &  wire7834 ) | ( n_n363  &  wire7835 ) ;
 assign wire7838 = ( wire493  &  n_n620 ) | ( n_n242  &  wire418 ) ;
 assign wire7840 = ( wire7838 ) | ( i_34_  &  i_36_  &  wire643 ) ;
 assign wire7842 = ( (~ i_27_)  &  (~ i_28_)  &  i_31_  &  (~ i_29_) ) ;
 assign wire7843 = ( (~ i_23_)  &  (~ i_34_)  &  i_35_  &  wire541 ) ;
 assign wire7844 = ( wire437  &  wire7842 ) | ( wire891  &  wire7842 ) ;
 assign wire7845 = ( (~ i_32_)  &  i_36_  &  n_n1441  &  wire7831 ) ;
 assign wire7849 = ( wire7843  &  wire7844 ) | ( n_n358  &  wire7845 ) ;
 assign wire7852 = ( wire7849 ) | ( _11326 ) | ( n_n576  &  wire540 ) ;
 assign wire7853 = ( wire7825 ) | ( wire7840 ) | ( _11354 ) ;
 assign wire7854 = ( (~ i_27_)  &  (~ i_23_)  &  (~ i_17_)  &  i_36_ ) ;
 assign wire7855 = ( wire214  &  wire7854 ) ;
 assign wire7856 = ( n_n1441  &  wire265  &  wire7831 ) ;
 assign wire7857 = ( (~ i_27_)  &  (~ i_28_)  &  (~ i_31_) ) ;
 assign wire7863 = ( wire227  &  wire267 ) ;
 assign wire7864 = ( n_n355  &  wire7855 ) | ( n_n358  &  wire7863 ) ;
 assign wire7867 = ( n_n1369  &  n_n1128  &  n_n576 ) ;
 assign wire7869 = ( (~ i_32_)  &  (~ i_34_)  &  i_35_  &  wire267 ) ;
 assign wire7870 = ( (~ i_27_)  &  (~ i_23_)  &  (~ i_17_)  &  wire214 ) ;
 assign wire7879 = ( n_n437  &  wire483 ) | ( n_n195  &  wire500 ) ;
 assign wire7881 = ( wire849 ) | ( wire7879 ) | ( wire86  &  wire543 ) ;
 assign wire7885 = ( i_36_  &  (~ i_35_)  &  n_n1433  &  n_n1375 ) ;
 assign wire7888 = ( i_34_  &  i_36_  &  n_n1375  &  n_n1400 ) ;
 assign wire7889 = ( (~ i_27_)  &  (~ i_23_)  &  (~ i_24_)  &  _11363 ) ;
 assign wire7893 = ( n_n608  &  wire7885 ) | ( n_n242  &  wire7888 ) ;
 assign wire7895 = ( wire7893 ) | ( _107 ) | ( wire7887  &  _11366 ) ;
 assign wire7896 = ( i_31_  &  (~ i_34_)  &  i_35_  &  wire267 ) ;
 assign wire7897 = ( i_36_  &  (~ i_35_)  &  n_n1369  &  n_n1128 ) ;
 assign wire7899 = ( i_31_  &  i_34_  &  n_n1429  &  n_n1375 ) ;
 assign wire7902 = ( (~ i_26_)  &  (~ i_23_)  &  (~ i_24_)  &  _11361 ) ;
 assign wire7906 = ( wire669  &  wire7896 ) | ( wire491  &  wire7897 ) ;
 assign wire7907 = ( wire833 ) | ( n_n712  &  wire7898  &  wire7899 ) ;
 assign wire7909 = ( wire7906 ) | ( wire7907 ) | ( n_n1147  &  wire383 ) ;
 assign wire7910 = ( (~ i_32_)  &  i_36_  &  n_n1375  &  n_n1213 ) ;
 assign wire7911 = ( n_n1314  &  wire80  &  wire86 ) ;
 assign wire7912 = ( (~ i_34_)  &  i_35_  &  (~ i_29_)  &  _11296 ) ;
 assign wire7913 = ( (~ i_27_)  &  (~ i_28_)  &  (~ i_26_)  &  _11309 ) ;
 assign wire7914 = ( (~ i_32_)  &  (~ i_31_)  &  i_34_  &  _11307 ) ;
 assign wire7915 = ( n_n608  &  wire7913 ) | ( n_n544  &  wire7914 ) ;
 assign wire7918 = ( wire825 ) | ( n_n1089  &  wire383 ) ;
 assign wire7921 = ( wire834 ) | ( wire843 ) | ( wire7895 ) | ( wire7909 ) ;
 assign wire7932 = ( (~ i_27_)  &  (~ i_28_)  &  (~ i_26_)  &  i_33_ ) ;
 assign wire7935 = ( wire512 ) | ( wire38  &  wire7932 ) ;
 assign wire7936 = ( wire112 ) | ( wire507 ) | ( wire372  &  wire7029 ) ;
 assign wire7941 = ( (~ i_30_)  &  (~ i_31_)  &  n_n1375  &  wire86 ) ;
 assign wire7947 = ( i_36_  &  (~ i_35_)  &  n_n1369  &  n_n1254 ) ;
 assign wire7957 = ( (~ i_2_)  &  i_36_  &  n_n1443 ) ;
 assign wire7958 = ( n_n1441  &  wire77  &  wire7831 ) ;
 assign wire7959 = ( n_n1441  &  n_n1390  &  wire6993 ) ;
 assign wire7960 = ( (~ i_30_)  &  (~ i_31_)  &  wire258  &  wire86 ) ;
 assign wire7969 = ( i_20_  &  (~ i_28_)  &  (~ i_21_)  &  i_29_ ) ;
 assign wire7986 = ( (~ i_30_)  &  (~ i_31_)  &  wire259  &  wire86 ) ;
 assign wire7994 = ( i_36_  &  (~ i_35_)  &  wire259  &  n_n1459 ) ;
 assign wire8014 = ( wire178 ) | ( wire7947  &  _11113 ) ;
 assign wire8019 = ( i_36_  &  (~ i_35_)  &  n_n1441  &  n_n1133 ) ;
 assign wire8023 = ( wire163 ) | ( n_n544  &  wire8019 ) ;
 assign wire8026 = ( _11205 ) | ( i_36_  &  wire712 ) ;
 assign wire8027 = ( (~ i_27_)  &  (~ i_23_)  &  (~ i_24_)  &  i_34_ ) ;
 assign wire8028 = ( (~ i_28_)  &  i_31_  &  (~ i_29_)  &  wire8027 ) ;
 assign wire8029 = ( (~ i_2_)  &  i_36_  &  n_n1408 ) ;
 assign wire8030 = ( n_n1441  &  wire77  &  wire7831 ) ;
 assign wire8031 = ( (~ i_13_)  &  (~ i_17_)  &  (~ i_16_)  &  wire305 ) ;
 assign wire8039 = ( (~ i_13_)  &  (~ i_12_)  &  (~ i_16_)  &  wire305 ) ;
 assign wire8041 = ( (~ i_26_)  &  (~ i_23_)  &  (~ i_24_)  &  _11170 ) ;
 assign wire8077 = ( n_n1580 ) | ( n_n1579 ) | ( n_n1581 ) | ( n_n1583 ) ;
 assign wire8082 = ( (~ i_7_)  &  (~ i_11_)  &  (~ i_19_) ) ;
 assign wire8084 = ( (~ i_23_)  &  (~ i_21_)  &  wire232  &  wire8082 ) ;
 assign wire8093 = ( wire34 ) | ( wire462  &  wire8084 ) ;
 assign wire8094 = ( wire22 ) | ( _3 ) | ( _4 ) ;
 assign _3 = ( (~ i_21_)  &  wire462  &  wire338  &  wire8091 ) ;
 assign _4 = ( (~ i_21_)  &  wire105  &  wire8090 ) | ( (~ i_21_)  &  wire107  &  wire8090 ) ;
 assign _31 = ( (~ i_30_)  &  (~ i_28_)  &  wire245  &  wire8056 ) ;
 assign _32 = ( n_n1425  &  wire8056  &  _11495 ) ;
 assign _41 = ( n_n1404  &  n_n1312  &  wire6996  &  _11479 ) ;
 assign _42 = ( n_n1404  &  n_n1257  &  wire47  &  _9318 ) ;
 assign _43 = ( n_n1404  &  n_n1406  &  n_n1213  &  _9325 ) ;
 assign _62 = ( wire79  &  n_n1489  &  n_n1141  &  n_n1263 ) ;
 assign _63 = ( wire79  &  n_n1489  &  wire260  &  _11443 ) ;
 assign _64 = ( (~ i_28_)  &  i_31_  &  n_n1369  &  wire555 ) ;
 assign _67 = ( wire43  &  n_n1369  &  n_n1282  &  _11428 ) ;
 assign _75 = ( wire415  &  n_n1369  &  n_n1254  &  _11428 ) ;
 assign _77 = ( n_n1322  &  n_n1323  &  wire80  &  _11422 ) ;
 assign _78 = ( n_n1315  &  n_n1314  &  wire80  &  _11424 ) ;
 assign _79 = ( n_n1408  &  n_n1312  &  wire6996  &  _11419 ) ;
 assign _80 = ( n_n1408  &  n_n1257  &  wire47  &  _9318 ) ;
 assign _81 = ( n_n1406  &  n_n1213  &  wire7491  &  wire8 ) ;
 assign _82 = ( n_n1429  &  n_n1406  &  n_n1213  &  wire7491 ) ;
 assign _90 = ( i_22_  &  wire1663 ) | ( i_22_  &  _1089 ) | ( i_22_  &  _1090 ) ;
 assign _96 = ( (~ i_7_)  &  i_36_  &  wire214  &  _11391 ) ;
 assign _97 = ( n_n1433  &  n_n1489  &  _11393  &  _11395 ) ;
 assign _107 = ( wire610  &  wire6959  &  _11372 ) ;
 assign _180 = ( i_21_  &  wire189 ) | ( i_21_  &  _188 ) | ( i_21_  &  _189 ) ;
 assign _188 = ( (~ i_16_)  &  n_n1216  &  n_n1384  &  wire7999 ) ;
 assign _189 = ( (~ i_16_)  &  n_n1285  &  n_n1511  &  wire7997 ) ;
 assign _221 = ( i_21_  &  wire151 ) | ( i_21_  &  _231 ) | ( i_21_  &  _232 ) ;
 assign _231 = ( (~ i_17_)  &  wire47  &  n_n1387  &  wire7058 ) ;
 assign _232 = ( (~ i_17_)  &  n_n793  &  n_n1285  &  wire8043 ) ;
 assign _240 = ( (~ i_30_)  &  (~ i_31_)  &  n_n1202  &  wire7969 ) ;
 assign _278 = ( (~ i_13_)  &  (~ i_26_)  &  (~ i_23_)  &  (~ i_24_) ) ;
 assign _279 = ( (~ i_14_)  &  (~ i_26_)  &  (~ i_23_)  &  (~ i_24_) ) ;
 assign _282 = ( i_34_  &  i_36_  &  wire261  &  _11053 ) ;
 assign _283 = ( i_34_  &  i_36_  &  wire7178  &  _11056 ) ;
 assign _292 = ( n_n1408  &  n_n1118  &  n_n1279  &  _11029 ) ;
 assign _293 = ( n_n461  &  wire265  &  wire7819  &  _11033 ) ;
 assign _294 = ( i_36_  &  wire956 ) | ( i_36_  &  wire958 ) | ( i_36_  &  _11024 ) ;
 assign _303 = ( i_36_  &  wire966 ) | ( i_36_  &  wire967 ) | ( i_36_  &  _10999 ) ;
 assign _322 = ( wire404  &  n_n1300  &  wire61  &  _10475 ) ;
 assign _335 = ( n_n1128  &  wire239  &  wire624  &  _10933 ) ;
 assign _336 = ( n_n1128  &  _338 ) | ( n_n1128  &  wire521  &  _10937 ) ;
 assign _338 = ( (~ i_24_)  &  wire404  &  wire7274  &  wire7311 ) ;
 assign _342 = ( wire404  &  n_n1419  &  wire344  &  _10475 ) ;
 assign _343 = ( (~ i_33_)  &  i_38_  &  wire406  &  _10918 ) ;
 assign _363 = ( wire7332  &  _364 ) | ( wire7332  &  _365 ) ;
 assign _364 = ( n_n1307  &  n_n1100  &  _10667  &  _10876 ) ;
 assign _365 = ( wire404  &  _10475  &  _10877 ) ;
 assign _390 = ( n_n586  &  wire7272  &  _10317  &  _10846 ) ;
 assign _400 = ( n_n316  &  _10828 ) | ( n_n316  &  _10829 ) ;
 assign _401 = ( n_n1523  &  wire423  &  _9998 ) ;
 assign _402 = ( n_n300  &  _10826 ) | ( n_n300  &  _10827 ) ;
 assign _406 = ( i_19_  &  n_n1118  &  n_n1279  &  n_n1048 ) ;
 assign _407 = ( i_19_  &  n_n461  &  wire7411  &  n_n1028 ) ;
 assign _410 = ( wire434  &  wire78  &  _10816 ) | ( wire78  &  _411  &  _10816 ) ;
 assign _411 = ( n_n1118  &  n_n1058  &  wire7415 ) ;
 assign _415 = ( n_n1523  &  _418  &  _9998 ) | ( n_n1523  &  _419  &  _9998 ) ;
 assign _418 = ( i_19_  &  wire7419  &  wire7420  &  _10491 ) ;
 assign _419 = ( i_19_  &  n_n1307  &  n_n1048  &  n_n1144 ) ;
 assign _439 = ( i_38_  &  wire627 ) ;
 assign _442 = ( (~ i_24_)  &  i_38_  &  wire78  &  wire346 ) ;
 assign _451 = ( n_n1197  &  wire1349 ) | ( n_n1197  &  wire1350 ) | ( n_n1197  &  wire1351 ) ;
 assign _460 = ( n_n1100  &  wire311  &  _9748  &  _10762 ) ;
 assign _490 = ( n_n1100  &  n_n1419  &  _9748  &  _10651 ) ;
 assign _495 = ( n_n853  &  wire7547  &  _9996  &  _10754 ) ;
 assign _510 = ( n_n819  &  wire344  &  wire7721  &  _10648 ) ;
 assign _526 = ( wire381  &  _10631 ) | ( wire381  &  _10632 ) ;
 assign _530 = ( i_19_  &  n_n1118  &  n_n1279  &  n_n1048 ) ;
 assign _531 = ( i_19_  &  n_n461  &  wire7411  &  n_n1028 ) ;
 assign _539 = ( wire254  &  _10606 ) | ( wire254  &  _10607 ) ;
 assign _543 = ( n_n1307  &  wire7423  &  wire381  &  _10524 ) ;
 assign _585 = ( wire430  &  _588  &  _10496 ) | ( wire430  &  _589  &  _10496 ) ;
 assign _588 = ( i_19_  &  wire7419  &  wire7420  &  _10491 ) ;
 assign _589 = ( i_19_  &  n_n1307  &  n_n1048  &  n_n1144 ) ;
 assign _595 = ( wire404  &  wire429  &  _10475  &  _10477 ) ;
 assign _606 = ( n_n1279  &  wire7266  &  _10425  &  _10457 ) ;
 assign _609 = ( n_n1307  &  n_n1303  &  wire78  &  _10324 ) ;
 assign _612 = ( n_n1425  &  n_n1197  &  n_n1192  &  _10445 ) ;
 assign _613 = ( n_n1478  &  n_n1192  &  _10445  &  _10448 ) ;
 assign _614 = ( n_n1306  &  wire7265  &  _10038  &  _10160 ) ;
 assign _615 = ( n_n1279  &  wire7265  &  _10160  &  _10176 ) ;
 assign _617 = ( n_n1307  &  n_n1303  &  wire288  &  _10324 ) ;
 assign _624 = ( n_n1454  &  n_n1279  &  _10176  &  _10430 ) ;
 assign _626 = ( n_n1306  &  wire7266  &  _10425  &  _10426 ) ;
 assign _627 = ( n_n1303  &  wire7266  &  _10034  &  _10425 ) ;
 assign _635 = ( n_n1225  &  n_n1303  &  wire239  &  _10034 ) ;
 assign _637 = ( wire71  &  wire12  &  wire7703 ) ;
 assign _655 = ( n_n1489  &  wire226  &  wire7704 ) ;
 assign _656 = ( n_n1489  &  n_n1179  &  _10377 ) ;
 assign _657 = ( i_38_  &  wire1017 ) | ( i_38_  &  _662 ) ;
 assign _658 = ( i_38_  &  _664 ) | ( i_38_  &  _665 ) ;
 assign _662 = ( n_n1439  &  n_n1438  &  n_n1437 ) ;
 assign _664 = ( (~ i_2_)  &  n_n1425  &  wire7276  &  _10370 ) ;
 assign _665 = ( (~ i_2_)  &  n_n1454  &  n_n1431  &  _10372 ) ;
 assign _668 = ( (~ i_32_)  &  n_n1425  &  wire226  &  _10341 ) ;
 assign _674 = ( n_n1454  &  n_n1306  &  n_n1288  &  _10038 ) ;
 assign _676 = ( n_n1305  &  n_n1306  &  n_n1497  &  _10038 ) ;
 assign _677 = ( n_n1305  &  n_n1279  &  n_n1497  &  _10176 ) ;
 assign _678 = ( (~ i_33_)  &  i_38_  &  n_n1425  &  _10313 ) ;
 assign _679 = ( (~ i_33_)  &  i_38_  &  wire7272  &  _10317 ) ;
 assign _683 = ( n_n805  &  n_n1466  &  n_n1359  &  _10290 ) ;
 assign _684 = ( n_n1478  &  n_n1472  &  n_n1359  &  _10292 ) ;
 assign _685 = ( n_n1489  &  n_n1340  &  n_n1359  &  _10294 ) ;
 assign _686 = ( n_n1454  &  n_n1489  &  n_n1353  &  _10286 ) ;
 assign _702 = ( wire447  &  wire35 ) ;
 assign _733 = ( i_27_  &  i_22_  &  _10216 ) | ( i_16_  &  i_22_  &  _10216 ) ;
 assign _744 = ( i_12_  &  (~ i_24_)  &  i_17_ ) ;
 assign _746 = ( (~ i_28_)  &  i_32_  &  i_34_  &  (~ i_29_) ) ;
 assign _747 = ( i_30_  &  (~ i_28_)  &  i_34_  &  (~ i_29_) ) ;
 assign _749 = ( i_30_  &  wire298  &  wire345 ) | ( i_32_  &  wire298  &  wire345 ) ;
 assign _750 = ( (~ i_24_)  &  i_34_  &  n_n1489  &  _10205 ) ;
 assign _756 = ( i_34_  &  n_n1489  &  wire239  &  _10190 ) ;
 assign _757 = ( i_34_  &  n_n1466  &  wire77  &  _10192 ) ;
 assign _758 = ( i_34_  &  wire7612  &  _10197 ) ;
 assign _761 = ( n_n1279  &  n_n1523  &  _9998  &  _10181 ) ;
 assign _763 = ( n_n1279  &  wire214  &  _10176  &  _10177 ) ;
 assign _767 = ( n_n1307  &  n_n1303  &  _9684  &  _10171 ) ;
 assign _781 = ( n_n1454  &  n_n1279  &  wire446  &  _10133 ) ;
 assign _782 = ( n_n1100  &  n_n1191  &  _9748  &  _10137 ) ;
 assign _788 = ( n_n1438  &  n_n1197  &  wire61  &  _10108 ) ;
 assign _789 = ( n_n1197  &  n_n1523  &  wire7466  &  _10112 ) ;
 assign _791 = ( n_n1307  &  n_n1144  &  wire226  &  wire457 ) ;
 assign _795 = ( i_9_  &  i_12_  &  wire1168 ) | ( i_9_  &  i_12_  &  _797 ) ;
 assign _796 = ( i_9_  &  i_12_  &  _799 ) | ( i_9_  &  i_12_  &  _800 ) ;
 assign _797 = ( n_n1454  &  n_n1179  &  wire7577 ) ;
 assign _799 = ( (~ i_10_)  &  n_n1425  &  n_n1179  &  wire7276 ) ;
 assign _800 = ( (~ i_10_)  &  n_n1197  &  n_n1523  &  n_n1431 ) ;
 assign _803 = ( n_n1144  &  wire7547  &  _9996  &  _10073 ) ;
 assign _816 = ( n_n1466  &  n_n1306  &  _10038  &  _10041 ) ;
 assign _817 = ( n_n1454  &  n_n1307  &  wire446  &  _10045 ) ;
 assign _818 = ( n_n1303  &  wire214  &  wire7555  &  _10034 ) ;
 assign _820 = ( n_n1486  &  wire18  &  n_n998  &  wire7559 ) ;
 assign _821 = ( (~ i_24_)  &  wire436  &  wire71  &  wire7559 ) ;
 assign _822 = ( n_n1307  &  n_n1303  &  n_n1059  &  _10022 ) ;
 assign _823 = ( n_n1307  &  n_n1306  &  n_n1288  &  n_n1059 ) ;
 assign _832 = ( n_n1144  &  _9999  &  _10004 ) ;
 assign _833 = ( (~ i_24_)  &  (~ i_29_)  &  wire223  &  wire311 ) ;
 assign _834 = ( n_n1279  &  wire7547  &  _9992  &  _9996 ) ;
 assign _835 = ( n_n1144  &  n_n1523  &  _9998  &  _9999 ) ;
 assign _844 = ( (~ i_33_)  &  i_37_  &  n_n18  &  _9913 ) ;
 assign _860 = ( (~ i_35_)  &  i_37_  &  wire604  &  wire6889 ) ;
 assign _881 = ( n_n1408  &  wire484  &  wire7219 ) | ( n_n1408  &  wire489  &  wire7219 ) ;
 assign _899 = ( n_n245  &  wire233  &  _9834 ) ;
 assign _927 = ( n_n1295  &  wire85  &  wire7178 ) | ( n_n1295  &  wire85  &  wire7179 ) ;
 assign _928 = ( i_34_  &  i_37_  &  wire261  &  _9754 ) ;
 assign _929 = ( i_34_  &  i_37_  &  wire223  &  _9755 ) ;
 assign _963 = ( n_n1213  &  _9659  &  _9674 ) ;
 assign _975 = ( i_37_  &  wire1634 ) | ( i_37_  &  _1002 ) | ( i_37_  &  _1003 ) ;
 assign _983 = ( wire7053  &  wire7084  &  wire7083  &  _9619 ) ;
 assign _993 = ( wire7072  &  _995 ) | ( wire7072  &  _996 ) ;
 assign _995 = ( n_n1431  &  wire7068  &  wire7069 ) ;
 assign _996 = ( wire7053  &  wire7069  &  _9404 ) ;
 assign _1002 = ( (~ i_0_)  &  wire1635 ) | ( (~ i_0_)  &  wire1637 ) ;
 assign _1003 = ( (~ i_0_)  &  _1005 ) | ( (~ i_0_)  &  _1006 ) ;
 assign _1005 = ( n_n1404  &  n_n1213  &  wire7053  &  _9644 ) ;
 assign _1006 = ( n_n1441  &  n_n1404  &  wire77  &  wire7055 ) ;
 assign _1015 = ( wire260  &  wire77  &  wire365  &  _9551 ) ;
 assign _1016 = ( n_n1263  &  wire365  &  _9551  &  _9553 ) ;
 assign _1020 = ( wire47  &  wire1678  &  _9542 ) ;
 assign _1021 = ( wire47  &  wire1677  &  _9542 ) ;
 assign _1027 = ( n_n1216  &  n_n1141  &  n_n1263  &  _9351 ) ;
 assign _1070 = ( wire7053  &  wire402  &  _9404  &  _9408 ) ;
 assign _1074 = ( n_n1404  &  n_n1406  &  wire245 ) ;
 assign _1076 = ( n_n1202  &  n_n1459  &  wire7014 ) ;
 assign _1082 = ( n_n1408  &  n_n1257  &  wire47  &  _9318 ) ;
 assign _1083 = ( n_n1408  &  wire6996  &  wire6997  &  _9322 ) ;
 assign _1084 = ( i_22_  &  wire1663 ) | ( i_22_  &  _1089 ) | ( i_22_  &  _1090 ) ;
 assign _1089 = ( wire54  &  wire44  &  wire29 ) | ( wire54  &  wire44  &  wire7027 ) ;
 assign _1090 = ( (~ i_23_)  &  (~ i_24_)  &  wire6984  &  _9379 ) ;
 assign _1098 = ( n_n1375  &  n_n1400  &  wire258  &  wire7004 ) ;
 assign _1099 = ( n_n1390  &  n_n1375  &  wire6993  &  wire7004 ) ;
 assign _1102 = ( n_n1216  &  wire260  &  _9351  &  _9354 ) ;
 assign _1103 = ( n_n1429  &  n_n1080  &  wire7009 ) ;
 assign _1104 = ( n_n1396  &  n_n1429  &  n_n1375  &  _9344 ) ;
 assign _1105 = ( n_n1441  &  n_n1400  &  wire258  &  wire6994 ) ;
 assign _1106 = ( n_n1441  &  n_n1390  &  wire6993  &  wire6994 ) ;
 assign _1108 = ( n_n1404  &  n_n1257  &  wire47  &  _9318 ) ;
 assign _1109 = ( n_n1404  &  wire6996  &  wire6997  &  _9322 ) ;
 assign _1110 = ( n_n1258  &  n_n1499  &  n_n1377  &  _9309 ) ;
 assign _1111 = ( n_n1499  &  n_n1251  &  wire661  &  _9314 ) ;
 assign _1114 = ( n_n1369  &  wire8  &  wire7033  &  _9290 ) ;
 assign _1115 = ( n_n1369  &  n_n1429  &  wire7033  &  _9290 ) ;
 assign _1134 = ( n_n1439  &  n_n1438  &  wire6971  &  _9202 ) ;
 assign _1135 = ( n_n1489  &  wire6971  &  wire6967  &  _9206 ) ;
 assign _9202 = ( (~ i_23_)  &  (~ i_14_) ) ;
 assign _9206 = ( (~ i_24_)  &  (~ i_23_) ) ;
 assign _9225 = ( wire1715 ) | ( wire1717 ) | ( _1134 ) | ( _1135 ) ;
 assign _9227 = ( (~ i_24_)  &  i_21_  &  (~ i_34_) ) ;
 assign _9290 = ( i_29_  &  (~ i_28_) ) ;
 assign _9309 = ( i_35_  &  (~ i_34_) ) ;
 assign _9314 = ( i_35_  &  (~ i_34_) ) ;
 assign _9318 = ( i_25_  &  (~ i_27_) ) ;
 assign _9322 = ( i_33_  &  i_34_ ) ;
 assign _9325 = ( (~ i_20_)  &  i_2_  &  (~ i_21_) ) ;
 assign _9328 = ( (~ i_13_)  &  (~ i_12_)  &  (~ i_16_) ) ;
 assign _9338 = ( wire1690 ) | ( _1110 ) | ( _1111 ) ;
 assign _9344 = ( i_33_  &  i_34_ ) ;
 assign _9347 = ( (~ i_14_)  &  (~ i_12_)  &  (~ i_16_) ) ;
 assign _9351 = ( (~ i_30_)  &  i_34_  &  (~ i_29_)  &  i_37_ ) ;
 assign _9354 = ( (~ i_8_)  &  (~ i_7_) ) ;
 assign _9361 = ( wire1683 ) | ( _1103 ) | ( _1104 ) ;
 assign _9379 = ( (~ i_32_)  &  (~ i_31_)  &  i_34_ ) ;
 assign _9399 = ( wire1668 ) | ( wire1672 ) | ( _1074 ) | ( _1076 ) ;
 assign _9404 = ( (~ i_8_)  &  (~ i_26_)  &  (~ i_23_)  &  (~ i_24_) ) ;
 assign _9408 = ( (~ i_33_)  &  (~ i_35_)  &  i_37_ ) ;
 assign _9409 = ( i_37_  &  (~ i_33_) ) ;
 assign _9456 = ( (~ i_27_)  &  (~ i_28_)  &  (~ i_24_) ) ;
 assign _9459 = ( (~ i_27_)  &  (~ i_23_)  &  (~ i_24_) ) ;
 assign _9463 = ( i_37_  &  i_34_ ) ;
 assign _9466 = ( n_n1429  &  n_n1307  &  n_n1303 ) ;
 assign _9470 = ( (~ i_27_)  &  (~ i_28_)  &  (~ i_23_)  &  i_37_ ) ;
 assign _9480 = ( (~ i_28_)  &  (~ i_32_)  &  (~ i_29_) ) ;
 assign _9483 = ( (~ i_27_)  &  (~ i_28_)  &  (~ i_29_) ) ;
 assign _9494 = ( (~ i_5_)  &  (~ i_4_)  &  (~ i_2_) ) ;
 assign _9495 = ( (~ i_27_)  &  (~ i_28_)  &  (~ i_26_)  &  (~ i_29_) ) ;
 assign _9498 = ( i_37_  &  (~ i_35_) ) ;
 assign _9499 = ( n_n841  &  n_n1400  &  _9494  &  _9495 ) ;
 assign _9511 = ( (~ i_32_)  &  (~ i_33_)  &  (~ i_29_) ) ;
 assign _9514 = ( (~ i_28_)  &  (~ i_33_)  &  (~ i_29_) ) ;
 assign _9542 = ( i_20_  &  (~ i_27_)  &  (~ i_28_)  &  i_31_ ) ;
 assign _9551 = ( i_35_  &  (~ i_34_) ) ;
 assign _9553 = ( (~ i_30_)  &  (~ i_7_)  &  (~ i_8_)  &  (~ i_12_) ) ;
 assign _9577 = ( i_34_  &  (~ i_35_)  &  i_37_  &  wire80 ) ;
 assign _9583 = ( (~ i_32_)  &  i_34_  &  (~ i_35_) ) ;
 assign _9584 = ( wire1632 ) | ( n_n608  &  wire365  &  _9583 ) ;
 assign _9587 = ( (~ i_8_)  &  (~ i_26_)  &  (~ i_23_)  &  (~ i_24_) ) ;
 assign _9598 = ( wire1623  &  wire7072 ) | ( wire1625  &  wire7072 ) ;
 assign _9607 = ( (~ i_28_)  &  (~ i_35_)  &  (~ i_29_)  &  i_37_ ) ;
 assign _9611 = ( (~ i_32_)  &  (~ i_35_)  &  (~ i_29_)  &  i_37_ ) ;
 assign _9613 = ( (~ i_30_)  &  (~ i_28_)  &  (~ i_32_) ) ;
 assign _9616 = ( n_n1369  &  wire7084  &  _9613 ) ;
 assign _9619 = ( (~ i_8_)  &  (~ i_26_)  &  (~ i_23_)  &  (~ i_24_) ) ;
 assign _9621 = ( (~ i_27_)  &  (~ i_23_)  &  (~ i_24_)  &  i_37_ ) ;
 assign _9636 = ( wire7075 ) | ( wire7076 ) | ( _993 ) | ( _9598 ) ;
 assign _9644 = ( (~ i_20_)  &  (~ i_7_)  &  (~ i_32_) ) ;
 assign _9652 = ( n_n1018  &  wire248  &  _9480 ) ;
 assign _9659 = ( (~ i_20_)  &  (~ i_27_)  &  (~ i_28_)  &  i_29_ ) ;
 assign _9673 = ( (~ i_7_)  &  (~ i_6_)  &  (~ i_12_) ) ;
 assign _9674 = ( wire268  &  wire7161  &  _9673 ) ;
 assign _9678 = ( wire1509 ) | ( _963 ) | ( wire708  &  wire7188 ) ;
 assign _9683 = ( (~ i_34_)  &  i_35_  &  n_n301  &  n_n1258 ) ;
 assign _9684 = ( (~ i_10_)  &  (~ i_9_) ) ;
 assign _9686 = ( i_35_  &  (~ i_34_) ) ;
 assign _9688 = ( (~ i_13_)  &  n_n1307  &  n_n1303  &  _9684 ) ;
 assign _9724 = ( (~ i_5_)  &  (~ i_4_)  &  (~ i_0_) ) ;
 assign _9733 = ( n_n1306  &  wire7161  &  wire7163 ) ;
 assign _9736 = ( wire508  &  wire470 ) | ( wire222  &  _9733 ) ;
 assign _9737 = ( i_35_  &  (~ i_34_) ) ;
 assign _9740 = ( n_n1278  &  n_n1279  &  wire259 ) ;
 assign _9748 = ( (~ i_5_)  &  (~ i_4_)  &  (~ i_2_)  &  (~ i_32_) ) ;
 assign _9751 = ( i_13_  &  (~ i_9_) ) ;
 assign _9753 = ( (~ i_14_)  &  (~ i_23_)  &  (~ i_17_)  &  (~ i_16_) ) ;
 assign _9754 = ( _9753  &  wire80 ) ;
 assign _9755 = ( wire80  &  wire260 ) ;
 assign _9758 = ( (~ i_10_)  &  (~ i_13_)  &  (~ i_16_) ) ;
 assign _9760 = ( n_n1307  &  n_n841  &  n_n504  &  _9758 ) ;
 assign _9781 = ( (~ i_9_)  &  (~ i_13_)  &  (~ i_11_) ) ;
 assign _9784 = ( n_n1307  &  n_n1303  &  n_n130  &  _9781 ) ;
 assign _9804 = ( n_n245  &  wire44  &  wire6899 ) ;
 assign _9821 = ( (~ i_9_)  &  (~ i_5_)  &  (~ i_4_)  &  (~ i_2_) ) ;
 assign _9834 = ( (~ i_14_)  &  i_13_  &  i_37_ ) ;
 assign _9836 = ( wire1565 ) | ( wire1566 ) | ( wire7120  &  _9804 ) ;
 assign _9847 = ( (~ i_14_)  &  (~ i_34_)  &  i_35_  &  n_n1322 ) ;
 assign _9851 = ( (~ i_14_)  &  (~ i_34_)  &  i_35_ ) ;
 assign _9857 = ( (~ i_34_)  &  i_35_  &  n_n1258  &  n_n916 ) ;
 assign _9868 = ( (~ i_5_)  &  (~ i_6_)  &  n_n152  &  wire7215 ) ;
 assign _9872 = ( (~ i_32_)  &  (~ i_35_)  &  (~ i_29_)  &  i_37_ ) ;
 assign _9876 = ( (~ i_34_)  &  i_35_  &  n_n1258  &  wire7216 ) ;
 assign _9880 = ( (~ i_13_)  &  n_n1307  &  n_n1303  &  _9684 ) ;
 assign _9882 = ( wire1490 ) | ( wire7221 ) | ( wire7214  &  _9868 ) ;
 assign _9889 = ( (~ i_20_)  &  (~ i_23_)  &  (~ i_24_)  &  wire44 ) ;
 assign _9890 = ( i_37_  &  (~ i_13_) ) ;
 assign _9892 = ( wire224  &  n_n152  &  n_n1458  &  _9890 ) ;
 assign _9895 = ( (~ i_32_)  &  i_34_  &  (~ i_29_)  &  n_n1216 ) ;
 assign _9896 = ( wire7224  &  _9889 ) | ( wire7214  &  _9892 ) ;
 assign _9898 = ( wire1484 ) | ( wire1576  &  wire7230 ) | ( wire1577  &  wire7230 ) ;
 assign _9899 = ( wire1493 ) | ( wire7234 ) | ( _9882 ) | ( _9898 ) ;
 assign _9901 = ( wire7238 ) | ( n_n1690 ) ;
 assign _9907 = ( (~ i_9_)  &  (~ i_13_)  &  (~ i_33_)  &  i_37_ ) ;
 assign _9908 = ( (~ i_20_)  &  (~ i_17_)  &  (~ i_19_) ) ;
 assign _9913 = ( n_n245  &  n_n178  &  wire6906 ) ;
 assign _9918 = ( (~ i_20_)  &  (~ i_23_)  &  n_n460  &  n_n1369 ) ;
 assign _9919 = ( (~ i_20_)  &  (~ i_18_)  &  (~ i_17_) ) ;
 assign _9922 = ( n_n1406  &  n_n180  &  n_n1213  &  _9919 ) ;
 assign _9929 = ( (~ i_9_)  &  (~ i_8_)  &  (~ i_6_)  &  (~ i_11_) ) ;
 assign _9934 = ( (~ i_14_)  &  (~ i_16_)  &  (~ i_35_)  &  i_37_ ) ;
 assign _9950 = ( n_n245  &  wire6906  &  wire6908 ) ;
 assign _9959 = ( wire508  &  wire6901 ) | ( n_n18  &  _9950 ) ;
 assign _9963 = ( wire7250 ) | ( wire7257 ) | ( wire7044 ) | ( wire7045 ) ;
 assign _9992 = ( (~ i_8_)  &  (~ i_5_)  &  (~ i_6_) ) ;
 assign _9996 = ( (~ i_31_)  &  i_34_  &  (~ i_35_)  &  i_38_ ) ;
 assign _9998 = ( (~ i_28_)  &  (~ i_33_)  &  (~ i_35_)  &  i_38_ ) ;
 assign _9999 = ( (~ i_5_)  &  (~ i_4_)  &  (~ i_2_)  &  (~ i_31_) ) ;
 assign _10003 = ( (~ i_28_)  &  (~ i_25_)  &  (~ i_24_) ) ;
 assign _10004 = ( (~ i_29_)  &  n_n805  &  _10003 ) ;
 assign _10022 = ( (~ i_28_)  &  (~ i_12_)  &  (~ i_29_) ) ;
 assign _10025 = ( _823 ) | ( _822 ) ;
 assign _10034 = ( (~ i_5_)  &  (~ i_4_)  &  (~ i_12_)  &  (~ i_2_) ) ;
 assign _10038 = ( (~ i_5_)  &  (~ i_4_)  &  (~ i_2_)  &  i_38_ ) ;
 assign _10041 = ( (~ i_32_)  &  (~ i_34_)  &  i_35_ ) ;
 assign _10045 = ( (~ i_6_)  &  (~ i_28_)  &  (~ i_12_)  &  (~ i_22_) ) ;
 assign _10051 = ( wire1173 ) | ( _818 ) | ( _820 ) | ( _821 ) ;
 assign _10053 = ( wire7553 ) | ( _832 ) | ( _833 ) | ( _10025 ) ;
 assign _10062 = ( wire503  &  i_13_ ) ;
 assign _10073 = ( (~ i_5_)  &  (~ i_4_)  &  (~ i_2_) ) ;
 assign _10075 = ( wire7588 ) | ( wire1152 ) | ( wire272  &  _10062 ) ;
 assign _10085 = ( (~ i_8_)  &  (~ i_31_)  &  (~ i_35_)  &  i_38_ ) ;
 assign _10108 = ( i_12_  &  i_9_ ) ;
 assign _10112 = ( i_12_  &  i_9_ ) ;
 assign _10125 = ( wire1162 ) | ( wire7580 ) | ( _795 ) | ( _796 ) ;
 assign _10130 = ( n_n1437  &  n_n1472  &  wire7308 ) ;
 assign _10132 = ( (~ i_24_)  &  i_34_  &  i_38_  &  n_n1466 ) ;
 assign _10133 = ( (~ i_5_)  &  (~ i_6_)  &  (~ i_28_)  &  (~ i_22_) ) ;
 assign _10137 = ( (~ i_28_)  &  (~ i_26_)  &  (~ i_33_)  &  i_38_ ) ;
 assign _10142 = ( i_38_  &  (~ i_33_) ) ;
 assign _10143 = ( wire529  &  _10130 ) | ( wire261  &  _10132 ) ;
 assign _10151 = ( (~ i_24_)  &  i_34_  &  i_38_ ) ;
 assign _10160 = ( (~ i_22_)  &  (~ i_24_) ) ;
 assign _10169 = ( (~ i_7_)  &  (~ i_5_)  &  (~ i_6_)  &  i_38_ ) ;
 assign _10171 = ( (~ i_24_)  &  i_34_  &  i_38_ ) ;
 assign _10173 = ( (~ i_28_)  &  (~ i_25_)  &  (~ i_29_) ) ;
 assign _10175 = ( (~ i_24_)  &  i_34_  &  i_38_  &  n_n1302 ) ;
 assign _10176 = ( (~ i_7_)  &  (~ i_5_)  &  (~ i_6_)  &  i_38_ ) ;
 assign _10177 = ( (~ i_25_)  &  (~ i_8_) ) ;
 assign _10181 = ( (~ i_8_)  &  (~ i_5_)  &  (~ i_6_)  &  (~ i_31_) ) ;
 assign _10184 = ( i_13_  &  wire286 ) | ( wire261  &  _10175 ) ;
 assign _10186 = ( wire7511 ) | ( wire7512 ) | ( wire1211 ) | ( _10143 ) ;
 assign _10188 = ( wire7591 ) | ( wire7595 ) | ( _10075 ) | ( _10125 ) ;
 assign _10190 = ( (~ i_32_)  &  (~ i_7_) ) ;
 assign _10192 = ( i_38_  &  (~ i_24_) ) ;
 assign _10197 = ( i_12_  &  (~ i_24_)  &  i_17_ ) ;
 assign _10205 = ( (~ i_7_)  &  (~ i_8_)  &  (~ i_33_)  &  i_38_ ) ;
 assign _10216 = ( (~ i_28_)  &  (~ i_24_)  &  i_31_  &  i_34_ ) ;
 assign _10232 = ( wire7631 ) | ( _733 ) | ( (~ i_24_)  &  wire1100 ) ;
 assign _10281 = ( i_29_  &  (~ i_28_) ) ;
 assign _10282 = ( wire1086 ) | ( wire1087 ) | ( wire1081 ) | ( _702 ) ;
 assign _10283 = ( wire1070 ) | ( wire1080 ) | ( wire739  &  _10281 ) ;
 assign _10286 = ( i_38_  &  (~ i_35_) ) ;
 assign _10288 = ( (~ i_30_)  &  i_34_  &  (~ i_35_)  &  i_38_ ) ;
 assign _10290 = ( (~ i_32_)  &  (~ i_30_) ) ;
 assign _10292 = ( i_38_  &  (~ i_35_) ) ;
 assign _10294 = ( i_38_  &  (~ i_35_) ) ;
 assign _10313 = ( (~ i_7_)  &  (~ i_8_)  &  (~ i_24_)  &  (~ i_22_) ) ;
 assign _10317 = ( (~ i_30_)  &  (~ i_28_)  &  (~ i_32_) ) ;
 assign _10319 = ( i_12_  &  i_9_ ) ;
 assign _10324 = ( (~ i_12_)  &  (~ i_24_)  &  i_38_ ) ;
 assign _10326 = ( i_38_  &  (~ i_24_) ) ;
 assign _10331 = ( wire1045 ) | ( wire1044 ) ;
 assign _10332 = ( wire1041 ) | ( _674 ) | ( _676 ) | ( _677 ) ;
 assign _10341 = ( (~ i_2_)  &  (~ i_24_)  &  (~ i_22_) ) ;
 assign _10353 = ( wire1043 ) | ( wire1053 ) | ( wire1054 ) | ( wire7661 ) ;
 assign _10370 = ( (~ i_8_)  &  (~ i_7_) ) ;
 assign _10372 = ( (~ i_22_)  &  (~ i_7_) ) ;
 assign _10377 = ( (~ i_25_)  &  (~ i_26_)  &  (~ i_24_)  &  (~ i_31_) ) ;
 assign _10386 = ( (~ i_8_)  &  (~ i_25_)  &  (~ i_24_)  &  (~ i_31_) ) ;
 assign _10408 = ( wire999 ) | ( wire1023 ) | ( wire1024 ) | ( _637 ) ;
 assign _10409 = ( wire7705 ) | ( _655 ) | ( _656 ) ;
 assign _10425 = ( (~ i_26_)  &  (~ i_24_)  &  (~ i_22_) ) ;
 assign _10426 = ( (~ i_5_)  &  (~ i_4_)  &  (~ i_2_)  &  (~ i_32_) ) ;
 assign _10430 = ( (~ i_28_)  &  (~ i_32_)  &  (~ i_29_) ) ;
 assign _10432 = ( i_9_  &  i_12_  &  (~ i_24_)  &  i_38_ ) ;
 assign _10445 = ( (~ i_10_)  &  (~ i_24_)  &  (~ i_22_) ) ;
 assign _10448 = ( (~ i_30_)  &  (~ i_35_)  &  i_38_ ) ;
 assign _10457 = ( (~ i_7_)  &  (~ i_8_)  &  (~ i_5_)  &  (~ i_6_) ) ;
 assign _10458 = ( _606 ) | ( _612 ) | ( _613 ) ;
 assign _10460 = ( wire7502 ) | ( wire7503 ) | ( wire7504 ) | ( wire1064 ) ;
 assign _10465 = ( wire7274  &  wire404 ) ;
 assign _10469 = ( (~ i_9_)  &  (~ i_11_)  &  (~ i_19_) ) ;
 assign _10475 = ( (~ i_7_)  &  (~ i_5_)  &  (~ i_6_)  &  (~ i_18_) ) ;
 assign _10477 = ( (~ i_28_)  &  (~ i_32_)  &  (~ i_29_) ) ;
 assign _10478 = ( _595 ) | ( wire521  &  wire7446 ) | ( wire7446  &  _10465 ) ;
 assign _10480 = ( i_34_  &  (~ i_35_)  &  i_38_ ) ;
 assign _10484 = ( (~ i_28_)  &  i_38_  &  n_n1523  &  n_n1458 ) ;
 assign _10485 = ( (~ i_31_)  &  wire1289 ) | ( (~ i_31_)  &  wire4  &  _10484 ) ;
 assign _10491 = ( (~ i_2_)  &  (~ i_4_) ) ;
 assign _10496 = ( (~ i_24_)  &  (~ i_35_)  &  i_38_ ) ;
 assign _10498 = ( (~ i_6_)  &  (~ i_13_)  &  (~ i_12_)  &  i_18_ ) ;
 assign _10504 = ( wire434  &  wire430  &  _10496 ) | ( wire430  &  wire422  &  _10496 ) ;
 assign _10524 = ( (~ i_12_)  &  (~ i_6_) ) ;
 assign _10526 = ( n_n315  &  wire254 ) | ( n_n317  &  wire254 ) ;
 assign _10531 = ( (~ i_11_)  &  (~ i_19_)  &  wire429 ) ;
 assign _10533 = ( (~ i_24_)  &  wire446  &  wire78 ) ;
 assign _10534 = ( wire272  &  _10531 ) | ( wire4  &  _10533 ) ;
 assign _10536 = ( wire1240 ) | ( _585 ) | ( _10504 ) ;
 assign _10560 = ( (~ i_8_)  &  (~ i_31_)  &  (~ i_35_)  &  i_38_ ) ;
 assign _10575 = ( i_38_  &  (~ i_35_) ) ;
 assign _10578 = ( n_n1055  &  n_n461  &  wire7411 ) ;
 assign _10586 = ( i_10_  &  (~ i_13_)  &  i_12_  &  (~ i_22_) ) ;
 assign _10606 = ( n_n1055  &  n_n461  &  wire7411 ) | ( n_n461  &  wire7411  &  wire7412 ) ;
 assign _10607 = ( n_n1279  &  n_n819  &  wire7413 ) | ( n_n1279  &  n_n819  &  n_n735 ) ;
 assign _10625 = ( (~ i_24_)  &  (~ i_35_)  &  i_38_ ) ;
 assign _10626 = ( wire430  &  wire423  &  _10625 ) | ( wire430  &  wire435  &  _10625 ) ;
 assign _10628 = ( (~ i_33_)  &  (~ i_35_)  &  i_38_ ) ;
 assign _10631 = ( n_n1055  &  n_n461  &  wire7411 ) | ( n_n461  &  wire7411  &  wire7412 ) ;
 assign _10632 = ( n_n1279  &  n_n819  &  wire7413 ) | ( n_n1279  &  n_n819  &  n_n735 ) ;
 assign _10634 = ( wire1268 ) | ( wire1271 ) | ( _539 ) | ( _543 ) ;
 assign _10635 = ( n_n1847 ) | ( wire1274 ) | ( wire7458 ) | ( _10634 ) ;
 assign _10646 = ( (~ i_28_)  &  (~ i_33_)  &  (~ i_35_)  &  i_38_ ) ;
 assign _10648 = ( (~ i_10_)  &  (~ i_4_)  &  (~ i_1_)  &  (~ i_2_) ) ;
 assign _10651 = ( (~ i_10_)  &  (~ i_28_)  &  (~ i_25_)  &  (~ i_29_) ) ;
 assign _10658 = ( (~ i_25_)  &  (~ i_26_)  &  (~ i_24_) ) ;
 assign _10663 = ( (~ i_5_)  &  (~ i_4_)  &  (~ i_2_)  &  (~ i_31_) ) ;
 assign _10665 = ( (~ i_34_)  &  i_35_  &  i_38_ ) ;
 assign _10667 = ( (~ i_19_)  &  (~ i_11_) ) ;
 assign _10679 = ( (~ i_28_)  &  (~ i_33_)  &  (~ i_29_) ) ;
 assign _10690 = ( (~ i_10_)  &  (~ i_5_)  &  (~ i_4_)  &  (~ i_2_) ) ;
 assign _10693 = ( (~ i_5_)  &  (~ i_4_)  &  (~ i_2_)  &  (~ i_31_) ) ;
 assign _10705 = ( (~ i_32_)  &  (~ i_33_)  &  i_38_ ) ;
 assign _10708 = ( (~ i_6_)  &  (~ i_12_)  &  (~ i_24_) ) ;
 assign _10715 = ( (~ i_5_)  &  i_13_  &  (~ i_4_)  &  (~ i_2_) ) ;
 assign _10716 = ( (~ i_10_)  &  (~ i_5_)  &  (~ i_4_)  &  (~ i_2_) ) ;
 assign _10717 = ( (~ i_5_)  &  (~ i_4_)  &  (~ i_2_)  &  (~ i_32_) ) ;
 assign _10721 = ( (~ i_30_)  &  (~ i_2_)  &  (~ i_32_) ) ;
 assign _10722 = ( wire343  &  wire61 ) ;
 assign _10731 = ( i_9_  &  (~ i_10_)  &  (~ i_6_)  &  (~ i_12_) ) ;
 assign _10746 = ( (~ i_35_)  &  i_38_  &  (~ i_29_) ) ;
 assign _10748 = ( (~ i_25_)  &  (~ i_26_)  &  (~ i_24_) ) ;
 assign _10754 = ( (~ i_5_)  &  (~ i_4_)  &  (~ i_2_)  &  (~ i_32_) ) ;
 assign _10759 = ( n_n1852 ) | ( n_n1821 ) | ( wire7485 ) | ( _10635 ) ;
 assign _10762 = ( (~ i_10_)  &  (~ i_24_)  &  (~ i_22_) ) ;
 assign _10782 = ( (~ i_5_)  &  (~ i_4_)  &  (~ i_2_) ) ;
 assign _10785 = ( (~ i_35_)  &  i_38_  &  (~ i_29_) ) ;
 assign _10790 = ( wire1325 ) | ( wire7394 ) | ( wire7395 ) | ( _442 ) ;
 assign _10811 = ( n_n1523  &  wire434  &  _9998 ) | ( n_n1523  &  wire422  &  _9998 ) ;
 assign _10814 = ( wire1317 ) | ( wire1319 ) | ( _415 ) | ( _10811 ) ;
 assign _10816 = ( (~ i_24_)  &  (~ i_35_)  &  i_38_ ) ;
 assign _10819 = ( i_19_  &  wire78  &  _10816 ) ;
 assign _10822 = ( (~ i_28_)  &  (~ i_33_)  &  (~ i_35_)  &  i_38_ ) ;
 assign _10823 = ( (~ i_26_)  &  (~ i_24_)  &  (~ i_22_)  &  _10822 ) ;
 assign _10826 = ( n_n1055  &  n_n461  &  wire7411 ) | ( n_n461  &  wire7411  &  wire7412 ) ;
 assign _10827 = ( n_n1279  &  n_n819  &  wire7413 ) | ( n_n1279  &  n_n819  &  n_n735 ) ;
 assign _10828 = ( n_n1055  &  n_n461  &  wire7411 ) | ( n_n461  &  wire7411  &  wire7412 ) ;
 assign _10829 = ( n_n1279  &  n_n819  &  wire7413 ) | ( n_n1279  &  n_n819  &  n_n735 ) ;
 assign _10830 = ( wire1303 ) | ( _410 ) | ( wire657  &  _10819 ) ;
 assign _10831 = ( wire1305 ) | ( _400 ) | ( _401 ) | ( _402 ) ;
 assign _10833 = ( wire7432 ) | ( wire7433 ) | ( n_n1843 ) | ( _10814 ) ;
 assign _10846 = ( i_10_  &  (~ i_3_)  &  (~ i_33_)  &  i_38_ ) ;
 assign _10849 = ( (~ i_24_)  &  (~ i_22_)  &  i_38_  &  wire7265 ) ;
 assign _10850 = ( (~ i_11_)  &  (~ i_32_)  &  (~ i_19_) ) ;
 assign _10870 = ( (~ i_24_)  &  (~ i_22_)  &  i_38_ ) ;
 assign _10876 = ( (~ i_28_)  &  (~ i_24_)  &  (~ i_32_)  &  (~ i_29_) ) ;
 assign _10877 = ( (~ i_28_)  &  (~ i_24_)  &  (~ i_32_)  &  (~ i_29_) ) ;
 assign _10879 = ( (~ i_31_)  &  (~ i_35_)  &  i_38_ ) ;
 assign _10885 = ( (~ i_5_)  &  (~ i_4_)  &  (~ i_2_)  &  (~ i_31_) ) ;
 assign _10889 = ( (~ i_28_)  &  (~ i_25_)  &  (~ i_29_) ) ;
 assign _10917 = ( (~ i_24_)  &  wire446  &  wire71 ) ;
 assign _10918 = ( (~ i_30_)  &  (~ i_28_)  &  (~ i_32_)  &  wire7272 ) ;
 assign _10933 = ( (~ i_32_)  &  i_34_  &  (~ i_35_) ) ;
 assign _10937 = ( wire7311  &  (~ i_24_) ) ;
 assign _10942 = ( wire1419 ) | ( wire7312 ) | ( _335 ) | ( _336 ) ;
 assign _10948 = ( (~ i_5_)  &  (~ i_4_)  &  (~ i_2_)  &  (~ i_31_) ) ;
 assign _10950 = ( (~ i_28_)  &  (~ i_22_)  &  (~ i_35_)  &  i_38_ ) ;
 assign _10962 = ( (~ i_32_)  &  (~ i_35_)  &  i_38_ ) ;
 assign _10970 = ( n_n1854 ) | ( wire4  &  _10917 ) ;
 assign _10972 = ( n_n1829 ) | ( n_n1825 ) | ( wire1392 ) | ( wire7339 ) ;
 assign _10974 = ( wire7714 ) | ( n_n1831 ) | ( wire7598 ) | ( _10188 ) ;
 assign _10984 = ( wire232  &  wire44  &  wire7749 ) ;
 assign _10985 = ( (~ i_28_)  &  (~ i_23_)  &  (~ i_21_)  &  i_29_ ) ;
 assign _10990 = ( (~ i_35_)  &  i_36_ ) ;
 assign _10991 = ( n_n1443  &  n_n1369  &  _10985  &  _10990 ) ;
 assign _10994 = ( (~ i_13_)  &  (~ i_11_)  &  (~ i_16_)  &  n_n177 ) ;
 assign _10995 = ( (~ i_14_)  &  n_n1307  &  n_n1303  &  _9751 ) ;
 assign _10998 = ( (~ i_34_)  &  i_35_  &  n_n1258  &  n_n916 ) ;
 assign _10999 = ( wire7757  &  _10994 ) | ( wire272  &  _10998 ) ;
 assign _11001 = ( wire7751  &  _10984 ) | ( wire547  &  _10991 ) ;
 assign _11016 = ( wire420  &  wire455 ) | ( wire363  &  wire7763 ) ;
 assign _11020 = ( n_n787  &  n_n180  &  n_n179 ) ;
 assign _11021 = ( (~ i_13_)  &  n_n1307  &  n_n1303  &  _9684 ) ;
 assign _11023 = ( (~ i_34_)  &  i_35_  &  n_n301  &  n_n1258 ) ;
 assign _11024 = ( wire7766  &  _11020 ) | ( wire272  &  _11023 ) ;
 assign _11027 = ( (~ i_27_)  &  (~ i_28_)  &  (~ i_29_) ) ;
 assign _11029 = ( n_n1213  &  wire265  &  _11027 ) ;
 assign _11033 = ( (~ i_8_)  &  (~ i_14_)  &  (~ i_12_) ) ;
 assign _11037 = ( i_36_  &  n_n1375  &  n_n1400  &  n_n301 ) ;
 assign _11051 = ( wire7874 ) | ( wire7875 ) | ( _292 ) | ( _293 ) ;
 assign _11052 = ( (~ i_14_)  &  (~ i_23_)  &  (~ i_17_)  &  (~ i_16_) ) ;
 assign _11053 = ( _11052  &  wire80 ) ;
 assign _11055 = ( (~ i_5_)  &  (~ i_4_)  &  (~ i_2_)  &  (~ i_32_) ) ;
 assign _11056 = ( (~ i_9_)  &  (~ i_7_)  &  (~ i_6_)  &  _11055 ) ;
 assign _11063 = ( (~ i_32_)  &  i_36_  &  (~ i_35_) ) ;
 assign _11077 = ( (~ i_27_)  &  (~ i_28_)  &  i_31_ ) ;
 assign _11087 = ( i_36_  &  i_34_ ) ;
 assign _11089 = ( (~ i_13_)  &  n_n1307  &  n_n1303  &  _9684 ) ;
 assign _11093 = ( wire864 ) | ( wire850 ) | ( wire7881 ) | ( _11051 ) ;
 assign _11094 = ( i_36_  &  n_n1213  &  _11027 ) ;
 assign _11097 = ( (~ i_13_)  &  (~ i_31_)  &  i_36_  &  (~ i_35_) ) ;
 assign _11113 = ( (~ i_8_)  &  (~ i_14_)  &  (~ i_12_)  &  n_n1345 ) ;
 assign _11117 = ( (~ i_28_)  &  (~ i_32_)  &  (~ i_29_) ) ;
 assign _11118 = ( wire172 ) | ( wire79  &  n_n620  &  _11117 ) ;
 assign _11119 = ( wire176 ) | ( (~ i_13_)  &  (~ i_16_)  &  wire295 ) ;
 assign _11120 = ( wire8014 ) | ( _11118 ) | ( _11119 ) ;
 assign _11141 = ( (~ i_24_)  &  i_21_  &  (~ i_34_) ) ;
 assign _11146 = ( wire234 ) | ( wire304 ) | ( wire336 ) | ( _240 ) ;
 assign _11170 = ( (~ i_27_)  &  (~ i_28_)  &  i_36_  &  (~ i_29_) ) ;
 assign _11202 = ( (~ i_14_)  &  (~ i_31_)  &  i_36_  &  (~ i_35_) ) ;
 assign _11205 = ( wire166 ) | ( (~ i_14_)  &  (~ i_16_)  &  wire295 ) ;
 assign _11215 = ( (~ i_23_)  &  (~ i_24_)  &  (~ i_16_) ) ;
 assign _11227 = ( (~ i_8_)  &  (~ i_13_)  &  (~ i_12_)  &  n_n1345 ) ;
 assign _11262 = ( (~ i_27_)  &  (~ i_28_)  &  (~ i_26_) ) ;
 assign _11294 = ( n_n1578 ) | ( n_n1576 ) | ( wire174 ) | ( _11120 ) ;
 assign _11296 = ( (~ i_27_)  &  (~ i_28_)  &  (~ i_23_)  &  i_36_ ) ;
 assign _11307 = ( (~ i_27_)  &  (~ i_28_)  &  (~ i_29_) ) ;
 assign _11309 = ( (~ i_32_)  &  (~ i_31_)  &  (~ i_29_) ) ;
 assign _11313 = ( (~ i_35_)  &  i_36_ ) ;
 assign _11315 = ( n_n1307  &  n_n841  &  n_n301  &  _11313 ) ;
 assign _11325 = ( (~ i_27_)  &  (~ i_26_)  &  (~ i_24_) ) ;
 assign _11326 = ( n_n1429  &  wire307 ) | ( wire458  &  _11315 ) ;
 assign _11333 = ( (~ i_8_)  &  (~ i_12_)  &  n_n461  &  wire7820 ) ;
 assign _11334 = ( (~ i_35_)  &  i_36_ ) ;
 assign _11336 = ( n_n1307  &  n_n841  &  n_n916  &  _11334 ) ;
 assign _11343 = ( wire7819  &  _11333 ) | ( wire458  &  _11336 ) ;
 assign _11350 = ( (~ i_27_)  &  (~ i_28_)  &  (~ i_23_)  &  i_36_ ) ;
 assign _11354 = ( wire906 ) | ( wire7836 ) | ( wire7837 ) | ( _11343 ) ;
 assign _11360 = ( (~ i_13_)  &  (~ i_16_)  &  i_36_ ) ;
 assign _11361 = ( (~ i_27_)  &  (~ i_28_)  &  (~ i_32_)  &  (~ i_29_) ) ;
 assign _11362 = ( (~ i_14_)  &  (~ i_16_)  &  i_36_ ) ;
 assign _11363 = ( (~ i_28_)  &  (~ i_32_)  &  i_34_  &  (~ i_29_) ) ;
 assign _11365 = ( (~ i_5_)  &  (~ i_4_)  &  (~ i_2_)  &  (~ i_31_) ) ;
 assign _11366 = ( (~ i_8_)  &  (~ i_6_)  &  (~ i_12_)  &  _11365 ) ;
 assign _11372 = ( (~ i_27_)  &  (~ i_28_)  &  (~ i_24_)  &  i_21_ ) ;
 assign _11388 = ( wire7916 ) | ( wire7917 ) | ( wire7920 ) | ( wire7852 ) ;
 assign _11391 = ( (~ i_30_)  &  (~ i_32_)  &  (~ i_31_) ) ;
 assign _11393 = ( (~ i_24_)  &  (~ i_23_) ) ;
 assign _11395 = ( i_36_  &  (~ i_7_) ) ;
 assign _11400 = ( wire7926 ) | ( wire196 ) ;
 assign _11419 = ( i_33_  &  i_34_ ) ;
 assign _11422 = ( i_34_  &  i_31_ ) ;
 assign _11424 = ( i_34_  &  i_31_ ) ;
 assign _11425 = ( (~ i_28_)  &  i_25_  &  i_21_ ) ;
 assign _11428 = ( (~ i_28_)  &  i_0_  &  i_29_ ) ;
 assign _11430 = ( wire117 ) | ( _75 ) | ( _81 ) | ( _82 ) ;
 assign _11431 = ( _77 ) | ( _78 ) | ( _79 ) | ( _80 ) ;
 assign _11443 = ( (~ i_8_)  &  (~ i_7_) ) ;
 assign _11479 = ( i_33_  &  i_34_ ) ;
 assign _11482 = ( (~ i_13_)  &  (~ i_12_)  &  (~ i_16_) ) ;
 assign _11489 = ( wire918 ) | ( _41 ) | ( _42 ) ;
 assign _11495 = ( (~ i_24_)  &  i_21_  &  (~ i_34_) ) ;
 assign _11510 = ( (~ i_10_)  &  (~ i_13_)  &  (~ i_17_)  &  (~ i_16_) ) ;
 assign _11519 = ( wire232  &  wire44  &  wire7749 ) ;
 assign _11521 = ( (~ i_28_)  &  i_36_  &  (~ i_35_)  &  (~ i_29_) ) ;
 assign _11531 = ( (~ i_27_)  &  (~ i_28_)  &  (~ i_23_)  &  i_36_ ) ;
 assign _11532 = ( n_n1307  &  n_n1303  &  n_n130  &  _9781 ) ;
 assign _11544 = ( wire7771 ) | ( _294 ) | ( _303 ) | ( _11001 ) ;


endmodule

