module C7552 (
	P_4528_206_, P_4526_205_, P_4437_204_, P_4432_203_, P_4427_202_, P_4420_201_, P_4415_200_, P_4410_199_, 
	P_4405_198_, P_4400_197_, P_4394_196_, P_4393_195_, P_3749_194_, P_3743_193_, P_3737_192_, P_3729_191_, P_3723_190_, P_3717_189_, 
	P_3711_188_, P_3705_187_, P_3701_186_, P_3698_185_, P_2256_184_, P_2253_183_, P_2247_182_, P_2239_181_, P_2236_180_, P_2230_179_, 
	P_2224_178_, P_2218_177_, P_2211_176_, P_2208_175_, P_2204_174_, P_1496_173_, P_1492_172_, P_1486_171_, P_1480_170_, P_1469_169_, 
	P_1462_168_, P_1459_167_, P_1455_166_, P_1197_165_, P_339_164_, P_240_163_, P_239_162_, P_238_161_, P_237_160_, P_236_159_, 
	P_235_158_, P_234_157_, P_233_156_, P_232_155_, P_231_154_, P_230_153_, P_229_152_, P_228_151_, P_227_150_, P_226_149_, 
	P_225_148_, P_224_147_, P_223_146_, P_222_145_, P_221_144_, P_220_143_, P_219_142_, P_218_141_, P_217_140_, P_216_139_, 
	P_215_138_, P_214_137_, P_213_136_, P_212_135_, P_211_134_, P_210_133_, P_209_132_, P_208_131_, P_207_130_, P_206_129_, 
	P_205_128_, P_204_127_, P_203_126_, P_202_125_, P_201_124_, P_200_123_, P_199_122_, P_198_121_, P_197_120_, P_196_119_, 
	P_195_118_, P_194_117_, P_193_116_, P_192_115_, P_191_114_, P_190_113_, P_189_112_, P_188_111_, P_187_110_, P_186_109_, 
	P_185_108_, P_184_107_, P_183_106_, P_182_105_, P_181_104_, P_180_103_, P_179_102_, P_178_101_, P_177_100_, P_176_99_, 
	P_175_98_, P_174_97_, P_173_96_, P_172_95_, P_171_94_, P_170_93_, P_169_92_, P_168_91_, P_167_90_, P_166_89_, 
	P_165_88_, P_164_87_, P_163_86_, P_162_85_, P_161_84_, P_160_83_, P_159_82_, P_158_81_, P_157_80_, P_156_79_, 
	P_155_78_, P_154_77_, P_153_76_, P_152_75_, P_151_74_, P_150_73_, P_147_72_, P_144_71_, P_141_70_, P_138_69_, 
	P_135_68_, P_134_67_, P_133_66_, P_130_65_, P_127_64_, P_124_63_, P_121_62_, P_118_61_, P_115_60_, P_114_59_, 
	P_113_58_, P_112_57_, P_111_56_, P_110_55_, P_109_54_, P_106_53_, P_103_52_, P_100_51_, P_97_50_, P_94_49_, 
	P_89_48_, P_88_47_, P_87_46_, P_86_45_, P_85_44_, P_84_43_, P_83_42_, P_82_41_, P_81_40_, P_80_39_, 
	P_79_38_, P_78_37_, P_77_36_, P_76_35_, P_75_34_, P_74_33_, P_73_32_, P_70_31_, P_69_30_, P_66_29_, 
	P_65_28_, P_64_27_, P_63_26_, P_62_25_, P_61_24_, P_60_23_, P_59_22_, P_58_21_, P_57_20_, P_56_19_, 
	P_55_18_, P_54_17_, P_53_16_, P_50_15_, P_47_14_, P_44_13_, P_41_12_, P_38_11_, P_35_10_, P_32_9_, 
	P_29_8_, P_26_7_, P_23_6_, P_18_5_, P_15_4_, P_12_3_, P_9_2_, P_5_1_, P_1_0_, P_560_248_, 
	P_558_244_, P_556_242_, P_554_240_, P_552_238_, P_550_236_, P_548_234_, P_546_232_, P_544_230_, P_542_246_, P_540_227_, 
	P_538_224_, P_536_222_, P_534_220_, P_532_218_, P_530_216_, P_528_214_, P_526_212_, P_524_210_, P_522_226_, P_496_271_, 
	P_494_267_, P_492_265_, P_490_263_, P_488_260_, P_486_258_, P_484_256_, P_482_253_, P_480_250_, P_478_269_, P_471_3445_, 
	P_469_3452_, P_453_596_, P_450_288_, P_448_284_, P_446_393_, P_444_282_, P_442_280_, P_440_277_, P_438_274_, P_436_286_, 
	P_432_428_, P_422_3451_, P_419_3444_, P_418_3449_, P_416_3368_, P_414_3338_, P_412_3369_, P_410_387_, P_408_385_, P_406_388_, 
	P_404_390_, P_402_395_, P_399_3717_, P_397_3097_, P_394_3095_, P_391_3094_, P_388_3093_, P_385_3151_, P_382_3148_, P_379_3207_, 
	P_376_3206_, P_373_2994_, P_370_3718_, P_368_3431_, P_365_3430_, P_362_3429_, P_359_3426_, P_356_3424_, P_353_3425_, P_350_3421_, 
	P_347_3420_, P_344_3382_, P_341_420_, P_338_3716_, P_336_3412_, P_333_3416_, P_330_3411_, P_327_3408_, P_324_3363_, P_321_3715_, 
	P_319_3398_, P_316_3397_, P_313_3396_, P_310_3393_, P_307_3389_, P_304_3390_, P_301_3388_, P_298_3387_, P_295_3352_, P_292_392_, 
	P_289_383_, P_286_419_, P_284_384_, P_281_547_, P_279_304_, P_278_536_, P_276_3401_, P_273_3402_, P_270_3109_, P_264_3121_, 
	P_258_3122_, P_252_3450_, P_249_3418_, P_246_3110_, P_3_312_, P_2_313_);

input P_4528_206_, P_4526_205_, P_4437_204_, P_4432_203_, P_4427_202_, P_4420_201_, P_4415_200_, P_4410_199_, P_4405_198_, P_4400_197_, P_4394_196_, P_4393_195_, P_3749_194_, P_3743_193_, P_3737_192_, P_3729_191_, P_3723_190_, P_3717_189_, P_3711_188_, P_3705_187_, P_3701_186_, P_3698_185_, P_2256_184_, P_2253_183_, P_2247_182_, P_2239_181_, P_2236_180_, P_2230_179_, P_2224_178_, P_2218_177_, P_2211_176_, P_2208_175_, P_2204_174_, P_1496_173_, P_1492_172_, P_1486_171_, P_1480_170_, P_1469_169_, P_1462_168_, P_1459_167_, P_1455_166_, P_1197_165_, P_339_164_, P_240_163_, P_239_162_, P_238_161_, P_237_160_, P_236_159_, P_235_158_, P_234_157_, P_233_156_, P_232_155_, P_231_154_, P_230_153_, P_229_152_, P_228_151_, P_227_150_, P_226_149_, P_225_148_, P_224_147_, P_223_146_, P_222_145_, P_221_144_, P_220_143_, P_219_142_, P_218_141_, P_217_140_, P_216_139_, P_215_138_, P_214_137_, P_213_136_, P_212_135_, P_211_134_, P_210_133_, P_209_132_, P_208_131_, P_207_130_, P_206_129_, P_205_128_, P_204_127_, P_203_126_, P_202_125_, P_201_124_, P_200_123_, P_199_122_, P_198_121_, P_197_120_, P_196_119_, P_195_118_, P_194_117_, P_193_116_, P_192_115_, P_191_114_, P_190_113_, P_189_112_, P_188_111_, P_187_110_, P_186_109_, P_185_108_, P_184_107_, P_183_106_, P_182_105_, P_181_104_, P_180_103_, P_179_102_, P_178_101_, P_177_100_, P_176_99_, P_175_98_, P_174_97_, P_173_96_, P_172_95_, P_171_94_, P_170_93_, P_169_92_, P_168_91_, P_167_90_, P_166_89_, P_165_88_, P_164_87_, P_163_86_, P_162_85_, P_161_84_, P_160_83_, P_159_82_, P_158_81_, P_157_80_, P_156_79_, P_155_78_, P_154_77_, P_153_76_, P_152_75_, P_151_74_, P_150_73_, P_147_72_, P_144_71_, P_141_70_, P_138_69_, P_135_68_, P_134_67_, P_133_66_, P_130_65_, P_127_64_, P_124_63_, P_121_62_, P_118_61_, P_115_60_, P_114_59_, P_113_58_, P_112_57_, P_111_56_, P_110_55_, P_109_54_, P_106_53_, P_103_52_, P_100_51_, P_97_50_, P_94_49_, P_89_48_, P_88_47_, P_87_46_, P_86_45_, P_85_44_, P_84_43_, P_83_42_, P_82_41_, P_81_40_, P_80_39_, P_79_38_, P_78_37_, P_77_36_, P_76_35_, P_75_34_, P_74_33_, P_73_32_, P_70_31_, P_69_30_, P_66_29_, P_65_28_, P_64_27_, P_63_26_, P_62_25_, P_61_24_, P_60_23_, P_59_22_, P_58_21_, P_57_20_, P_56_19_, P_55_18_, P_54_17_, P_53_16_, P_50_15_, P_47_14_, P_44_13_, P_41_12_, P_38_11_, P_35_10_, P_32_9_, P_29_8_, P_26_7_, P_23_6_, P_18_5_, P_15_4_, P_12_3_, P_9_2_, P_5_1_, P_1_0_;

output P_560_248_, P_558_244_, P_556_242_, P_554_240_, P_552_238_, P_550_236_, P_548_234_, P_546_232_, P_544_230_, P_542_246_, P_540_227_, P_538_224_, P_536_222_, P_534_220_, P_532_218_, P_530_216_, P_528_214_, P_526_212_, P_524_210_, P_522_226_, P_496_271_, P_494_267_, P_492_265_, P_490_263_, P_488_260_, P_486_258_, P_484_256_, P_482_253_, P_480_250_, P_478_269_, P_471_3445_, P_469_3452_, P_453_596_, P_450_288_, P_448_284_, P_446_393_, P_444_282_, P_442_280_, P_440_277_, P_438_274_, P_436_286_, P_432_428_, P_422_3451_, P_419_3444_, P_418_3449_, P_416_3368_, P_414_3338_, P_412_3369_, P_410_387_, P_408_385_, P_406_388_, P_404_390_, P_402_395_, P_399_3717_, P_397_3097_, P_394_3095_, P_391_3094_, P_388_3093_, P_385_3151_, P_382_3148_, P_379_3207_, P_376_3206_, P_373_2994_, P_370_3718_, P_368_3431_, P_365_3430_, P_362_3429_, P_359_3426_, P_356_3424_, P_353_3425_, P_350_3421_, P_347_3420_, P_344_3382_, P_341_420_, P_338_3716_, P_336_3412_, P_333_3416_, P_330_3411_, P_327_3408_, P_324_3363_, P_321_3715_, P_319_3398_, P_316_3397_, P_313_3396_, P_310_3393_, P_307_3389_, P_304_3390_, P_301_3388_, P_298_3387_, P_295_3352_, P_292_392_, P_289_383_, P_286_419_, P_284_384_, P_281_547_, P_279_304_, P_278_536_, P_276_3401_, P_273_3402_, P_270_3109_, P_264_3121_, P_258_3122_, P_252_3450_, P_249_3418_, P_246_3110_, P_3_312_, P_2_313_;

wire wire43, wire93, wire101, n98, n99, n103, n106, n109, n112, n114, n116, n118, n122, n120, n123, n129, n130, n128, n126, n134, n133, n131, n138, n139, n137, n135, n143, n142, n140, n147, n145, n146, n144, n151, n152, n150, n148, n156, n153, n161, n159, n157, n165, n166, n164, n162, n170, n167, n174, n173, n171, n178, n175, n182, n179, n184, n185, n183, n187, n188, n186, n192, n193, n191, n189, n194, n196, n197, n198, n199, n195, n201, n202, n203, n204, n200, n206, n207, n208, n209, n205, n211, n212, n213, n214, n210, n215, n221, n222, n223, n224, n220, n226, n227, n228, n229, n225, n231, n232, n233, n234, n230, n236, n237, n238, n239, n235, n241, n242, n243, n244, n240, n246, n247, n248, n249, n245, n253, n251, n252, n250, n257, n256, n254, n261, n259, n260, n258, n265, n264, n262, n269, n267, n266, n273, n272, n270, n276, n277, n275, n274, n281, n282, n279, n278, n285, n286, n284, n283, n289, n290, n288, n287, n291, n292, n293, n294, n295, n296, n297, n298, n300, n301, n302, n303, n304, n305, n307, n312, n310, n311, n309, n313, n314, n315, n319, n317, n316, n322, n323, n320, n321, n327, n324, n325, n328, n329, n330, n331, n332, n336, n334, n340, n337, n341, n346, n343, n347, n349, n352, n354, n359, n356, n360, n362, n364, n369, n366, n370, n375, n372, n376, n381, n378, n382, n387, n384, n391, n388, n395, n392, n396, n400, n399, n403, n402, n408, n406, n405, n412, n410, n409, n416, n414, n413, n418, n417, n424, n422, n421, n426, n425, n432, n430, n429, n434, n433, n439, n437, n436, n441, n440, n445, n444, n449, n448, n452, n451, n453, n455, n457, n460, n462, n459, n463, n465, n467, n469, n471, n474, n476, n473, n477, n483, n479, n484, n486, n487, n485, n491, n492, n488, n493, n495, n496, n494, n498, n499, n500, n497, n504, n502, n503, n501, n506, n505, n507, n515, n513, n514, n512, n517, n526, n523, n524, n522, n532, n534, n531, n538, n536, n535, n542, n540, n539, n546, n544, n543, n547, n552, n551, n557, n554, n561, n559, n558, n563, n568, n567, n573, n571, n576, n577, n578, n580, n583, n581, n584, n586, n587, n589, n588, n593, n590, n595, n598, n600, n603, n606, n605, n607, n610, n609, n611, n613, n615, n616, n619, n620, n622, n621, n624, n623, n625, n626, n627, n629, n630, n628, n631, n633, n634, n632, n635, n636, n638, n639, n637, n640, n642, n641, n644, n643, n646, n645, n647, n649, n648, n650, n651, n652, n654, n655, n653, n657, n658, n656, n660, n659, n662, n661, n663, n667, n668, n671, n670, n673, n672, n676, n677, n679, n678, n681, n680, n683, n684, n686, n685, n689, n687, n690, n692, n693, n695, n696, n694, n697, n698, n699, n700, n703, n702, n706, n707, n710, n711, n712, n713, n715, n717, n718, n720, n722, n723, n724, n726, n728, n729, n730, n731, n732, n735, n734, n736, n737, n740, n739, n745, n746, n744, n750, n749, n751, n752, n753, n754, n755, n756, n757, n760, n762, n761, n763, n764, n765, n766, n767, n769, n770, n771, n772, n775, n776, n778, n779, n781, n783, n784, n785, n786, n789, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n808, n809, n807, n810, n811, n812, n813, n814, n815, n817, n818, n816, n819, n820, n821, n822, n823, n824, n826, n827, n825, n828, n830, n831, n829, n832, n834, n835, n833, n836, n838, n839, n837, n840, n842, n843, n841, n844, n846, n847, n845, n848, n850, n851, n849, n852, n853, n854, n855, n856, n857, n858, n859, n861, n863, n870, n872, n873, n874, n876, n877, n878, n880, n881, n882, n883, n884, n885, n886, n888, n889, n891, n892, n893, n895, n900, n901, n903, n904, n905, n906, n907, n908, n909, n910, n912, n913, n914, n915, n916, n918, n919, n917, n920, n921, n922, n923, n924, n925, n927, n928, n926, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n942, n943, n941, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n961, n962, n960, n963, n964, n966, n967, n968, n970, n971, n972, n976, n977, n978, n981, n984, n987, n988, n990, n991, n993, n994, n996, n997, n999, n1000, n1001, n1002, n1004, n1007, n1008, n1010, n1012, n1014, n1015, n1017, n1019, n1020, n1021, n1022, n1024, n1023, n1026, n1027, n1028, n1030, n1031, n1032, n1034, n1033, n1035, n1036, n1037, n1039, n1040, n1043, n1042, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1059, n1060, n1061, n1062, n1063, n1064, n1068, n1089;

assign P_469_3452_ = ( (~ n882) ) ;
 assign P_422_3451_ = ( (~ n882) ) ;
 assign wire43 = ( n590  &  n707 ) | ( (~ n590)  &  (~ n707) ) ;
 assign P_418_3449_ = ( P_416_3368_ ) | ( P_414_3338_ ) | ( P_412_3369_ ) | ( (~ n328) ) | ( (~ n329) ) | ( (~ n330) ) | ( (~ n331) ) ;
 assign P_416_3368_ = ( n300 ) | ( n301 ) | ( n302 ) | ( (~ n816) ) ;
 assign P_414_3338_ = ( n303 ) | ( n304 ) | ( n305 ) | ( (~ n807) ) ;
 assign P_412_3369_ = ( n295 ) | ( n296 ) | ( n297 ) | ( n298 ) ;
 assign P_410_387_ = ( (~ n331) ) ;
 assign P_408_385_ = ( (~ n330) ) ;
 assign P_406_388_ = ( (~ n329) ) ;
 assign P_404_390_ = ( (~ n328) ) ;
 assign P_402_395_ = ( P_57_20_ ) | ( P_5_1_ ) ;
 assign P_399_3717_ = ( n283  &  n1035 ) | ( (~ n283)  &  (~ n1035) ) ;
 assign P_397_3097_ = ( n448  &  n620 ) | ( (~ n448)  &  (~ n620) ) ;
 assign P_394_3095_ = ( n444  &  n619 ) | ( (~ n444)  &  (~ n619) ) ;
 assign P_391_3094_ = ( n186  &  n440 ) | ( (~ n186)  &  (~ n440) ) ;
 assign P_388_3093_ = ( n183  &  n436 ) | ( (~ n183)  &  (~ n436) ) ;
 assign P_385_3151_ = ( n194  &  n739 ) | ( (~ n194)  &  (~ n739) ) ;
 assign P_382_3148_ = ( (~ n873) ) ;
 assign P_379_3207_ = ( (~ n872) ) ;
 assign P_376_3206_ = ( n399  &  n623 ) | ( (~ n399)  &  (~ n623) ) ;
 assign P_373_2994_ = ( (~ P_4526_205_)  &  n702 ) | ( P_4526_205_  &  (~ n702) ) ;
 assign P_370_3718_ = ( n287  &  n1031 ) | ( (~ n287)  &  (~ n1031) ) ;
 assign P_368_3431_ = ( n433  &  n677 ) | ( (~ n433)  &  (~ n677) ) ;
 assign P_365_3430_ = ( n429  &  n676 ) | ( (~ n429)  &  (~ n676) ) ;
 assign P_362_3429_ = ( n270  &  n425 ) | ( (~ n270)  &  (~ n425) ) ;
 assign P_359_3426_ = ( n266  &  n421 ) | ( (~ n266)  &  (~ n421) ) ;
 assign P_356_3424_ = ( (~ n744)  &  n600 ) | ( n744  &  (~ n600) ) ;
 assign P_353_3425_ = ( (~ n881) ) ;
 assign P_350_3421_ = ( (~ n880) ) ;
 assign P_347_3420_ = ( n409  &  n680 ) | ( (~ n409)  &  (~ n680) ) ;
 assign P_344_3382_ = ( (~ n598)  &  n749 ) | ( n598  &  (~ n749) ) ;
 assign P_341_420_ = ( (~ P_15_4_) ) ;
 assign P_338_3716_ = ( n274  &  n1027 ) | ( (~ n274)  &  (~ n1027) ) ;
 assign P_336_3412_ = ( n349  &  n588 ) | ( (~ n349)  &  (~ n588) ) ;
 assign P_333_3416_ = ( n356  &  n587 ) | ( (~ n356)  &  (~ n587) ) ;
 assign P_330_3411_ = ( n262  &  n343 ) | ( (~ n262)  &  (~ n343) ) ;
 assign P_327_3408_ = ( n258  &  n337 ) | ( (~ n258)  &  (~ n337) ) ;
 assign P_324_3363_ = ( (~ n259)  &  n606 ) | ( n259  &  (~ n606) ) ;
 assign P_321_3715_ = ( n278  &  n1022 ) | ( (~ n278)  &  (~ n1022) ) ;
 assign P_319_3398_ = ( n396  &  n668 ) | ( (~ n396)  &  (~ n668) ) ;
 assign P_316_3397_ = ( n392  &  n667 ) | ( (~ n392)  &  (~ n667) ) ;
 assign P_313_3396_ = ( n254  &  n388 ) | ( (~ n254)  &  (~ n388) ) ;
 assign P_310_3393_ = ( n250  &  n384 ) | ( (~ n250)  &  (~ n384) ) ;
 assign P_307_3389_ = ( n173  &  n595 ) | ( (~ n173)  &  (~ n595) ) ;
 assign P_304_3390_ = ( (~ n877) ) ;
 assign P_301_3388_ = ( (~ n876) ) ;
 assign P_298_3387_ = ( n366  &  n672 ) | ( (~ n366)  &  (~ n672) ) ;
 assign P_295_3352_ = ( n251  &  n734 ) | ( (~ n251)  &  (~ n734) ) ;
 assign P_292_392_ = ( (~ n332) ) ;
 assign P_286_419_ = ( (~ P_15_4_) ) ;
 assign wire93 = ( (~ P_1197_165_) ) | ( P_5_1_ ) ;
 assign P_281_547_ = ( (~ n332) ) ;
 assign P_279_304_ = ( (~ P_15_4_) ) ;
 assign P_278_536_ = ( P_163_86_  &  P_1_0_ ) ;
 assign P_276_3401_ = ( (~ n120) ) | ( n613 ) ;
 assign P_273_3402_ = ( (~ n294) ) ;
 assign P_270_3109_ = ( (~ n307) ) ;
 assign wire101 = ( n292 ) | ( n293 ) ;
 assign P_252_3450_ = ( (~ n291) ) ;
 assign P_246_3110_ = ( (~ n307) ) ;
 assign n98 = ( P_12_3_  &  P_9_2_ ) ;
 assign n99 = ( (~ P_180_103_)  &  (~ n1050) ) | ( (~ P_18_5_)  &  (~ n1050) ) ;
 assign n103 = ( (~ P_179_102_)  &  (~ n1049) ) | ( (~ P_18_5_)  &  (~ n1049) ) ;
 assign n106 = ( (~ P_178_101_)  &  (~ n1051) ) | ( (~ P_18_5_)  &  (~ n1051) ) ;
 assign n109 = ( (~ P_171_94_)  &  (~ n1048) ) | ( (~ P_18_5_)  &  (~ n1048) ) ;
 assign n112 = ( (~ P_160_83_)  &  (~ n1050) ) | ( (~ P_18_5_)  &  (~ n1050) ) ;
 assign n114 = ( (~ P_159_82_)  &  (~ n1049) ) | ( (~ P_18_5_)  &  (~ n1049) ) ;
 assign n116 = ( (~ P_158_81_)  &  (~ n1051) ) | ( (~ P_18_5_)  &  (~ n1051) ) ;
 assign n118 = ( (~ P_151_74_)  &  (~ n1048) ) | ( (~ P_18_5_)  &  (~ n1048) ) ;
 assign n122 = ( (~ P_38_11_) ) | ( (~ n706) ) ;
 assign n120 = ( P_1496_173_  &  n122 ) | ( (~ P_38_11_)  &  n122 ) ;
 assign n123 = ( (~ n707)  &  (~ n854) ) ;
 assign n129 = ( (~ n384) ) | ( n391  &  n728 ) ;
 assign n130 = ( n387  &  (~ n384) ) | ( n387  &  n731 ) ;
 assign n128 = ( (~ n388) ) | ( n729 ) ;
 assign n126 = ( n129  &  n130  &  n128 ) | ( n129  &  n130  &  (~ n384) ) ;
 assign n134 = ( n112 ) | ( P_2218_177_ ) ;
 assign n133 = ( n118 ) | ( P_2211_176_ ) ;
 assign n131 = ( n134  &  n133 ) | ( n134  &  (~ n396) ) ;
 assign n138 = ( (~ n337) ) | ( n346  &  n711 ) ;
 assign n139 = ( n340  &  (~ n337) ) | ( n340  &  n713 ) ;
 assign n137 = ( (~ n343) ) | ( n712 ) ;
 assign n135 = ( n138  &  n139  &  n137 ) | ( n138  &  n139  &  (~ n337) ) ;
 assign n143 = ( P_1469_169_ ) | ( n347 ) ;
 assign n142 = ( P_1462_168_ ) | ( n352 ) ;
 assign n140 = ( n143  &  n142 ) | ( n143  &  (~ n349) ) ;
 assign n147 = ( n322  &  n323  &  n320 ) | ( n322  &  n323  &  n321 ) ;
 assign n145 = ( (~ P_3729_191_)  &  P_53_16_ ) | ( (~ P_3729_191_)  &  P_18_5_ ) | ( P_53_16_  &  (~ P_18_5_) ) ;
 assign n146 = ( P_203_126_  &  P_130_65_ ) | ( P_203_126_  &  P_18_5_ ) | ( P_130_65_  &  (~ P_18_5_) ) ;
 assign n144 = ( n147  &  n145 ) | ( n147  &  n146 ) ;
 assign n151 = ( (~ n421) ) | ( (~ n779)  &  n781 ) ;
 assign n152 = ( n424  &  (~ n421) ) | ( n424  &  n786 ) ;
 assign n150 = ( (~ n425) ) | ( n783 ) ;
 assign n148 = ( n151  &  n152  &  n150 ) | ( n151  &  n152  &  (~ n421) ) ;
 assign n156 = ( P_4400_197_ ) | ( (~ n434) ) ;
 assign n153 = ( n156  &  (~ n433) ) | ( n156  &  (~ n784) ) ;
 assign n161 = ( (~ n399) ) | ( n760  &  n764 ) ;
 assign n159 = ( P_3743_193_ ) | ( (~ n403) ) ;
 assign n157 = ( n161  &  n159  &  (~ n1052) ) | ( n161  &  (~ n399)  &  (~ n1052) ) ;
 assign n165 = ( (~ n436) ) | ( (~ n765)  &  n767 ) ;
 assign n166 = ( n439  &  (~ n436) ) | ( n439  &  n772 ) ;
 assign n164 = ( (~ n440) ) | ( n769 ) ;
 assign n162 = ( n165  &  n166  &  n164 ) | ( n165  &  n166  &  (~ n436) ) ;
 assign n170 = ( P_3705_187_ ) | ( (~ n449) ) ;
 assign n167 = ( n170  &  (~ n448) ) | ( n170  &  (~ n770) ) ;
 assign n174 = ( n381  &  n723 ) ;
 assign n173 = ( (~ n722) ) | ( n726 ) ;
 assign n171 = ( n174  &  n173 ) | ( n174  &  (~ n378) ) ;
 assign n178 = ( (~ n775)  &  n778 ) ;
 assign n175 = ( n178  &  (~ n417) ) | ( n178  &  (~ n744) ) ;
 assign n182 = ( n408  &  n763 ) ;
 assign n179 = ( n182  &  (~ n405) ) | ( n182  &  (~ n739) ) ;
 assign n184 = ( n164  &  (~ n765)  &  n767  &  n772 ) ;
 assign n185 = ( n188 ) | ( (~ n440) ) ;
 assign n183 = ( n184  &  n185 ) ;
 assign n187 = ( (~ n766)  &  n769  &  n771 ) ;
 assign n188 = ( (~ n444) ) | ( n793 ) ;
 assign n186 = ( n187  &  n188 ) ;
 assign n192 = ( n148 ) | ( (~ n409) ) | ( n753 ) ;
 assign n193 = ( n412  &  (~ n409)  &  n883 ) | ( n412  &  n776  &  n883 ) ;
 assign n191 = ( (~ n413) ) | ( n778 ) ;
 assign n189 = ( n192  &  n193  &  n191 ) | ( n192  &  n193  &  (~ n409) ) ;
 assign n194 = ( n162  &  n185 ) | ( n162  &  (~ n436) ) ;
 assign n196 = ( (~ n647) ) | ( (~ n648) ) | ( n1000 ) ;
 assign n197 = ( n647 ) | ( (~ n648) ) | ( (~ n1000) ) ;
 assign n198 = ( (~ n647) ) | ( n648 ) | ( (~ n1000) ) ;
 assign n199 = ( n647 ) | ( n648 ) | ( n1000 ) ;
 assign n195 = ( n196  &  n197  &  n198  &  n199 ) ;
 assign n201 = ( (~ n643) ) | ( (~ n645) ) | ( n997 ) ;
 assign n202 = ( n643 ) | ( (~ n645) ) | ( (~ n997) ) ;
 assign n203 = ( (~ n643) ) | ( n645 ) | ( (~ n997) ) ;
 assign n204 = ( n643 ) | ( n645 ) | ( n997 ) ;
 assign n200 = ( n201  &  n202  &  n203  &  n204 ) ;
 assign n206 = ( (~ n663) ) | ( n1015 ) | ( n1040 ) ;
 assign n207 = ( (~ n663) ) | ( (~ n1015) ) | ( (~ n1040) ) ;
 assign n208 = ( n663 ) | ( (~ n1015) ) | ( n1040 ) ;
 assign n209 = ( n663 ) | ( n1015 ) | ( (~ n1040) ) ;
 assign n205 = ( n206  &  n207  &  n208  &  n209 ) ;
 assign n211 = ( (~ n636) ) | ( n988 ) | ( (~ n1037) ) ;
 assign n212 = ( (~ n636) ) | ( (~ n988) ) | ( n1037 ) ;
 assign n213 = ( n636 ) | ( (~ n988) ) | ( (~ n1037) ) ;
 assign n214 = ( n636 ) | ( n1037 ) | ( n988 ) ;
 assign n210 = ( n211  &  n212  &  n213  &  n214 ) ;
 assign n215 = ( (~ n157)  &  (~ n451)  &  (~ n755) ) | ( (~ n162)  &  (~ n451)  &  (~ n755) ) ;
 assign n221 = ( (~ n632) ) | ( (~ n635) ) | ( (~ n984) ) ;
 assign n222 = ( n632 ) | ( (~ n635) ) | ( n984 ) ;
 assign n223 = ( (~ n632) ) | ( n635 ) | ( n984 ) ;
 assign n224 = ( n632 ) | ( n635 ) | ( (~ n984) ) ;
 assign n220 = ( n221  &  n222  &  n223  &  n224 ) ;
 assign n226 = ( (~ n659) ) | ( (~ n661) ) | ( n1012 ) ;
 assign n227 = ( n659 ) | ( (~ n661) ) | ( (~ n1012) ) ;
 assign n228 = ( (~ n659) ) | ( n661 ) | ( (~ n1012) ) ;
 assign n229 = ( n659 ) | ( n661 ) | ( n1012 ) ;
 assign n225 = ( n226  &  n227  &  n228  &  n229 ) ;
 assign n231 = ( (~ n628) ) | ( (~ n631) ) | ( (~ n981) ) ;
 assign n232 = ( n628 ) | ( (~ n631) ) | ( n981 ) ;
 assign n233 = ( (~ n628) ) | ( n631 ) | ( n981 ) ;
 assign n234 = ( n628 ) | ( n631 ) | ( (~ n981) ) ;
 assign n230 = ( n231  &  n232  &  n233  &  n234 ) ;
 assign n236 = ( (~ n640) ) | ( (~ n641) ) | ( n994 ) ;
 assign n237 = ( n640 ) | ( (~ n641) ) | ( (~ n994) ) ;
 assign n238 = ( (~ n640) ) | ( n641 ) | ( (~ n994) ) ;
 assign n239 = ( n640 ) | ( n641 ) | ( n994 ) ;
 assign n235 = ( n236  &  n237  &  n238  &  n239 ) ;
 assign n241 = ( (~ n637) ) | ( n991 ) | ( n1039 ) ;
 assign n242 = ( (~ n637) ) | ( (~ n991) ) | ( (~ n1039) ) ;
 assign n243 = ( n637 ) | ( n991 ) | ( (~ n1039) ) ;
 assign n244 = ( n637 ) | ( (~ n991) ) | ( n1039 ) ;
 assign n240 = ( n241  &  n242  &  n243  &  n244 ) ;
 assign n246 = ( (~ n653) ) | ( (~ n656) ) | ( n1010 ) ;
 assign n247 = ( n653 ) | ( (~ n656) ) | ( (~ n1010) ) ;
 assign n248 = ( (~ n653) ) | ( n656 ) | ( (~ n1010) ) ;
 assign n249 = ( n653 ) | ( n656 ) | ( n1010 ) ;
 assign n245 = ( n246  &  n247  &  n248  &  n249 ) ;
 assign n253 = ( n128  &  n731  &  n391  &  n728 ) ;
 assign n251 = ( n189  &  (~ n215)  &  n756 ) ;
 assign n252 = ( (~ n388) ) | ( n736 ) ;
 assign n250 = ( n253  &  n251 ) | ( n253  &  n252 ) ;
 assign n257 = ( n395  &  n729  &  n730 ) ;
 assign n256 = ( (~ n396) ) | ( n794 ) ;
 assign n254 = ( n257  &  n256 ) | ( n257  &  (~ n392) ) ;
 assign n261 = ( n137  &  n713  &  n346  &  n711 ) ;
 assign n259 = ( n313  &  n314  &  n315 ) ;
 assign n260 = ( (~ n343) ) | ( n717 ) ;
 assign n258 = ( n261  &  n259 ) | ( n261  &  n260 ) ;
 assign n265 = ( n359  &  n710  &  n712 ) ;
 assign n264 = ( (~ n349) ) | ( n589 ) ;
 assign n262 = ( n265  &  n264 ) | ( n265  &  (~ n356) ) ;
 assign n269 = ( n150  &  (~ n779)  &  n781  &  n786 ) ;
 assign n267 = ( (~ n425) ) | ( n751 ) ;
 assign n266 = ( n269  &  n267 ) | ( n269  &  (~ n598) ) ;
 assign n273 = ( n432  &  n783  &  n785 ) ;
 assign n272 = ( (~ n433) ) | ( n795 ) ;
 assign n270 = ( n273  &  n272 ) | ( n273  &  (~ n429) ) ;
 assign n276 = ( (~ n135) ) | ( (~ n259) ) | ( n1042 ) ;
 assign n277 = ( n259  &  n1026 ) | ( n275  &  n1026 ) | ( (~ n593)  &  n1026 ) ;
 assign n275 = ( (~ n854)  &  n1024 ) | ( n707  &  n1024  &  n1023 ) ;
 assign n274 = ( n276  &  n277  &  n135 ) | ( n276  &  n277  &  n275 ) ;
 assign n281 = ( n251 ) | ( n685 ) | ( n1021 ) ;
 assign n282 = ( n1020  &  n126 ) | ( n1020  &  n685 ) ;
 assign n279 = ( (~ n683)  &  n684 ) | ( n683  &  (~ n684) ) ;
 assign n278 = ( n281  &  n282  &  n279 ) | ( n281  &  n282  &  (~ n1021) ) ;
 assign n285 = ( P_4526_205_ ) | ( (~ n162) ) | ( n694 ) ;
 assign n286 = ( (~ P_4526_205_)  &  n1032 ) | ( n284  &  n1032 ) | ( n609  &  n1032 ) ;
 assign n284 = ( (~ n697)  &  n698 ) | ( n697  &  (~ n698) ) ;
 assign n283 = ( n285  &  n286  &  n162 ) | ( n285  &  n286  &  n284 ) ;
 assign n289 = ( (~ n148) ) | ( n687 ) | ( n796 ) ;
 assign n290 = ( n288  &  n1030 ) | ( (~ n796)  &  n1030 ) | ( n1028  &  n1030 ) ;
 assign n288 = ( (~ n692)  &  n693 ) | ( n692  &  (~ n693) ) ;
 assign n287 = ( n289  &  n290  &  n148 ) | ( n289  &  n290  &  n288 ) ;
 assign n291 = ( (~ n522)  &  (~ n856)  &  (~ n1061) ) | ( (~ n522)  &  (~ n857)  &  (~ n1061) ) ;
 assign n292 = ( (~ P_4528_206_)  &  n576 ) | ( P_2204_174_  &  n576 ) | ( P_38_11_  &  n576 ) ;
 assign n293 = ( (~ P_4528_206_)  &  P_38_11_ ) | ( P_2204_174_  &  P_38_11_ ) | ( P_1455_166_  &  P_38_11_ ) ;
 assign n294 = ( n120  &  (~ n123) ) | ( n120  &  (~ n590) ) ;
 assign n295 = ( (~ n801)  &  n802 ) | ( n801  &  (~ n802) ) ;
 assign n296 = ( (~ n803)  &  n804 ) | ( n803  &  (~ n804) ) ;
 assign n297 = ( (~ n580)  &  n627 ) | ( n580  &  (~ n627) ) ;
 assign n298 = ( (~ n799)  &  n800 ) | ( n799  &  (~ n800) ) ;
 assign n300 = ( (~ n819)  &  n820 ) | ( n819  &  (~ n820) ) ;
 assign n301 = ( (~ n586)  &  n652 ) | ( n586  &  (~ n652) ) ;
 assign n302 = ( (~ n814)  &  n815 ) | ( n814  &  (~ n815) ) ;
 assign n303 = ( (~ n810)  &  n811 ) | ( n810  &  (~ n811) ) ;
 assign n304 = ( (~ n812)  &  n813 ) | ( n812  &  (~ n813) ) ;
 assign n305 = ( (~ n805)  &  n806 ) | ( n805  &  (~ n806) ) ;
 assign n307 = ( n360  &  n259 ) | ( n360  &  n577 ) ;
 assign n312 = ( n327  &  n324  &  (~ n888) ) | ( n327  &  n325  &  (~ n888) ) ;
 assign n310 = ( (~ P_3705_187_)  &  P_74_33_ ) | ( (~ P_3705_187_)  &  P_18_5_ ) | ( P_74_33_  &  (~ P_18_5_) ) ;
 assign n311 = ( P_207_130_  &  P_29_8_ ) | ( P_207_130_  &  P_18_5_ ) | ( P_29_8_  &  (~ P_18_5_) ) ;
 assign n309 = ( n312  &  n310 ) | ( n312  &  n311 ) ;
 assign n313 = ( n757 ) | ( n189  &  (~ n215) ) ;
 assign n314 = ( n126  &  n885 ) | ( (~ n366)  &  n885 ) | ( n732  &  n885 ) ;
 assign n315 = ( n369  &  (~ n366)  &  n884 ) | ( n369  &  n375  &  n884 ) ;
 assign n319 = ( (~ n467) ) | ( n855 ) ;
 assign n317 = ( (~ P_2253_183_)  &  P_109_54_ ) | ( (~ P_2253_183_)  &  P_18_5_ ) | ( P_109_54_  &  (~ P_18_5_) ) ;
 assign n316 = ( n319  &  n317 ) | ( n319  &  (~ n465) ) ;
 assign n322 = ( n487 ) | ( n486 ) ;
 assign n323 = ( n863 ) | ( n861 ) ;
 assign n320 = ( (~ P_3737_192_)  &  P_54_17_ ) | ( (~ P_3737_192_)  &  P_18_5_ ) | ( P_54_17_  &  (~ P_18_5_) ) ;
 assign n321 = ( P_202_125_  &  P_127_64_ ) | ( P_202_125_  &  P_18_5_ ) | ( P_127_64_  &  (~ P_18_5_) ) ;
 assign n327 = ( n639 ) | ( n658 ) ;
 assign n324 = ( (~ P_3711_188_)  &  P_76_35_ ) | ( (~ P_3711_188_)  &  P_18_5_ ) | ( P_76_35_  &  (~ P_18_5_) ) ;
 assign n325 = ( P_206_129_  &  P_26_7_ ) | ( P_206_129_  &  P_18_5_ ) | ( P_26_7_  &  (~ P_18_5_) ) ;
 assign n328 = ( P_150_73_  &  P_184_107_  &  P_228_151_  &  P_240_163_ ) ;
 assign n329 = ( P_210_133_  &  P_152_75_  &  P_218_141_  &  P_230_153_ ) ;
 assign n330 = ( P_183_106_  &  P_182_105_  &  P_185_108_  &  P_186_109_ ) ;
 assign n331 = ( P_162_85_  &  P_172_95_  &  P_188_111_  &  P_199_122_ ) ;
 assign n332 = ( P_134_67_  &  P_133_66_  &  (~ P_5_1_) ) ;
 assign n336 = ( n98 ) | ( P_18_5_ ) ;
 assign n334 = ( (~ P_213_136_)  &  n336 ) | ( n98  &  n336 ) ;
 assign n340 = ( P_1486_171_ ) | ( n334 ) ;
 assign n337 = ( (~ P_1486_171_)  &  n340 ) | ( (~ n334)  &  n340 ) ;
 assign n341 = ( (~ P_214_137_)  &  n336 ) | ( n98  &  n336 ) ;
 assign n346 = ( P_1480_170_ ) | ( n341 ) ;
 assign n343 = ( (~ P_1480_170_)  &  n346 ) | ( (~ n341)  &  n346 ) ;
 assign n347 = ( (~ P_216_139_)  &  n336 ) | ( n98  &  n336 ) ;
 assign n349 = ( (~ P_1469_169_)  &  n143 ) | ( n143  &  (~ n347) ) ;
 assign n352 = ( (~ P_209_132_)  &  n336 ) | ( n98  &  n336 ) ;
 assign n354 = ( (~ P_215_138_)  &  n336 ) | ( n98  &  n336 ) ;
 assign n359 = ( P_106_53_ ) | ( n354 ) ;
 assign n356 = ( (~ P_106_53_)  &  n359 ) | ( (~ n354)  &  n359 ) ;
 assign n360 = ( n120  &  (~ n123) ) | ( n120  &  n135 ) ;
 assign n362 = ( (~ P_153_76_)  &  n336 ) | ( n98  &  n336 ) ;
 assign n364 = ( (~ P_154_77_)  &  n336 ) | ( n98  &  n336 ) ;
 assign n369 = ( P_2256_184_ ) | ( n362 ) ;
 assign n366 = ( (~ P_2256_184_)  &  n369 ) | ( (~ n362)  &  n369 ) ;
 assign n370 = ( (~ P_155_78_)  &  n336 ) | ( n98  &  n336 ) ;
 assign n375 = ( P_2253_183_ ) | ( n364 ) ;
 assign n372 = ( (~ P_2253_183_)  &  n375 ) | ( (~ n364)  &  n375 ) ;
 assign n376 = ( (~ P_156_79_)  &  n336 ) | ( n98  &  n336 ) ;
 assign n381 = ( P_2247_182_ ) | ( n370 ) ;
 assign n378 = ( (~ P_2247_182_)  &  n381 ) | ( (~ n370)  &  n381 ) ;
 assign n382 = ( (~ P_157_80_)  &  n336 ) | ( n98  &  n336 ) ;
 assign n387 = ( P_2236_180_ ) | ( n382 ) ;
 assign n384 = ( (~ P_2236_180_)  &  n387 ) | ( (~ n382)  &  n387 ) ;
 assign n391 = ( n116 ) | ( P_2230_179_ ) ;
 assign n388 = ( (~ P_2230_179_)  &  n391 ) | ( (~ n116)  &  n391 ) ;
 assign n395 = ( n114 ) | ( P_2224_178_ ) ;
 assign n392 = ( (~ P_2224_178_)  &  n395 ) | ( (~ n114)  &  n395 ) ;
 assign n396 = ( (~ P_2218_177_)  &  n134 ) | ( (~ n112)  &  n134 ) ;
 assign n400 = ( P_231_154_  &  P_100_51_ ) | ( P_231_154_  &  P_18_5_ ) | ( P_100_51_  &  (~ P_18_5_) ) ;
 assign n399 = ( (~ P_3749_194_)  &  (~ n1052) ) | ( n400  &  (~ n1052) ) ;
 assign n403 = ( P_232_155_  &  P_124_63_ ) | ( P_232_155_  &  P_18_5_ ) | ( P_124_63_  &  (~ P_18_5_) ) ;
 assign n402 = ( (~ P_3743_193_)  &  n159 ) | ( n159  &  n403 ) ;
 assign n408 = ( P_3737_192_ ) | ( (~ n406) ) ;
 assign n406 = ( P_233_156_  &  P_127_64_ ) | ( P_233_156_  &  P_18_5_ ) | ( P_127_64_  &  (~ P_18_5_) ) ;
 assign n405 = ( (~ P_3737_192_)  &  n408 ) | ( n408  &  n406 ) ;
 assign n412 = ( P_4437_204_ ) | ( (~ n410) ) ;
 assign n410 = ( P_219_142_  &  P_66_29_ ) | ( P_219_142_  &  P_18_5_ ) | ( P_66_29_  &  (~ P_18_5_) ) ;
 assign n409 = ( (~ P_4437_204_)  &  n412 ) | ( n412  &  n410 ) ;
 assign n416 = ( P_4432_203_ ) | ( (~ n414) ) ;
 assign n414 = ( P_220_143_  &  P_50_15_ ) | ( P_220_143_  &  P_18_5_ ) | ( P_50_15_  &  (~ P_18_5_) ) ;
 assign n413 = ( (~ P_4432_203_)  &  n416 ) | ( n416  &  n414 ) ;
 assign n418 = ( P_221_144_  &  P_32_9_ ) | ( P_221_144_  &  P_18_5_ ) | ( P_32_9_  &  (~ P_18_5_) ) ;
 assign n417 = ( (~ P_4427_202_)  &  (~ n775) ) | ( n418  &  (~ n775) ) ;
 assign n424 = ( P_4415_200_ ) | ( (~ n422) ) ;
 assign n422 = ( P_223_146_  &  P_47_14_ ) | ( P_223_146_  &  P_18_5_ ) | ( P_47_14_  &  (~ P_18_5_) ) ;
 assign n421 = ( (~ P_4415_200_)  &  n424 ) | ( n424  &  n422 ) ;
 assign n426 = ( P_224_147_  &  P_121_62_ ) | ( P_224_147_  &  P_18_5_ ) | ( P_121_62_  &  (~ P_18_5_) ) ;
 assign n425 = ( (~ P_4410_199_)  &  (~ n779) ) | ( n426  &  (~ n779) ) ;
 assign n432 = ( P_4405_198_ ) | ( (~ n430) ) ;
 assign n430 = ( P_225_148_  &  P_94_49_ ) | ( P_225_148_  &  P_18_5_ ) | ( P_94_49_  &  (~ P_18_5_) ) ;
 assign n429 = ( (~ P_4405_198_)  &  n432 ) | ( n432  &  n430 ) ;
 assign n434 = ( P_226_149_  &  P_97_50_ ) | ( P_226_149_  &  P_18_5_ ) | ( P_97_50_  &  (~ P_18_5_) ) ;
 assign n433 = ( (~ P_4400_197_)  &  n156 ) | ( n156  &  n434 ) ;
 assign n439 = ( P_3723_190_ ) | ( (~ n437) ) ;
 assign n437 = ( P_235_158_  &  P_103_52_ ) | ( P_235_158_  &  P_18_5_ ) | ( P_103_52_  &  (~ P_18_5_) ) ;
 assign n436 = ( (~ P_3723_190_)  &  n439 ) | ( n439  &  n437 ) ;
 assign n441 = ( P_236_159_  &  P_23_6_ ) | ( P_236_159_  &  P_18_5_ ) | ( P_23_6_  &  (~ P_18_5_) ) ;
 assign n440 = ( (~ P_3717_189_)  &  (~ n765) ) | ( n441  &  (~ n765) ) ;
 assign n445 = ( P_237_160_  &  P_26_7_ ) | ( P_237_160_  &  P_18_5_ ) | ( P_26_7_  &  (~ P_18_5_) ) ;
 assign n444 = ( (~ P_3711_188_)  &  (~ n766) ) | ( n445  &  (~ n766) ) ;
 assign n449 = ( P_238_161_  &  P_29_8_ ) | ( P_238_161_  &  P_18_5_ ) | ( P_29_8_  &  (~ P_18_5_) ) ;
 assign n448 = ( (~ P_3705_187_)  &  n170 ) | ( n170  &  n449 ) ;
 assign n452 = ( (~ n402) ) | ( (~ n405) ) | ( (~ n739) ) ;
 assign n451 = ( n157  &  (~ n399) ) | ( n157  &  n452 ) ;
 assign n453 = ( (~ P_166_89_)  &  n336 ) | ( n98  &  n336 ) ;
 assign n455 = ( (~ P_167_90_)  &  n336 ) | ( n98  &  n336 ) ;
 assign n457 = ( (~ P_168_91_)  &  n336 ) | ( n98  &  n336 ) ;
 assign n460 = ( (~ n455) ) | ( n568 ) ;
 assign n462 = ( (~ P_106_53_)  &  P_87_46_ ) | ( (~ P_106_53_)  &  P_18_5_ ) | ( P_87_46_  &  (~ P_18_5_) ) ;
 assign n459 = ( (~ n457)  &  n460  &  n462 ) ;
 assign n463 = ( (~ P_169_92_)  &  n336 ) | ( n98  &  n336 ) ;
 assign n465 = ( (~ P_174_97_)  &  n336 ) | ( n98  &  n336 ) ;
 assign n467 = ( (~ P_173_96_)  &  n336 ) | ( n98  &  n336 ) ;
 assign n469 = ( (~ P_175_98_)  &  n336 ) | ( n98  &  n336 ) ;
 assign n471 = ( (~ P_176_99_)  &  n336 ) | ( n98  &  n336 ) ;
 assign n474 = ( (~ n469) ) | ( n552 ) ;
 assign n476 = ( (~ P_2239_181_)  &  P_63_26_ ) | ( (~ P_2239_181_)  &  P_18_5_ ) | ( P_63_26_  &  (~ P_18_5_) ) ;
 assign n473 = ( (~ n471)  &  n474  &  n476 ) ;
 assign n477 = ( (~ P_177_100_)  &  n336 ) | ( n98  &  n336 ) ;
 assign n483 = ( (~ n639)  &  n886 ) | ( (~ n658)  &  n886 ) | ( n886  &  n888 ) ;
 assign n479 = ( n483  &  (~ n638)  &  (~ n1054) ) | ( n483  &  (~ n657)  &  (~ n1054) ) ;
 assign n484 = ( n320  &  n322  &  n321 ) ;
 assign n486 = ( P_201_124_  &  P_124_63_ ) | ( P_201_124_  &  P_18_5_ ) | ( P_124_63_  &  (~ P_18_5_) ) ;
 assign n487 = ( (~ P_3743_193_)  &  P_55_18_ ) | ( (~ P_3743_193_)  &  P_18_5_ ) | ( P_55_18_  &  (~ P_18_5_) ) ;
 assign n485 = ( n323  &  n484 ) | ( n323  &  n486  &  n487 ) ;
 assign n491 = ( (~ P_4394_196_)  &  P_77_36_ ) | ( (~ P_4394_196_)  &  P_18_5_ ) | ( P_77_36_  &  (~ P_18_5_) ) ;
 assign n492 = ( P_187_110_  &  P_118_61_ ) | ( P_187_110_  &  P_18_5_ ) | ( P_118_61_  &  (~ P_18_5_) ) ;
 assign n488 = ( n491  &  (~ n892) ) | ( n492  &  (~ n892) ) | ( n491  &  (~ n893) ) | ( n492  &  (~ n893) ) ;
 assign n493 = ( n492  &  n491 ) ;
 assign n495 = ( (~ P_4400_197_)  &  P_78_37_ ) | ( (~ P_4400_197_)  &  P_18_5_ ) | ( P_78_37_  &  (~ P_18_5_) ) ;
 assign n496 = ( P_196_119_  &  P_97_50_ ) | ( P_196_119_  &  P_18_5_ ) | ( P_97_50_  &  (~ P_18_5_) ) ;
 assign n494 = ( n488  &  n495 ) | ( n493  &  n495 ) | ( n488  &  n496 ) | ( n493  &  n496 ) ;
 assign n498 = ( (~ P_4405_198_)  &  P_59_22_ ) | ( (~ P_4405_198_)  &  P_18_5_ ) | ( P_59_22_  &  (~ P_18_5_) ) ;
 assign n499 = ( n503 ) | ( n502 ) ;
 assign n500 = ( P_195_118_  &  P_94_49_ ) | ( P_195_118_  &  P_18_5_ ) | ( P_94_49_  &  (~ P_18_5_) ) ;
 assign n497 = ( n498  &  n499  &  n500 ) ;
 assign n504 = ( n642 ) | ( n662 ) ;
 assign n502 = ( P_194_117_  &  P_121_62_ ) | ( P_194_117_  &  P_18_5_ ) | ( P_121_62_  &  (~ P_18_5_) ) ;
 assign n503 = ( (~ P_4410_199_)  &  P_81_40_ ) | ( (~ P_4410_199_)  &  P_18_5_ ) | ( P_81_40_  &  (~ P_18_5_) ) ;
 assign n501 = ( n504  &  n497 ) | ( n504  &  n502  &  n503 ) ;
 assign n506 = ( n504  &  n494 ) | ( n504  &  n496  &  n495 ) ;
 assign n505 = ( n499  &  n506  &  n498 ) | ( n499  &  n506  &  n500 ) ;
 assign n507 = ( (~ n501)  &  (~ n505)  &  (~ n642) ) | ( (~ n501)  &  (~ n505)  &  (~ n662) ) ;
 assign n515 = ( n858 ) | ( n859 ) ;
 assign n513 = ( (~ P_4420_201_)  &  P_79_38_ ) | ( (~ P_4420_201_)  &  P_18_5_ ) | ( P_79_38_  &  (~ P_18_5_) ) ;
 assign n514 = ( P_192_115_  &  P_35_10_ ) | ( P_192_115_  &  P_18_5_ ) | ( P_35_10_  &  (~ P_18_5_) ) ;
 assign n512 = ( (~ n507)  &  n515  &  n513 ) | ( (~ n507)  &  n515  &  n514 ) ;
 assign n517 = ( (~ n512)  &  (~ n858)  &  (~ n1060) ) | ( (~ n512)  &  (~ n859)  &  (~ n1060) ) ;
 assign n526 = ( n857 ) | ( n856 ) ;
 assign n523 = ( (~ P_4432_203_)  &  P_61_24_ ) | ( (~ P_4432_203_)  &  P_18_5_ ) | ( P_61_24_  &  (~ P_18_5_) ) ;
 assign n524 = ( P_190_113_  &  P_50_15_ ) | ( P_190_113_  &  P_18_5_ ) | ( P_50_15_  &  (~ P_18_5_) ) ;
 assign n522 = ( (~ n517)  &  n526  &  n523 ) | ( (~ n517)  &  n526  &  n524 ) ;
 assign n532 = ( (~ n99) ) | ( n536 ) ;
 assign n534 = ( (~ P_2211_176_)  &  P_65_28_ ) | ( (~ P_2211_176_)  &  P_18_5_ ) | ( P_65_28_  &  (~ P_18_5_) ) ;
 assign n531 = ( (~ n109)  &  n532  &  n534 ) ;
 assign n538 = ( (~ n103) ) | ( n540 ) ;
 assign n536 = ( (~ P_2218_177_)  &  P_83_42_ ) | ( (~ P_2218_177_)  &  P_18_5_ ) | ( P_83_42_  &  (~ P_18_5_) ) ;
 assign n535 = ( n531  &  n538 ) | ( (~ n99)  &  n538  &  n536 ) ;
 assign n542 = ( (~ n106) ) | ( n544 ) ;
 assign n540 = ( (~ P_2224_178_)  &  P_84_43_ ) | ( (~ P_2224_178_)  &  P_18_5_ ) | ( P_84_43_  &  (~ P_18_5_) ) ;
 assign n539 = ( n535  &  n542 ) | ( (~ n103)  &  n542  &  n540 ) ;
 assign n546 = ( (~ n477) ) | ( n649 ) ;
 assign n544 = ( (~ P_2230_179_)  &  P_85_44_ ) | ( (~ P_2230_179_)  &  P_18_5_ ) | ( P_85_44_  &  (~ P_18_5_) ) ;
 assign n543 = ( n539  &  n546 ) | ( (~ n106)  &  n546  &  n544 ) ;
 assign n547 = ( n477  &  (~ n543)  &  (~ n1062) ) | ( (~ n543)  &  (~ n649)  &  (~ n1062) ) ;
 assign n552 = ( (~ P_2247_182_)  &  P_86_45_ ) | ( (~ P_2247_182_)  &  P_18_5_ ) | ( P_86_45_  &  (~ P_18_5_) ) ;
 assign n551 = ( n316  &  n473 ) | ( n316  &  (~ n469)  &  n552 ) ;
 assign n557 = ( (~ n474)  &  (~ n551) ) | ( n547  &  (~ n551) ) | ( (~ n551)  &  (~ n895) ) ;
 assign n554 = ( n467  &  n557  &  (~ n1063) ) | ( n557  &  (~ n855)  &  (~ n1063) ) ;
 assign n561 = ( (~ n463) ) | ( n644 ) ;
 assign n559 = ( (~ P_1462_168_)  &  P_113_58_ ) | ( (~ P_1462_168_)  &  P_18_5_ ) | ( P_113_58_  &  (~ P_18_5_) ) ;
 assign n558 = ( (~ n98)  &  (~ n554)  &  n561 ) | ( (~ n554)  &  n561  &  n559 ) ;
 assign n563 = ( n463  &  (~ n558)  &  (~ n1064) ) | ( (~ n558)  &  (~ n644)  &  (~ n1064) ) ;
 assign n568 = ( (~ P_1480_170_)  &  P_112_57_ ) | ( (~ P_1480_170_)  &  P_18_5_ ) | ( P_112_57_  &  (~ P_18_5_) ) ;
 assign n567 = ( n459  &  (~ n1059) ) | ( (~ n455)  &  n568  &  (~ n1059) ) ;
 assign n573 = ( (~ n460) ) | ( n563 ) | ( (~ n616) ) | ( n1059 ) ;
 assign n571 = ( n453  &  (~ n567)  &  n573 ) | ( (~ n567)  &  n573  &  (~ n646) ) ;
 assign n576 = ( (~ P_4528_206_)  &  (~ n571) ) | ( P_1455_166_  &  (~ n571) ) | ( P_38_11_  &  (~ n571) ) ;
 assign n577 = ( (~ n123) ) | ( n718 ) ;
 assign n578 = ( (~ P_212_135_)  &  n336 ) | ( n98  &  n336 ) ;
 assign n580 = ( P_211_134_  &  (~ n98) ) | ( (~ P_18_5_)  &  (~ n98) ) ;
 assign n583 = ( P_70_31_ ) | ( P_18_5_ ) ;
 assign n581 = ( (~ P_3701_186_)  &  n583 ) | ( (~ P_18_5_)  &  n583 ) ;
 assign n584 = ( (~ P_165_88_)  &  n336 ) | ( n98  &  n336 ) ;
 assign n586 = ( P_164_87_  &  (~ n98) ) | ( (~ P_18_5_)  &  (~ n98) ) ;
 assign n587 = ( n140  &  n264 ) ;
 assign n589 = ( n259 ) | ( n606 ) ;
 assign n588 = ( n142  &  n589 ) ;
 assign n593 = ( (~ n135) ) | ( (~ n718) ) ;
 assign n590 = ( (~ n135)  &  n593 ) | ( (~ n259)  &  n593 ) ;
 assign n595 = ( (~ n126)  &  (~ n1021) ) | ( (~ n251)  &  (~ n1021) ) ;
 assign n598 = ( (~ n157)  &  (~ n451) ) | ( (~ n194)  &  (~ n451) ) ;
 assign n600 = ( (~ n148)  &  (~ n1028) ) | ( n598  &  (~ n1028) ) ;
 assign n603 = ( n131  &  (~ n396) ) | ( n131  &  (~ n734) ) ;
 assign n606 = ( (~ n142) ) | ( n715 ) ;
 assign n605 = ( n140  &  (~ n349) ) | ( n140  &  n606 ) ;
 assign n607 = ( n153  &  (~ n433) ) | ( n153  &  (~ n749) ) ;
 assign n610 = ( (~ n440) ) | ( n754 ) ;
 assign n609 = ( (~ n436) ) | ( n610 ) ;
 assign n611 = ( n167  &  (~ n448) ) | ( n167  &  (~ n702) ) ;
 assign n613 = ( n123  &  (~ n135) ) | ( n123  &  (~ n259)  &  (~ n718) ) ;
 assign n615 = ( (~ n109) ) | ( n534 ) ;
 assign n616 = ( (~ n457) ) | ( n462 ) ;
 assign n619 = ( n793  &  n167 ) ;
 assign n620 = ( (~ n770)  &  n792 ) ;
 assign n622 = ( n764  &  n760 ) ;
 assign n621 = ( n159  &  n622 ) ;
 assign n624 = ( n452  &  n621 ) ;
 assign n623 = ( n621  &  n624 ) | ( n621  &  n194 ) ;
 assign n625 = ( (~ n347)  &  n354 ) | ( n347  &  (~ n354) ) ;
 assign n626 = ( (~ n334)  &  n341 ) | ( n334  &  (~ n341) ) ;
 assign n627 = ( (~ n578)  &  n1056 ) | ( n578  &  (~ n1056) ) ;
 assign n629 = ( (~ P_239_162_)  &  (~ P_44_13_) ) | ( (~ P_239_162_)  &  P_18_5_ ) | ( (~ P_44_13_)  &  (~ P_18_5_) ) ;
 assign n630 = ( P_229_152_  &  P_41_12_ ) | ( P_229_152_  &  P_18_5_ ) | ( P_41_12_  &  (~ P_18_5_) ) ;
 assign n628 = ( (~ n629)  &  n630 ) | ( n629  &  (~ n630) ) ;
 assign n631 = ( (~ n441)  &  n437 ) | ( n441  &  (~ n437) ) ;
 assign n633 = ( (~ P_227_150_)  &  (~ P_115_60_) ) | ( (~ P_227_150_)  &  P_18_5_ ) | ( (~ P_115_60_)  &  (~ P_18_5_) ) ;
 assign n634 = ( P_217_140_  &  P_118_61_ ) | ( P_217_140_  &  P_18_5_ ) | ( P_118_61_  &  (~ P_18_5_) ) ;
 assign n632 = ( (~ n633)  &  n634 ) | ( n633  &  (~ n634) ) ;
 assign n635 = ( (~ n426)  &  n422 ) | ( n426  &  (~ n422) ) ;
 assign n636 = ( (~ n382)  &  n116 ) | ( n382  &  (~ n116) ) ;
 assign n638 = ( (~ P_3723_190_)  &  P_73_32_ ) | ( (~ P_3723_190_)  &  P_18_5_ ) | ( P_73_32_  &  (~ P_18_5_) ) ;
 assign n639 = ( (~ P_3717_189_)  &  P_75_34_ ) | ( (~ P_3717_189_)  &  P_18_5_ ) | ( P_75_34_  &  (~ P_18_5_) ) ;
 assign n637 = ( (~ n638)  &  n639 ) | ( n638  &  (~ n639) ) ;
 assign n640 = ( (~ n498)  &  n495 ) | ( n498  &  (~ n495) ) ;
 assign n642 = ( (~ P_4415_200_)  &  P_80_39_ ) | ( (~ P_4415_200_)  &  P_18_5_ ) | ( P_80_39_  &  (~ P_18_5_) ) ;
 assign n641 = ( (~ n642)  &  n503 ) | ( n642  &  (~ n503) ) ;
 assign n644 = ( (~ P_1469_169_)  &  P_111_56_ ) | ( (~ P_1469_169_)  &  P_18_5_ ) | ( P_111_56_  &  (~ P_18_5_) ) ;
 assign n643 = ( (~ n644)  &  n462 ) | ( n644  &  (~ n462) ) ;
 assign n646 = ( (~ P_1486_171_)  &  P_88_47_ ) | ( (~ P_1486_171_)  &  P_18_5_ ) | ( P_88_47_  &  (~ P_18_5_) ) ;
 assign n645 = ( (~ n646)  &  n568 ) | ( n646  &  (~ n568) ) ;
 assign n647 = ( (~ n540)  &  n536 ) | ( n540  &  (~ n536) ) ;
 assign n649 = ( (~ P_2236_180_)  &  P_64_27_ ) | ( (~ P_2236_180_)  &  P_18_5_ ) | ( P_64_27_  &  (~ P_18_5_) ) ;
 assign n648 = ( (~ n649)  &  n544 ) | ( n649  &  (~ n544) ) ;
 assign n650 = ( (~ n453)  &  n455 ) | ( n453  &  (~ n455) ) ;
 assign n651 = ( n457  &  n463 ) | ( (~ n457)  &  (~ n463) ) ;
 assign n652 = ( (~ n584)  &  n1055 ) | ( n584  &  (~ n1055) ) ;
 assign n654 = ( (~ P_208_131_)  &  (~ P_44_13_) ) | ( (~ P_208_131_)  &  P_18_5_ ) | ( (~ P_44_13_)  &  (~ P_18_5_) ) ;
 assign n655 = ( P_198_121_  &  P_41_12_ ) | ( P_198_121_  &  P_18_5_ ) | ( P_41_12_  &  (~ P_18_5_) ) ;
 assign n653 = ( (~ n654)  &  n655 ) | ( n654  &  (~ n655) ) ;
 assign n657 = ( P_204_127_  &  P_103_52_ ) | ( P_204_127_  &  P_18_5_ ) | ( P_103_52_  &  (~ P_18_5_) ) ;
 assign n658 = ( P_205_128_  &  P_23_6_ ) | ( P_205_128_  &  P_18_5_ ) | ( P_23_6_  &  (~ P_18_5_) ) ;
 assign n656 = ( (~ n657)  &  n658 ) | ( n657  &  (~ n658) ) ;
 assign n660 = ( (~ P_197_120_)  &  (~ P_115_60_) ) | ( (~ P_197_120_)  &  P_18_5_ ) | ( (~ P_115_60_)  &  (~ P_18_5_) ) ;
 assign n659 = ( (~ n660)  &  n492 ) | ( n660  &  (~ n492) ) ;
 assign n662 = ( P_193_116_  &  P_47_14_ ) | ( P_193_116_  &  P_18_5_ ) | ( P_47_14_  &  (~ P_18_5_) ) ;
 assign n661 = ( (~ n662)  &  n502 ) | ( n662  &  (~ n502) ) ;
 assign n663 = ( (~ n106)  &  n477 ) | ( n106  &  (~ n477) ) ;
 assign n667 = ( n256  &  n131 ) ;
 assign n668 = ( n794  &  n133 ) ;
 assign n671 = ( n724  &  n720 ) ;
 assign n670 = ( n375  &  n671 ) ;
 assign n673 = ( n732  &  n670 ) ;
 assign n672 = ( (~ n595)  &  n670 ) | ( n670  &  n673 ) ;
 assign n676 = ( n272  &  n153 ) ;
 assign n677 = ( (~ n784)  &  n795 ) ;
 assign n679 = ( n191  &  n776 ) ;
 assign n678 = ( n416  &  n679 ) ;
 assign n681 = ( n753  &  n678 ) ;
 assign n680 = ( (~ n600)  &  n678 ) | ( n678  &  n681 ) ;
 assign n683 = ( (~ n915)  &  n916 ) | ( n915  &  (~ n916) ) ;
 assign n684 = ( (~ n914)  &  n173 ) | ( n914  &  (~ n173) ) ;
 assign n686 = ( (~ n912)  &  n913 ) | ( n912  &  (~ n913) ) ;
 assign n685 = ( (~ n686)  &  n684 ) | ( n686  &  (~ n684) ) ;
 assign n689 = ( n744  &  n940 ) | ( (~ n744)  &  (~ n940) ) ;
 assign n687 = ( n689  &  n939 ) | ( (~ n689)  &  (~ n939) ) ;
 assign n690 = ( (~ n162)  &  (~ n451) ) | ( P_4526_205_  &  (~ n451)  &  (~ n609) ) ;
 assign n692 = ( (~ n935)  &  n936 ) | ( n935  &  (~ n936) ) ;
 assign n693 = ( (~ n940)  &  n744 ) | ( n940  &  (~ n744) ) ;
 assign n695 = ( (~ n950)  &  n951 ) | ( n950  &  (~ n951) ) ;
 assign n696 = ( n739  &  n952 ) | ( (~ n739)  &  (~ n952) ) ;
 assign n694 = ( (~ n695)  &  n696 ) | ( n695  &  (~ n696) ) ;
 assign n697 = ( (~ n953)  &  n954 ) | ( n953  &  (~ n954) ) ;
 assign n698 = ( n739  &  n955 ) | ( (~ n739)  &  (~ n955) ) ;
 assign n699 = ( (~ P_3701_186_) ) | ( P_18_5_ ) ;
 assign n700 = ( (~ P_18_5_)  &  n630 ) ;
 assign n703 = ( n700 ) | ( n699 ) ;
 assign n702 = ( n703  &  (~ n770) ) ;
 assign n706 = ( (~ P_4528_206_) ) | ( (~ P_1492_172_) ) ;
 assign n707 = ( (~ n122) ) | ( (~ n1023) ) ;
 assign n710 = ( n143 ) | ( (~ n356) ) ;
 assign n711 = ( (~ n343) ) | ( n710 ) ;
 assign n712 = ( n142 ) | ( (~ n349) ) | ( (~ n356) ) ;
 assign n713 = ( (~ n343) ) | ( n359 ) ;
 assign n715 = ( n352  &  P_1462_168_ ) ;
 assign n717 = ( (~ n349) ) | ( (~ n356) ) | ( n606 ) ;
 assign n718 = ( n260 ) | ( (~ n337) ) ;
 assign n720 = ( (~ n372) ) | ( n381 ) ;
 assign n722 = ( P_2239_181_ ) | ( n376 ) ;
 assign n723 = ( (~ n378) ) | ( n722 ) ;
 assign n724 = ( (~ n372) ) | ( n723 ) ;
 assign n726 = ( n376  &  P_2239_181_ ) ;
 assign n728 = ( (~ n388) ) | ( n395 ) ;
 assign n729 = ( n134 ) | ( (~ n392) ) ;
 assign n730 = ( n133 ) | ( (~ n392) ) | ( (~ n396) ) ;
 assign n731 = ( (~ n388) ) | ( n730 ) ;
 assign n732 = ( n173 ) | ( (~ n372) ) | ( (~ n378) ) ;
 assign n735 = ( (~ P_2211_176_) ) | ( (~ n118) ) ;
 assign n734 = ( n735  &  n133 ) ;
 assign n736 = ( (~ n392) ) | ( (~ n396) ) | ( (~ n734) ) ;
 assign n737 = ( n252 ) | ( (~ n384) ) ;
 assign n740 = ( (~ P_3729_191_) ) | ( n762 ) ;
 assign n739 = ( n740  &  (~ n761) ) ;
 assign n745 = ( (~ P_4420_201_) ) | ( n967 ) ;
 assign n746 = ( P_4420_201_ ) | ( (~ n967) ) ;
 assign n744 = ( n745  &  n746 ) ;
 assign n750 = ( (~ P_4394_196_) ) | ( n634 ) ;
 assign n749 = ( n750  &  (~ n784) ) ;
 assign n751 = ( (~ n429) ) | ( (~ n433) ) | ( (~ n749) ) ;
 assign n752 = ( n267 ) | ( (~ n421) ) ;
 assign n753 = ( (~ n413) ) | ( (~ n417) ) | ( (~ n744) ) ;
 assign n754 = ( (~ n444) ) | ( (~ n448) ) | ( (~ n702) ) ;
 assign n755 = ( (~ n409) ) | ( n752 ) | ( n753 ) ;
 assign n756 = ( (~ P_4526_205_) ) | ( (~ n399) ) | ( n452 ) | ( n609 ) | ( n755 ) ;
 assign n757 = ( (~ n366) ) | ( n732 ) | ( n737 ) ;
 assign n760 = ( (~ n402) ) | ( n408 ) ;
 assign n762 = ( P_234_157_  &  P_130_65_ ) | ( P_234_157_  &  P_18_5_ ) | ( P_130_65_  &  (~ P_18_5_) ) ;
 assign n761 = ( (~ P_3729_191_)  &  n762 ) ;
 assign n763 = ( (~ n405) ) | ( (~ n761) ) ;
 assign n764 = ( (~ n402) ) | ( n763 ) ;
 assign n765 = ( (~ P_3717_189_)  &  n441 ) ;
 assign n766 = ( (~ P_3711_188_)  &  n445 ) ;
 assign n767 = ( (~ n440) ) | ( (~ n766) ) ;
 assign n769 = ( n170 ) | ( (~ n444) ) ;
 assign n770 = ( n699  &  n700 ) ;
 assign n771 = ( (~ n444) ) | ( (~ n448) ) | ( (~ n770) ) ;
 assign n772 = ( (~ n440) ) | ( n771 ) ;
 assign n775 = ( (~ P_4427_202_)  &  n418 ) ;
 assign n776 = ( (~ n413) ) | ( (~ n775) ) ;
 assign n778 = ( (~ n417) ) | ( n746 ) ;
 assign n779 = ( (~ P_4410_199_)  &  n426 ) ;
 assign n781 = ( (~ n425) ) | ( n432 ) ;
 assign n783 = ( n156 ) | ( (~ n429) ) ;
 assign n784 = ( (~ P_4394_196_)  &  n634 ) ;
 assign n785 = ( (~ n429) ) | ( (~ n433) ) | ( (~ n784) ) ;
 assign n786 = ( (~ n425) ) | ( n785 ) ;
 assign n789 = ( (~ P_18_5_)  &  n655 ) ;
 assign n792 = ( (~ P_4526_205_) ) | ( (~ n702) ) ;
 assign n793 = ( (~ n448) ) | ( n792 ) ;
 assign n794 = ( n251 ) | ( (~ n734) ) ;
 assign n795 = ( (~ n598) ) | ( (~ n749) ) ;
 assign n796 = ( (~ n157) ) | ( n690 ) ;
 assign n797 = ( (~ n179)  &  n402 ) | ( n179  &  (~ n402) ) ;
 assign n798 = ( n405  &  n740 ) | ( (~ n405)  &  (~ n740) ) ;
 assign n799 = ( (~ n762)  &  n900 ) | ( n762  &  (~ n900) ) ;
 assign n800 = ( (~ n406)  &  n403 ) | ( n406  &  (~ n403) ) ;
 assign n801 = ( n901  &  n967 ) | ( (~ n901)  &  (~ n967) ) ;
 assign n802 = ( (~ n418)  &  n414 ) | ( n418  &  (~ n414) ) ;
 assign n803 = ( (~ n364)  &  n903 ) | ( n364  &  (~ n903) ) ;
 assign n804 = ( (~ n370)  &  n376 ) | ( n370  &  (~ n376) ) ;
 assign n805 = ( (~ n145)  &  n904 ) | ( n145  &  (~ n904) ) ;
 assign n806 = ( (~ n487)  &  n320 ) | ( n487  &  (~ n320) ) ;
 assign n808 = ( (~ n523)  &  n905 ) | ( n523  &  (~ n905) ) ;
 assign n809 = ( (~ n858)  &  n513 ) | ( n858  &  (~ n513) ) ;
 assign n807 = ( (~ n808)  &  n809 ) | ( n808  &  (~ n809) ) ;
 assign n810 = ( (~ P_1492_172_)  &  P_1455_166_ ) | ( (~ P_1492_172_)  &  P_18_5_ ) | ( P_1455_166_  &  (~ P_18_5_) ) ;
 assign n811 = ( (~ n200)  &  n906 ) | ( n200  &  (~ n906) ) ;
 assign n812 = ( (~ n317)  &  n907 ) | ( n317  &  (~ n907) ) ;
 assign n813 = ( (~ n552)  &  n476 ) | ( n552  &  (~ n476) ) ;
 assign n814 = ( (~ n146)  &  n908 ) | ( n146  &  (~ n908) ) ;
 assign n815 = ( (~ n486)  &  n321 ) | ( n486  &  (~ n321) ) ;
 assign n817 = ( (~ n524)  &  n909 ) | ( n524  &  (~ n909) ) ;
 assign n818 = ( (~ n859)  &  n514 ) | ( n859  &  (~ n514) ) ;
 assign n816 = ( (~ n817)  &  n818 ) | ( n817  &  (~ n818) ) ;
 assign n819 = ( n467  &  n910 ) | ( (~ n467)  &  (~ n910) ) ;
 assign n820 = ( (~ n469)  &  n471 ) | ( n469  &  (~ n471) ) ;
 assign n821 = ( (~ n171)  &  n372 ) | ( n171  &  (~ n372) ) ;
 assign n822 = ( (~ n726)  &  n378 ) | ( n726  &  (~ n378) ) ;
 assign n823 = ( (~ n175)  &  n413 ) | ( n175  &  (~ n413) ) ;
 assign n824 = ( n417  &  n745 ) | ( (~ n417)  &  (~ n745) ) ;
 assign n826 = ( (~ n923)  &  n924 ) | ( n923  &  (~ n924) ) ;
 assign n827 = ( (~ n922)  &  n925 ) | ( n922  &  (~ n925) ) ;
 assign n825 = ( (~ n826)  &  n827 ) | ( n826  &  (~ n827) ) ;
 assign n828 = ( n388  &  n825 ) | ( (~ n388)  &  (~ n825) ) ;
 assign n830 = ( (~ n917)  &  n920 ) | ( n917  &  (~ n920) ) ;
 assign n831 = ( (~ n922)  &  n921 ) | ( n922  &  (~ n921) ) ;
 assign n829 = ( (~ n830)  &  n831 ) | ( n830  &  (~ n831) ) ;
 assign n832 = ( (~ n388)  &  n829 ) | ( n388  &  (~ n829) ) ;
 assign n834 = ( (~ n932)  &  n933 ) | ( n932  &  (~ n933) ) ;
 assign n835 = ( (~ n931)  &  n934 ) | ( n931  &  (~ n934) ) ;
 assign n833 = ( (~ n834)  &  n835 ) | ( n834  &  (~ n835) ) ;
 assign n836 = ( (~ n343)  &  n833 ) | ( n343  &  (~ n833) ) ;
 assign n838 = ( (~ n926)  &  n929 ) | ( n926  &  (~ n929) ) ;
 assign n839 = ( (~ n931)  &  n930 ) | ( n931  &  (~ n930) ) ;
 assign n837 = ( (~ n838)  &  n839 ) | ( n838  &  (~ n839) ) ;
 assign n840 = ( (~ n343)  &  n837 ) | ( n343  &  (~ n837) ) ;
 assign n842 = ( (~ n947)  &  n948 ) | ( n947  &  (~ n948) ) ;
 assign n843 = ( (~ n946)  &  n949 ) | ( n946  &  (~ n949) ) ;
 assign n841 = ( (~ n842)  &  n843 ) | ( n842  &  (~ n843) ) ;
 assign n844 = ( (~ n425)  &  n841 ) | ( n425  &  (~ n841) ) ;
 assign n846 = ( (~ n941)  &  n944 ) | ( n941  &  (~ n944) ) ;
 assign n847 = ( (~ n946)  &  n945 ) | ( n946  &  (~ n945) ) ;
 assign n845 = ( (~ n846)  &  n847 ) | ( n846  &  (~ n847) ) ;
 assign n848 = ( (~ n425)  &  n845 ) | ( n425  &  (~ n845) ) ;
 assign n850 = ( (~ n956)  &  n957 ) | ( n956  &  (~ n957) ) ;
 assign n851 = ( (~ n958)  &  n959 ) | ( n958  &  (~ n959) ) ;
 assign n849 = ( (~ n850)  &  n851 ) | ( n850  &  (~ n851) ) ;
 assign n852 = ( n440  &  n849 ) | ( (~ n440)  &  (~ n849) ) ;
 assign n853 = ( n122  &  n854 ) | ( (~ n122)  &  (~ n854) ) ;
 assign n854 = ( n968  &  P_38_11_ ) | ( n968  &  P_1496_173_  &  P_4528_206_ ) ;
 assign n855 = ( (~ P_2256_184_)  &  P_110_55_ ) | ( (~ P_2256_184_)  &  P_18_5_ ) | ( P_110_55_  &  (~ P_18_5_) ) ;
 assign n856 = ( P_189_112_  &  P_66_29_ ) | ( P_189_112_  &  P_18_5_ ) | ( P_66_29_  &  (~ P_18_5_) ) ;
 assign n857 = ( (~ P_4437_204_)  &  P_62_25_ ) | ( (~ P_4437_204_)  &  P_18_5_ ) | ( P_62_25_  &  (~ P_18_5_) ) ;
 assign n858 = ( (~ P_4427_202_)  &  P_60_23_ ) | ( (~ P_4427_202_)  &  P_18_5_ ) | ( P_60_23_  &  (~ P_18_5_) ) ;
 assign n859 = ( P_191_114_  &  P_32_9_ ) | ( P_191_114_  &  P_18_5_ ) | ( P_32_9_  &  (~ P_18_5_) ) ;
 assign n861 = ( (~ P_3749_194_)  &  P_56_19_ ) | ( (~ P_3749_194_)  &  P_18_5_ ) | ( P_56_19_  &  (~ P_18_5_) ) ;
 assign n863 = ( P_200_123_  &  P_100_51_ ) | ( P_200_123_  &  P_18_5_ ) | ( P_100_51_  &  (~ P_18_5_) ) ;
 assign n870 = ( (~ n182)  &  n622 ) | ( n402  &  n622 ) ;
 assign n872 = ( (~ n194)  &  n797 ) | ( n194  &  (~ n870) ) | ( n797  &  (~ n870) ) ;
 assign n873 = ( (~ n194)  &  n798 ) | ( n194  &  n970 ) | ( n798  &  n970 ) ;
 assign n874 = ( (~ n174)  &  n671 ) | ( n372  &  n671 ) ;
 assign n876 = ( n595  &  n821 ) | ( (~ n595)  &  (~ n874) ) | ( n821  &  (~ n874) ) ;
 assign n877 = ( n595  &  n822 ) | ( (~ n595)  &  n1017 ) | ( n822  &  n1017 ) ;
 assign n878 = ( (~ n178)  &  n679 ) | ( n413  &  n679 ) ;
 assign n880 = ( n600  &  n823 ) | ( (~ n600)  &  (~ n878) ) | ( n823  &  (~ n878) ) ;
 assign n881 = ( n600  &  n824 ) | ( (~ n600)  &  n1019 ) | ( n824  &  n1019 ) ;
 assign n882 = ( (~ n590)  &  n853 ) | ( n590  &  n1036 ) | ( n853  &  n1036 ) ;
 assign n883 = ( (~ n409) ) | ( n416 ) ;
 assign n884 = ( (~ n366) ) | ( n720  &  n724 ) ;
 assign n885 = ( n756 ) | ( n757 ) ;
 assign n886 = ( (~ n312)  &  (~ n1053) ) | ( (~ n310)  &  (~ n1053) ) | ( (~ n311)  &  (~ n1053) ) ;
 assign n888 = ( (~ n638)  &  (~ n657) ) ;
 assign n889 = ( n309  &  n789 ) | ( n309  &  n583 ) ;
 assign n891 = ( (~ n144)  &  (~ n861) ) | ( n479  &  (~ n861) ) | ( (~ n144)  &  (~ n863) ) | ( n479  &  (~ n863) ) ;
 assign n892 = ( (~ P_89_48_)  &  n891 ) | ( (~ n144)  &  n891 ) | ( (~ n889)  &  n891 ) ;
 assign n893 = ( (~ n147)  &  (~ n485) ) | ( (~ n145)  &  (~ n485) ) | ( (~ n146)  &  (~ n485) ) ;
 assign n895 = ( n316  &  (~ n471) ) | ( n316  &  n476 ) ;
 assign n900 = ( (~ n230)  &  n400 ) | ( n230  &  (~ n400) ) ;
 assign n901 = ( n220  &  n410 ) | ( (~ n220)  &  (~ n410) ) ;
 assign n903 = ( (~ n210)  &  n362 ) | ( n210  &  (~ n362) ) ;
 assign n904 = ( (~ n240)  &  n861 ) | ( n240  &  (~ n861) ) ;
 assign n905 = ( n235  &  n857 ) | ( (~ n235)  &  (~ n857) ) ;
 assign n906 = ( P_2204_174_  &  (~ P_1496_173_) ) | ( (~ P_1496_173_)  &  P_18_5_ ) | ( P_2204_174_  &  (~ P_18_5_) ) ;
 assign n907 = ( (~ n195)  &  n855 ) | ( n195  &  (~ n855) ) ;
 assign n908 = ( (~ n245)  &  n863 ) | ( n245  &  (~ n863) ) ;
 assign n909 = ( n225  &  n856 ) | ( (~ n225)  &  (~ n856) ) ;
 assign n910 = ( n205  &  n465 ) | ( (~ n205)  &  (~ n465) ) ;
 assign n912 = ( (~ n171)  &  n673 ) | ( n171  &  (~ n673) ) ;
 assign n913 = ( (~ n726)  &  n366 ) | ( n726  &  (~ n366) ) ;
 assign n914 = ( (~ n372)  &  n378 ) | ( n372  &  (~ n378) ) ;
 assign n915 = ( n670  &  n722 ) | ( (~ n670)  &  (~ n722) ) ;
 assign n916 = ( (~ n366)  &  n174 ) | ( n366  &  (~ n174) ) ;
 assign n918 = ( n736  &  n257 ) ;
 assign n919 = ( n252  &  n253 ) ;
 assign n917 = ( (~ n918)  &  n919 ) | ( n918  &  (~ n919) ) ;
 assign n920 = ( n384  &  n735 ) | ( (~ n384)  &  (~ n735) ) ;
 assign n921 = ( (~ n734)  &  n603 ) | ( n734  &  (~ n603) ) ;
 assign n922 = ( (~ n392)  &  n396 ) | ( n392  &  (~ n396) ) ;
 assign n923 = ( (~ n133)  &  n131 ) | ( n133  &  (~ n131) ) ;
 assign n924 = ( (~ n384)  &  n253 ) | ( n384  &  (~ n253) ) ;
 assign n925 = ( (~ n257)  &  n734 ) | ( n257  &  (~ n734) ) ;
 assign n927 = ( n717  &  n265 ) ;
 assign n928 = ( n260  &  n261 ) ;
 assign n926 = ( (~ n927)  &  n928 ) | ( n927  &  (~ n928) ) ;
 assign n929 = ( (~ n715)  &  n337 ) | ( n715  &  (~ n337) ) ;
 assign n930 = ( (~ n356)  &  n605 ) | ( n356  &  (~ n605) ) ;
 assign n931 = ( n349  &  n606 ) | ( (~ n349)  &  (~ n606) ) ;
 assign n932 = ( n142  &  n140 ) | ( (~ n142)  &  (~ n140) ) ;
 assign n933 = ( (~ n337)  &  n261 ) | ( n337  &  (~ n261) ) ;
 assign n934 = ( (~ n265)  &  n356 ) | ( n265  &  (~ n356) ) ;
 assign n935 = ( (~ n175)  &  n681 ) | ( n175  &  (~ n681) ) ;
 assign n936 = ( (~ n745)  &  n409 ) | ( n745  &  (~ n409) ) ;
 assign n937 = ( (~ n678)  &  n746 ) | ( n678  &  (~ n746) ) ;
 assign n938 = ( (~ n409)  &  n178 ) | ( n409  &  (~ n178) ) ;
 assign n939 = ( (~ n937)  &  n938 ) | ( n937  &  (~ n938) ) ;
 assign n940 = ( (~ n413)  &  n417 ) | ( n413  &  (~ n417) ) ;
 assign n942 = ( n751  &  n273 ) ;
 assign n943 = ( n267  &  n269 ) ;
 assign n941 = ( (~ n942)  &  n943 ) | ( n942  &  (~ n943) ) ;
 assign n944 = ( n421  &  n750 ) | ( (~ n421)  &  (~ n750) ) ;
 assign n945 = ( (~ n749)  &  n607 ) | ( n749  &  (~ n607) ) ;
 assign n946 = ( (~ n429)  &  n433 ) | ( n429  &  (~ n433) ) ;
 assign n947 = ( (~ n784)  &  n153 ) | ( n784  &  (~ n153) ) ;
 assign n948 = ( (~ n421)  &  n269 ) | ( n421  &  (~ n269) ) ;
 assign n949 = ( (~ n273)  &  n749 ) | ( n273  &  (~ n749) ) ;
 assign n950 = ( (~ n621)  &  n761 ) | ( n621  &  (~ n761) ) ;
 assign n951 = ( (~ n399)  &  n182 ) | ( n399  &  (~ n182) ) ;
 assign n952 = ( (~ n402)  &  n405 ) | ( n402  &  (~ n405) ) ;
 assign n953 = ( (~ n179)  &  n624 ) | ( n179  &  (~ n624) ) ;
 assign n954 = ( n399  &  n740 ) | ( (~ n399)  &  (~ n740) ) ;
 assign n955 = ( (~ n402)  &  n405 ) | ( n402  &  (~ n405) ) ;
 assign n956 = ( (~ n770)  &  n167 ) | ( n770  &  (~ n167) ) ;
 assign n957 = ( n184  &  n702 ) | ( (~ n184)  &  (~ n702) ) ;
 assign n958 = ( (~ n436)  &  n444 ) | ( n436  &  (~ n444) ) ;
 assign n959 = ( (~ n187)  &  n448 ) | ( n187  &  (~ n448) ) ;
 assign n961 = ( n754  &  n187 ) ;
 assign n962 = ( n610  &  n184 ) ;
 assign n960 = ( (~ n961)  &  n962 ) | ( n961  &  (~ n962) ) ;
 assign n963 = ( (~ n436)  &  n440 ) | ( n436  &  (~ n440) ) ;
 assign n964 = ( n960  &  n963 ) | ( (~ n960)  &  (~ n963) ) ;
 assign n966 = ( (~ n444)  &  n448 ) | ( n444  &  (~ n448) ) ;
 assign n967 = ( P_222_145_  &  P_35_10_ ) | ( P_222_145_  &  P_18_5_ ) | ( P_35_10_  &  (~ P_18_5_) ) ;
 assign n968 = ( (~ P_4528_206_) ) | ( (~ P_1496_173_) ) | ( (~ P_38_11_) ) ;
 assign n970 = ( n405  &  n761 ) | ( (~ n405)  &  (~ n761) ) ;
 assign n971 = ( (~ n98)  &  n352 ) ;
 assign n972 = ( (~ n625)  &  (~ n626)  &  (~ n971) ) ;
 assign n976 = ( n625  &  (~ n626)  &  n971 ) ;
 assign n977 = ( (~ n625)  &  n626  &  n971 ) ;
 assign n978 = ( n625  &  n626  &  (~ n971) ) ;
 assign n981 = ( n445  &  n449 ) | ( (~ n445)  &  (~ n449) ) ;
 assign n984 = ( n430  &  n434 ) | ( (~ n430)  &  (~ n434) ) ;
 assign n987 = ( (~ P_161_84_)  &  (~ P_141_70_) ) | ( (~ P_161_84_)  &  P_18_5_ ) | ( (~ P_141_70_)  &  (~ P_18_5_) ) ;
 assign n988 = ( (~ n112)  &  n114 ) | ( n112  &  (~ n114) ) ;
 assign n990 = ( (~ P_3698_185_)  &  P_69_30_ ) | ( (~ P_3698_185_)  &  P_18_5_ ) | ( P_69_30_  &  (~ P_18_5_) ) ;
 assign n991 = ( (~ n324)  &  n310 ) | ( n324  &  (~ n310) ) ;
 assign n993 = ( P_4393_195_  &  (~ P_58_21_) ) | ( P_4393_195_  &  P_18_5_ ) | ( (~ P_58_21_)  &  (~ P_18_5_) ) ;
 assign n994 = ( (~ n993)  &  n491 ) | ( n993  &  (~ n491) ) ;
 assign n996 = ( P_1459_167_  &  (~ P_114_59_) ) | ( P_1459_167_  &  P_18_5_ ) | ( (~ P_114_59_)  &  (~ P_18_5_) ) ;
 assign n997 = ( (~ n996)  &  n559 ) | ( n996  &  (~ n559) ) ;
 assign n999 = ( P_2208_175_  &  (~ P_82_41_) ) | ( P_2208_175_  &  P_18_5_ ) | ( (~ P_82_41_)  &  (~ P_18_5_) ) ;
 assign n1000 = ( (~ n999)  &  n534 ) | ( n999  &  (~ n534) ) ;
 assign n1001 = ( P_170_93_ ) | ( (~ P_18_5_) ) | ( n98 ) ;
 assign n1002 = ( (~ n650)  &  n651  &  n1001 ) ;
 assign n1004 = ( (~ n650)  &  (~ n651)  &  (~ n1001) ) ;
 assign n1007 = ( n650  &  (~ n651)  &  n1001 ) ;
 assign n1008 = ( n650  &  n651  &  (~ n1001) ) ;
 assign n1010 = ( (~ n325)  &  n311 ) | ( n325  &  (~ n311) ) ;
 assign n1012 = ( (~ n500)  &  n496 ) | ( n500  &  (~ n496) ) ;
 assign n1014 = ( (~ P_181_104_)  &  (~ P_141_70_) ) | ( (~ P_181_104_)  &  P_18_5_ ) | ( (~ P_141_70_)  &  (~ P_18_5_) ) ;
 assign n1015 = ( (~ n99)  &  n103 ) | ( n99  &  (~ n103) ) ;
 assign n1017 = ( (~ n378)  &  n722 ) | ( n378  &  (~ n722) ) ;
 assign n1019 = ( (~ n417)  &  n746 ) | ( n417  &  (~ n746) ) ;
 assign n1020 = ( (~ n126) ) | ( (~ n251) ) | ( n279 ) ;
 assign n1021 = ( n737  &  n126 ) ;
 assign n1022 = ( n251  &  n828 ) | ( (~ n251)  &  n832 ) | ( n828  &  n832 ) ;
 assign n1024 = ( (~ n707) ) | ( n854 ) | ( (~ n1023) ) ;
 assign n1023 = ( P_38_11_ ) | ( n706 ) ;
 assign n1026 = ( n1042 ) | ( n593 ) ;
 assign n1027 = ( n259  &  n836 ) | ( (~ n259)  &  n840 ) | ( n836  &  n840 ) ;
 assign n1028 = ( n752  &  n148 ) ;
 assign n1030 = ( n687 ) | ( (~ n1028) ) ;
 assign n1031 = ( (~ n796)  &  n844 ) | ( n796  &  n848 ) | ( n844  &  n848 ) ;
 assign n1032 = ( (~ n162) ) | ( (~ n609) ) | ( n694 ) ;
 assign n1034 = ( (~ n966)  &  n1089 ) | ( n966  &  (~ n1089) ) ;
 assign n1033 = ( (~ n964)  &  n1034 ) | ( n964  &  (~ n1034) ) ;
 assign n1035 = ( (~ P_4526_205_)  &  n852 ) | ( P_4526_205_  &  n1033 ) | ( n852  &  n1033 ) ;
 assign n1036 = ( (~ n854)  &  n1023 ) | ( n854  &  (~ n1023) ) ;
 assign n1037 = ( n118  &  n987 ) | ( (~ n118)  &  (~ n987) ) ;
 assign n1039 = ( (~ n581)  &  n990 ) | ( n581  &  (~ n990) ) ;
 assign n1040 = ( (~ n1014)  &  n109 ) | ( n1014  &  (~ n109) ) ;
 assign n1043 = ( (~ n122) ) | ( (~ n707) ) ;
 assign n1042 = ( (~ n854)  &  n1043 ) | ( n854  &  (~ n1043) ) ;
 assign n1048 = ( P_147_72_  &  (~ P_18_5_) ) ;
 assign n1049 = ( P_144_71_  &  (~ P_18_5_) ) ;
 assign n1050 = ( P_138_69_  &  (~ P_18_5_) ) ;
 assign n1051 = ( P_135_68_  &  (~ P_18_5_) ) ;
 assign n1052 = ( (~ P_3749_194_)  &  n400 ) ;
 assign n1053 = ( n327  &  n324  &  n325  &  (~ n888) ) ;
 assign n1054 = ( n583  &  n309  &  n789 ) ;
 assign n1055 = ( n1007 ) | ( n1008 ) | ( n1002 ) | ( n1004 ) ;
 assign n1056 = ( n977 ) | ( n978 ) | ( n972 ) | ( n976 ) ;
 assign n1059 = ( n453  &  (~ n646) ) ;
 assign n1060 = ( n515  &  n513  &  n514 ) ;
 assign n1061 = ( n526  &  n523  &  n524 ) ;
 assign n1062 = ( (~ n291)  &  n532  &  n538  &  n542  &  n546  &  n615 ) ;
 assign n1063 = ( n319  &  n317  &  (~ n465) ) ;
 assign n1064 = ( (~ n98)  &  n561  &  n559 ) ;
 assign n1068 = ( n703  &  (~ n702) ) ;
 assign n1089 = ( (~ n611)  &  n1068 ) | ( n611  &  (~ n1068) ) ;
 assign P_560_248_ = ( P_3698_185_ ) ;
 assign P_558_244_ = ( P_3705_187_ ) ;
 assign P_556_242_ = ( P_3711_188_ ) ;
 assign P_554_240_ = ( P_3717_189_ ) ;
 assign P_552_238_ = ( P_3723_190_ ) ;
 assign P_550_236_ = ( P_3729_191_ ) ;
 assign P_548_234_ = ( P_3737_192_ ) ;
 assign P_546_232_ = ( P_3743_193_ ) ;
 assign P_544_230_ = ( P_3749_194_ ) ;
 assign P_542_246_ = ( P_3701_186_ ) ;
 assign P_540_227_ = ( P_4393_195_ ) ;
 assign P_538_224_ = ( P_4400_197_ ) ;
 assign P_536_222_ = ( P_4405_198_ ) ;
 assign P_534_220_ = ( P_4410_199_ ) ;
 assign P_532_218_ = ( P_4415_200_ ) ;
 assign P_530_216_ = ( P_4420_201_ ) ;
 assign P_528_214_ = ( P_4427_202_ ) ;
 assign P_526_212_ = ( P_4432_203_ ) ;
 assign P_524_210_ = ( P_4437_204_ ) ;
 assign P_522_226_ = ( P_4394_196_ ) ;
 assign P_496_271_ = ( P_2208_175_ ) ;
 assign P_494_267_ = ( P_2218_177_ ) ;
 assign P_492_265_ = ( P_2224_178_ ) ;
 assign P_490_263_ = ( P_2230_179_ ) ;
 assign P_488_260_ = ( P_2236_180_ ) ;
 assign P_486_258_ = ( P_2239_181_ ) ;
 assign P_484_256_ = ( P_2247_182_ ) ;
 assign P_482_253_ = ( P_2253_183_ ) ;
 assign P_480_250_ = ( P_2256_184_ ) ;
 assign P_478_269_ = ( P_2211_176_ ) ;
 assign P_471_3445_ = ( wire43 ) ;
 assign P_453_596_ = ( P_1_0_ ) ;
 assign P_450_288_ = ( P_1459_167_ ) ;
 assign P_448_284_ = ( P_1469_169_ ) ;
 assign P_446_393_ = ( P_106_53_ ) ;
 assign P_444_282_ = ( P_1480_170_ ) ;
 assign P_442_280_ = ( P_1486_171_ ) ;
 assign P_440_277_ = ( P_1492_172_ ) ;
 assign P_438_274_ = ( P_1496_173_ ) ;
 assign P_436_286_ = ( P_1462_168_ ) ;
 assign P_432_428_ = ( P_1_0_ ) ;
 assign P_419_3444_ = ( wire43 ) ;
 assign P_289_383_ = ( wire93 ) ;
 assign P_284_384_ = ( wire93 ) ;
 assign P_264_3121_ = ( wire101 ) ;
 assign P_258_3122_ = ( wire101 ) ;
 assign P_249_3418_ = ( wire101 ) ;
 assign P_3_312_ = ( P_1_0_ ) ;
 assign P_2_313_ = ( P_1_0_ ) ;


endmodule

