module C3540 (
	_77_9_, _87_10_, _169_22_, _238_31_, _2897_49_, _68_8_, _128_16_, _226_29_, 
	_294_39_, _326_44_, _58_7_, _190_24_, _264_35_, _283_38_, _250_33_, _329_45_, _213_26_, _257_34_, 
	_20_2_, _223_28_, _159_21_, _232_30_, _41_4_, _124_14_, _13_1_, _50_6_, _222_27_, _97_11_, 
	_125_15_, _322_43_, _244_32_, _274_37_, _317_42_, _1_0_, _33_3_, _270_36_, _200_25_, _343_47_, 
	_330_46_, _1698_48_, _132_17_, _45_5_, _116_13_, _143_19_, _303_40_, _311_41_, _107_12_, _137_18_, 
	_150_20_, _179_23_, _381_1626_, _351_1247_, _353_405_, _375_1624_, _393_1605_, _364_1484_, _369_1321_, _384_1553_, 
	_387_1616_, _358_1161_, _355_399_, _399_1428_, _402_1718_, _372_1243_, _396_1504_, _405_1717_, _409_1670_, _378_1597_, 
	_390_1603_, _361_940_, _367_1585_, _407_1657_);

input _77_9_, _87_10_, _169_22_, _238_31_, _2897_49_, _68_8_, _128_16_, _226_29_, _294_39_, _326_44_, _58_7_, _190_24_, _264_35_, _283_38_, _250_33_, _329_45_, _213_26_, _257_34_, _20_2_, _223_28_, _159_21_, _232_30_, _41_4_, _124_14_, _13_1_, _50_6_, _222_27_, _97_11_, _125_15_, _322_43_, _244_32_, _274_37_, _317_42_, _1_0_, _33_3_, _270_36_, _200_25_, _343_47_, _330_46_, _1698_48_, _132_17_, _45_5_, _116_13_, _143_19_, _303_40_, _311_41_, _107_12_, _137_18_, _150_20_, _179_23_;

output _381_1626_, _351_1247_, _353_405_, _375_1624_, _393_1605_, _364_1484_, _369_1321_, _384_1553_, _387_1616_, _358_1161_, _355_399_, _399_1428_, _402_1718_, _372_1243_, _396_1504_, _405_1717_, _409_1670_, _378_1597_, _390_1603_, _361_940_, _367_1585_, _407_1657_;

wire n_n1710, n_n1709, n_n1697, n_n1688, n_n1670, n_n1711, n_n1703, n_n1690, n_n1680, n_n1675, n_n1712, n_n1695, n_n1684, n_n1681, n_n1686, n_n1674, n_n1693, n_n1685, n_n1717, n_n1691, n_n1698, n_n1689, n_n1715, n_n1705, n_n1718, n_n1713, n_n1692, n_n1708, n_n1704, n_n1676, n_n1687, n_n1682, n_n1677, n_n1719, n_n1716, n_n1683, n_n1694, n_n1672, n_n1673, n_n1671, n_n1702, n_n1714, n_n1706, n_n1700, n_n1679, n_n1678, n_n1707, n_n1701, n_n1699, n_n1696, n_n613, n_n1419, n_n595, n_n1304, n_n1293, n_n1282, n_n1271, n_n1218, n_n1207, n_n1189, n_n571, n_n1166, n_n1155, n_n1144, n_n1133, n_n545, n_n1083, n_n1071, n_n1058, n_n534, n_n1033, n_n1017, n_n512, n_n502, n_n937, n_n477, n_n910, n_n466, n_n460, n_n453, n_n445, n_n435, n_n430, n_n813, n_n414, n_n785, n_n385, n_n378, n_n707, n_n368, n_n1663, n_n704, n_n756, n_n778, n_n790, n_n804, n_n818, n_n827, n_n844, n_n856, n_n863, n_n327, n_n320, n_n905, n_n703, n_n315, n_n304, n_n943, n_n970, n_n981, n_n994, n_n1004, n_n1018, n_n1030, n_n1043, n_n285, n_n1052, n_n274, n_n267, n_n1100, n_n251, n_n243, n_n235, n_n227, n_n220, n_n1125, n_n1177, n_n202, n_n191, n_n169, n_n158, n_n1202, n_n146, n_n135, n_n124, n_n113, n_n102, n_n77, n_n1308, n_n64, n_n56, n_n1380, n_n52, n_n47, n_n19, n_n1440, n_n1459, n_n1669, n_n1509, n_n700, n_n612, n_n607, n_n594, n_n1305, n_n1292, n_n1283, n_n1261, n_n1217, n_n1208, n_n1188, n_n572, n_n1165, n_n1156, n_n1143, n_n1134, n_n553, n_n1082, n_n1072, n_n1057, n_n535, n_n528, n_n520, n_n511, n_n503, n_n936, n_n478, n_n909, n_n467, n_n459, n_n454, n_n444, n_n436, n_n429, n_n421, n_n413, n_n407, n_n384, n_n379, n_n708, n_n369, n_n729, n_n366, n_n766, n_n781, n_n789, n_n805, n_n817, n_n828, n_n841, n_n857, n_n862, n_n326, n_n321, n_n906, n_n319, n_n314, n_n305, n_n945, n_n967, n_n993, n_n995, n_n1002, n_n1019, n_n1029, n_n1044, n_n1048, n_n1053, n_n275, n_n266, n_n260, n_n259, n_n1108, n_n236, n_n1114, n_n1117, n_n1126, n_n211, n_n201, n_n192, n_n168, n_n159, n_n1203, n_n147, n_n134, n_n125, n_n112, n_n103, n_n1237, n_n71, n_n65, n_n55, n_n1377, n_n51, n_n48, n_n18, n_n11, n_n1460, n_n1479, n_n1510, n_n1532, n_n1545, n_n1433, n_n608, n_n1317, n_n586, n_n1291, n_n1273, n_n1262, n_n1220, n_n1209, n_n1187, n_n569, n_n1168, n_n1157, n_n565, n_n554, n_n1081, n_n1068, n_n1060, n_n536, n_n527, n_n1011, n_n513, n_n504, n_n961, n_n489, n_n908, n_n464, n_n462, n_n873, n_n860, n_n437, n_n826, n_n420, n_n801, n_n408, n_n387, n_n380, n_n709, n_n716, n_n727, n_n738, n_n355, n_n347, n_n340, n_n807, n_n820, n_n825, n_n840, n_n872, n_n884, n_n322, n_n916, n_n925, n_n317, n_n306, n_n946, n_n979, n_n992, n_n1020, n_n1032, n_n1037, n_n286, n_n277, n_n273, n_n268, n_n261, n_n242, n_n1111, n_n1113, n_n221, n_n216, n_n210, n_n204, n_n193, n_n167, n_n156, n_n1200, n_n148, n_n133, n_n122, n_n115, n_n104, n_n83, n_n75, n_n1311, n_n1315, n_n1382, n_n1389, n_n49, n_n33, n_n1431, n_n1461, n_n701, n_n1507, n_n1531, n_n642, n_n614, n_n609, n_n596, n_n587, n_n1281, n_n1272, n_n1263, n_n1219, n_n1210, n_n1186, n_n570, n_n1167, n_n1158, n_n564, n_n555, n_n1080, n_n1069, n_n1059, n_n537, n_n526, n_n519, n_n1003, n_n505, n_n960, n_n950, n_n907, n_n465, n_n461, n_n874, n_n446, n_n849, n_n427, n_n812, n_n799, n_n788, n_n386, n_n719, n_n710, n_n367, n_n728, n_n737, n_n348, n_n346, n_n341, n_n808, n_n819, n_n428, n_n839, n_n330, n_n883, n_n885, n_n918, n_n479, n_n316, n_n307, n_n971, n_n980, n_n991, n_n1021, n_n1031, n_n1040, n_n287, n_n276, n_n1093, n_n1096, n_n1099, n_n241, n_n234, n_n228, n_n222, n_n215, n_n1178, n_n203, n_n194, n_n166, n_n157, n_n1201, n_n149, n_n132, n_n123, n_n114, n_n105, n_n82, n_n76, n_n1307, n_n54, n_n1381, n_n1390, n_n1404, n_n32, n_n26, n_n1462, n_n1484, n_n1508, n_n1526, n_n649, n_n643, n_n1435, n_n1423, n_n1319, n_n588, n_n582, n_n580, n_n1231, n_n1185, n_n1174, n_n1148, n_n1137, n_n567, n_n556, n_n1079, n_n541, n_n1054, n_n1041, n_n532, n_n522, n_n515, n_n506, n_n959, n_n487, n_n933, n_n473, n_n889, n_n875, n_n441, n_n433, n_n837, n_n424, n_n416, n_n409, n_n724, n_n374, n_n705, n_n714, n_n723, n_n736, n_n343, n_n339, n_n798, n_n814, n_n337, n_n834, n_n887, n_n897, n_n922, n_n932, n_n308, n_n996, n_n1009, n_n1035, n_n1047, n_n256, n_n248, n_n1116, n_n214, n_n187, n_n176, n_n131, n_n120, n_n98, n_n1229, n_n53, n_n1384, n_n1392, n_n44, n_n38, n_n1465, n_n1492, n_n1515, n_n1537, n_n1656, n_n1546, n_n1533, n_n615, n_n1424, n_n1318, n_n589, n_n1252, n_n1243, n_n1221, n_n1184, n_n1175, n_n1147, n_n1138, n_n566, n_n557, n_n1078, n_n1067, n_n540, n_n1042, n_n531, n_n523, n_n514, n_n507, n_n958, n_n488, n_n482, n_n474, n_n463, n_n876, n_n440, n_n842, n_n836, n_n425, n_n415, n_n410, n_n382, n_n375, n_n371, n_n713, n_n726, n_n735, n_n342, n_n794, n_n800, n_n811, n_n336, n_n833, n_n888, n_n896, n_n901, n_n318, n_n309, n_n997, n_n1007, n_n1036, n_n288, n_n255, n_n1105, n_n229, n_n209, n_n186, n_n177, n_n130, n_n121, n_n97, n_n1222, n_n1316, n_n1383, n_n45, n_n1407, n_n39, n_n1467, n_n1489, n_n1518, n_n1536, n_n651, n_n644, n_n1437, n_n1425, n_n590, n_n1251, n_n1233, n_n575, n_n1164, n_n1153, n_n1146, n_n1135, n_n1128, n_n558, n_n1077, n_n1063, n_n1056, n_n533, n_n530, n_n521, n_n1008, n_n508, n_n957, n_n944, n_n935, n_n475, n_n912, n_n468, n_n443, n_n843, n_n835, n_n422, n_n806, n_n792, n_n383, n_n376, n_n1662, n_n370, n_n721, n_n733, n_n345, n_n793, n_n802, n_n816, n_n823, n_n832, n_n1664, n_n895, n_n902, n_n924, n_n310, n_n295, n_n1006, n_n1015, n_n1028, n_n258, n_n249, n_n1110, n_n200, n_n189, n_n178, n_n111, n_n100, n_n89, n_n1370, n_n50, n_n46, n_n702, n_n1499, n_n1511, n_n1534, n_n650, n_n1535, n_n616, n_n610, n_n1320, n_n1241, n_n1232, n_n1223, n_n1163, n_n1154, n_n568, n_n1136, n_n1127, n_n559, n_n1076, n_n1064, n_n1055, n_n1045, n_n529, n_n1023, n_n516, n_n509, n_n956, n_n486, n_n934, n_n476, n_n911, n_n469, n_n442, n_n434, n_n431, n_n423, n_n417, n_n411, n_n725, n_n377, n_n706, n_n715, n_n722, n_n732, n_n344, n_n791, n_n803, n_n815, n_n338, n_n831, n_n886, n_n894, n_n903, n_n923, n_n931, n_n294, n_n1005, n_n1016, n_n1027, n_n257, n_n250, n_n244, n_n190, n_n188, n_n179, n_n110, n_n101, n_n99, n_n1385, n_n1391, n_n1406, n_n7, n_n1495, n_n1512, n_n6, n_n685, n_n640, n_n1514, n_n1503, n_n626, n_n1481, n_n1416, n_n1405, n_n598, n_n1365, n_n1354, n_n1343, n_n1332, n_n1321, n_n1290, n_n1279, n_n584, n_n1257, n_n1246, n_n1235, n_n1224, n_n1152, n_n1141, n_n1130, n_n560, n_n548, n_n1086, n_n1000, n_n498, n_n966, n_n782, n_n770, n_n755, n_n391, n_n743, n_n760, n_n768, n_n776, n_n847, n_n335, n_n866, n_n878, n_n323, n_n947, n_n297, n_n984, n_n1666, n_n1014, n_n272, n_n265, n_n253, n_n1107, n_n237, n_n199, n_n183, n_n172, n_n161, n_n1199, n_n94, n_n86, n_n78, n_n1269, n_n66, n_n43, n_n35, n_n29, n_n21, n_n13, n_n1453, n_n693, n_n686, n_n1524, n_n637, n_n1502, n_n1493, n_n1471, n_n1415, n_n601, n_n597, n_n1366, n_n1353, n_n1344, n_n1331, n_n1322, n_n1300, n_n1278, n_n585, n_n1256, n_n581, n_n1234, n_n1225, n_n1151, n_n1142, n_n1129, n_n561, n_n547, n_n1087, n_n517, n_n497, n_n492, n_n780, n_n771, n_n753, n_n742, n_n744, n_n758, n_n359, n_n352, n_n848, n_n858, n_n867, n_n877, n_n900, n_n300, n_n296, n_n983, n_n1001, n_n1013, n_n1094, n_n1097, n_n252, n_n1106, n_n230, n_n208, n_n182, n_n173, n_n160, n_n1198, n_n93, n_n1230, n_n1247, n_n72, n_n59, n_n42, n_n36, n_n1430, n_n22, n_n12, n_n1452, n_n1658, n_n677, n_n1614, n_n1523, n_n636, n_n629, n_n1494, n_n1454, n_n1414, n_n1403, n_n1395, n_n1367, n_n1352, n_n1341, n_n1334, n_n1323, n_n1299, n_n1288, n_n1270, n_n1255, n_n1244, n_n579, n_n1226, n_n1212, n_n1194, n_n1150, n_n1139, n_n1132, n_n562, n_n550, n_n1088, n_n524, n_n986, n_n968, n_n779, n_n401, n_n398, n_n392, n_n381, n_n745, n_n364, n_n361, n_n353, n_n786, n_n797, n_n850, n_n333, n_n864, n_n328, n_n325, n_n899, n_n939, n_n949, n_n982, n_n998, n_n1012, n_n281, n_n1066, n_n1103, n_n246, n_n223, n_n1145, n_n185, n_n174, n_n151, n_n140, n_n96, n_n87, n_n1253, n_n1310, n_n1313, n_n1408, n_n37, n_n28, n_n1434, n_n14, n_n1447, n_n1657, n_n676, n_n1615, n_n639, n_n1513, n_n1504, n_n627, n_n618, n_n1413, n_n600, n_n599, n_n1368, n_n1351, n_n1342, n_n1333, n_n1324, n_n1298, n_n1289, n_n1280, n_n1254, n_n1245, n_n578, n_n1227, n_n1211, n_n573, n_n1149, n_n1140, n_n1131, n_n563, n_n549, n_n1089, n_n1038, n_n985, n_n969, n_n406, n_n769, n_n397, n_n393, n_n373, n_n746, n_n365, n_n360, n_n773, n_n787, n_n796, n_n851, n_n334, n_n865, n_n329, n_n324, n_n898, n_n940, n_n948, n_n973, n_n999, n_n1010, n_n1050, n_n1065, n_n254, n_n247, n_n1119, n_n1120, n_n184, n_n175, n_n150, n_n141, n_n95, n_n88, n_n1306, n_n67, n_n60, n_n1410, n_n1420, n_n27, n_n20, n_n1438, n_n1443, n_n692, n_n1600, n_n1589, n_n1521, n_n1485, n_n1474, n_n1457, n_n1441, n_n1412, n_n1401, n_n1374, n_n1361, n_n1358, n_n1347, n_n1336, n_n1325, n_n591, n_n1297, n_n1286, n_n1275, n_n1264, n_n1250, n_n1239, n_n1228, n_n1214, n_n574, n_n1193, n_n1182, n_n1170, n_n1159, n_n1101, n_n542, n_n538, n_n500, n_n493, n_n405, n_n765, n_n750, n_n388, n_n711, n_n747, n_n761, n_n772, n_n777, n_n809, n_n822, n_n852, n_n332, n_n870, n_n882, n_n919, n_n927, n_n311, n_n299, n_n954, n_n977, n_n990, n_n1022, n_n292, n_n290, n_n282, n_n280, n_n1075, n_n1095, n_n262, n_n240, n_n232, n_n1115, n_n217, n_n1121, n_n1176, n_n206, n_n195, n_n165, n_n1668, n_n153, n_n142, n_n139, n_n128, n_n117, n_n106, n_n90, n_n81, n_n1268, n_n69, n_n61, n_n1372, n_n1387, n_n1398, n_n1417, n_n34, n_n1427, n_n24, n_n16, n_n8, n_n1505, n_n1525, n_n695, n_n665, n_n661, n_n635, n_n624, n_n622, n_n1456, n_n619, n_n605, n_n1402, n_n1373, n_n1362, n_n1357, n_n1348, n_n1335, n_n1326, n_n1301, n_n1296, n_n1287, n_n1274, n_n1265, n_n583, n_n1238, n_n576, n_n1213, n_n1204, n_n1192, n_n1183, n_n1169, n_n1160, n_n551, n_n543, n_n1061, n_n987, n_n494, n_n404, n_n767, n_n396, n_n389, n_n717, n_n748, n_n363, n_n356, n_n349, n_n810, n_n821, n_n853, n_n859, n_n871, n_n881, n_n920, n_n926, n_n301, n_n298, n_n953, n_n978, n_n989, n_n1024, n_n293, n_n289, n_n283, n_n279, n_n1070, n_n269, n_n263, n_n1109, n_n233, n_n224, n_n218, n_n1122, n_n1173, n_n205, n_n196, n_n164, n_n1195, n_n152, n_n143, n_n138, n_n129, n_n116, n_n107, n_n1236, n_n1242, n_n1260, n_n68, n_n62, n_n58, n_n1388, n_n1394, n_n40, n_n1426, n_n1429, n_n25, n_n15, n_n9, n_n1506, n_n1522, n_n696, n_n1579, n_n1562, n_n1501, n_n1483, n_n1472, n_n1464, n_n1444, n_n604, n_n1399, n_n1379, n_n1363, n_n1356, n_n1345, n_n1338, n_n1327, n_n593, n_n1302, n_n1295, n_n1284, n_n1277, n_n1266, n_n1259, n_n1248, n_n577, n_n1216, n_n1205, n_n1191, n_n1180, n_n1172, n_n1161, n_n552, n_n1092, n_n1073, n_n775, n_n762, n_n752, n_n390, n_n730, n_n749, n_n764, n_n358, n_n350, n_n829, n_n846, n_n854, n_n861, n_n868, n_n880, n_n921, n_n313, n_n302, n_n941, n_n964, n_n974, n_n988, n_n1025, n_n1034, n_n1667, n_n1049, n_n278, n_n1091, n_n271, n_n1098, n_n1104, n_n239, n_n1112, n_n226, n_n1118, n_n1123, n_n212, n_n1179, n_n197, n_n181, n_n170, n_n163, n_n1197, n_n155, n_n144, n_n137, n_n126, n_n119, n_n108, n_n92, n_n84, n_n80, n_n73, n_n70, n_n1312, n_n1314, n_n1376, n_n1393, n_n41, n_n1422, n_n31, n_n1432, n_n17, n_n10, n_n1455, n_n1475, n_n1660, n_n1578, n_n1563, n_n1491, n_n1482, n_n621, n_n1463, n_n1445, n_n1409, n_n1400, n_n1378, n_n1364, n_n1355, n_n1346, n_n1337, n_n1328, n_n592, n_n1303, n_n1294, n_n1285, n_n1276, n_n1267, n_n1258, n_n1249, n_n1240, n_n1215, n_n1206, n_n1190, n_n1181, n_n1171, n_n1162, n_n1102, n_n544, n_n1084, n_n774, n_n400, n_n751, n_n739, n_n740, n_n754, n_n763, n_n357, n_n351, n_n830, n_n845, n_n855, n_n331, n_n869, n_n879, n_n929, n_n312, n_n303, n_n942, n_n1665, n_n975, n_n499, n_n1026, n_n291, n_n1046, n_n284, n_n1051, n_n1090, n_n270, n_n264, n_n245, n_n238, n_n231, n_n225, n_n219, n_n1124, n_n213, n_n207, n_n198, n_n180, n_n171, n_n162, n_n1196, n_n154, n_n145, n_n136, n_n127, n_n118, n_n109, n_n91, n_n85, n_n79, n_n74, n_n1309, n_n63, n_n57, n_n1375, n_n1386, n_n1411, n_n1421, n_n30, n_n23, n_n1436, n_n1442, n_n1458, n_n1473, n_n1659, n_n690, n_n682, n_n673, n_n668, n_n662, n_n658, n_n654, n_n1500, n_n625, n_n1478, n_n620, n_n1446, n_n1340, n_n1329, n_n1544, n_n1559, n_n1577, n_n5, n_n1613, n_n694, n_n1638, n_n674, n_n667, n_n1594, n_n1580, n_n655, n_n634, n_n1488, n_n623, n_n1466, n_n1448, n_n1339, n_n1330, n_n1542, n_n1561, n_n1576, n_n1603, n_n1612, n_n1651, n_n684, n_n1623, n_n1602, n_n1591, n_n1584, n_n1567, n_n1520, n_n1487, n_n1476, n_n1469, n_n1449, n_n1360, n_n1349, n_n1541, n_n1564, n_n1583, n_n1599, n_n1611, n_n689, n_n683, n_n675, n_n666, n_n1592, n_n1582, n_n656, n_n1530, n_n1486, n_n1477, n_n1468, n_n1450, n_n1359, n_n1350, n_n1540, n_n1565, n_n1581, n_n1601, n_n1610, n_n1661, n_n688, n_n679, n_n1616, n_n670, n_n664, n_n659, n_n1572, n_n1529, n_n638, n_n631, n_n1496, n_n1451, n_n1397, n_n1369, n_n495, n_n962, n_n399, n_n394, n_n354, n_n1539, n_n4, n_n1634, n_n1644, n_n1655, n_n1650, n_n678, n_n671, n_n1609, n_n1598, n_n1585, n_n1573, n_n1528, n_n1519, n_n630, n_n1497, n_n1470, n_n1396, n_n1371, n_n972, n_n963, n_n759, n_n395, n_n362, n_n1538, n_n1625, n_n1633, n_n1645, n_n691, n_n687, n_n681, n_n672, n_n1607, n_n663, n_n660, n_n657, n_n1527, n_n1516, n_n633, n_n1498, n_n1480, n_n1418, n_n602, n_n546, n_n976, n_n491, n_n784, n_n402, n_n757, n_n1626, n_n1636, n_n2, n_n1654, n_n1647, n_n680, n_n1619, n_n669, n_n1596, n_n1587, n_n1575, n_n641, n_n1517, n_n632, n_n628, n_n1490, n_n606, n_n603, n_n1085, n_n496, n_n965, n_n783, n_n403, n_n741, n_n3, n_n1635, n_n1, n_n697, n_n652, n_n645, n_n1439, n_n611, n_n1074, n_n955, n_n484, n_n481, n_n913, n_n419, n_n795, n_n731, n_n1586, n_n1604, n_n1620, n_n1630, n_n1642, n_n1653, n_n1550, n_n646, n_n617, n_n1428, n_n1062, n_n490, n_n485, n_n480, n_n914, n_n418, n_n412, n_n718, n_n1588, n_n699, n_n1621, n_n1629, n_n1643, n_n0, n_n653, n_n647, n_n539, n_n952, n_n938, n_n930, n_n915, n_n432, n_n426, n_n712, n_n1552, n_n1568, n_n1622, n_n1632, n_n1640, n_n1652, n_n1556, n_n648, n_n1039, n_n951, n_n483, n_n928, n_n917, n_n838, n_n824, n_n372, n_n1553, n_n1566, n_n1624, n_n1631, n_n1641, n_n1649, n_n1543, n_n525, n_n472, n_n892, n_n456, n_n449, n_n448, n_n438, n_n720, n_n1551, n_n1554, n_n1570, n_n1595, n_n698, n_n1637, n_n1648, n_n1560, n_n518, n_n904, n_n893, n_n455, n_n450, n_n447, n_n439, n_n734, n_n1549, n_n1555, n_n1569, n_n1597, n_n1608, n_n1639, n_n1646, n_n510, n_n471, n_n890, n_n458, n_n451, n_n1548, n_n1557, n_n1574, n_n1590, n_n1606, n_n1617, n_n1628, n_n501, n_n470, n_n891, n_n457, n_n452, n_n1547, n_n1558, n_n1571, n_n1593, n_n1605, n_n1618, n_n1627;

assign n_n1710 = ( _77_9_ ) ;
 assign _381_1626_ = ( n_n751 ) ;
 assign n_n1709 = ( _87_10_ ) ;
 assign n_n1697 = ( _169_22_ ) ;
 assign n_n1688 = ( _238_31_ ) ;
 assign _351_1247_ = ( n_n1666 ) ;
 assign n_n1670 = ( _2897_49_ ) ;
 assign n_n1711 = ( _68_8_ ) ;
 assign n_n1703 = ( _128_16_ ) ;
 assign _353_405_ = ( n_n1669 ) ;
 assign _375_1624_ = ( n_n752 ) ;
 assign n_n1690 = ( _226_29_ ) ;
 assign n_n1680 = ( _294_39_ ) ;
 assign n_n1675 = ( _326_44_ ) ;
 assign n_n1712 = ( _58_7_ ) ;
 assign n_n1695 = ( _190_24_ ) ;
 assign n_n1684 = ( _264_35_ ) ;
 assign n_n1681 = ( _283_38_ ) ;
 assign n_n1686 = ( _250_33_ ) ;
 assign n_n1674 = ( _329_45_ ) ;
 assign _393_1605_ = ( n_n765 ) ;
 assign n_n1693 = ( _213_26_ ) ;
 assign _364_1484_ = ( n_n849 ) ;
 assign n_n1685 = ( _257_34_ ) ;
 assign n_n1717 = ( _20_2_ ) ;
 assign n_n1691 = ( _223_28_ ) ;
 assign n_n1698 = ( _159_21_ ) ;
 assign n_n1689 = ( _232_30_ ) ;
 assign n_n1715 = ( _41_4_ ) ;
 assign _369_1321_ = ( n_n1665 ) ;
 assign _384_1553_ = ( n_n801 ) ;
 assign n_n1705 = ( _124_14_ ) ;
 assign _387_1616_ = ( n_n759 ) ;
 assign n_n1718 = ( _13_1_ ) ;
 assign n_n1713 = ( _50_6_ ) ;
 assign n_n1692 = ( _222_27_ ) ;
 assign n_n1708 = ( _97_11_ ) ;
 assign n_n1704 = ( _125_15_ ) ;
 assign n_n1676 = ( _322_43_ ) ;
 assign n_n1687 = ( _244_32_ ) ;
 assign n_n1682 = ( _274_37_ ) ;
 assign n_n1677 = ( _317_42_ ) ;
 assign _358_1161_ = ( n_n1667 ) ;
 assign n_n1719 = ( _1_0_ ) ;
 assign n_n1716 = ( _33_3_ ) ;
 assign n_n1683 = ( _270_36_ ) ;
 assign _355_399_ = ( n_n1569 ) ;
 assign _399_1428_ = ( n_n1664 ) ;
 assign n_n1694 = ( _200_25_ ) ;
 assign n_n1672 = ( _343_47_ ) ;
 assign _402_1718_ = ( n_n1662 ) ;
 assign n_n1673 = ( _330_46_ ) ;
 assign _372_1243_ = ( n_n1003 ) ;
 assign _396_1504_ = ( n_n835 ) ;
 assign n_n1671 = ( _1698_48_ ) ;
 assign n_n1702 = ( _132_17_ ) ;
 assign _405_1717_ = ( n_n705 ) ;
 assign n_n1714 = ( _45_5_ ) ;
 assign n_n1706 = ( _116_13_ ) ;
 assign n_n1700 = ( _143_19_ ) ;
 assign n_n1679 = ( _303_40_ ) ;
 assign n_n1678 = ( _311_41_ ) ;
 assign n_n1707 = ( _107_12_ ) ;
 assign _409_1670_ = ( n_n1663 ) ;
 assign n_n1701 = ( _137_18_ ) ;
 assign n_n1699 = ( _150_20_ ) ;
 assign _378_1597_ = ( n_n769 ) ;
 assign _390_1603_ = ( n_n767 ) ;
 assign _361_940_ = ( n_n1668 ) ;
 assign _367_1585_ = ( n_n775 ) ;
 assign n_n1696 = ( _179_23_ ) ;
 assign _407_1657_ = ( n_n704 ) ;
 assign n_n613 = ( n_n27  &  n_n26  &  n_n28 ) ;
 assign n_n1419 = ( n_n1463  &  n_n1658 ) ;
 assign n_n595 = ( n_n56  &  n_n55  &  n_n57 ) ;
 assign n_n1304 = ( n_n1385  &  n_n1698 ) ;
 assign n_n1293 = ( n_n1382  &  n_n1699 ) ;
 assign n_n1282 = ( n_n1386  &  n_n1701 ) ;
 assign n_n1271 = ( n_n1385  &  n_n1704 ) ;
 assign n_n1218 = ( n_n1382  &  n_n1713 ) ;
 assign n_n1207 = ( n_n128  &  n_n127  &  n_n130  &  n_n129  &  n_n131  &  n_n124  &  n_n126  &  n_n125 ) ;
 assign n_n1189 = ( n_n1222  &  n_n658 ) ;
 assign n_n571 = ( n_n1253  &  n_n1268 ) ;
 assign n_n1166 = ( n_n585  &  n_n1203  &  n_n1695 ) ;
 assign n_n1155 = ( n_n1236  &  n_n1198  &  n_n1696 ) ;
 assign n_n1144 = ( n_n1461  &  n_n1204 ) ;
 assign n_n1133 = ( n_n1716  &  n_n1209 ) ;
 assign n_n545 = ( n_n272  &  n_n273 ) ;
 assign n_n1083 = ( n_n1105  &  n_n658 ) ;
 assign n_n1071 = ( n_n1105  &  n_n1197  &  n_n1696 ) ;
 assign n_n1058 = ( n_n1394  &  n_n1097 ) ;
 assign n_n534 = ( n_n1065  &  n_n1176 ) ;
 assign n_n1033 = ( n_n1399  &  n_n1047 ) ;
 assign n_n1017 = ( n_n1073  &  n_n1038  &  n_n1072  &  n_n1069 ) ;
 assign n_n512 = ( n_n1024  &  n_n1037  &  n_n1021  &  n_n1075 ) ;
 assign n_n502 = ( n_n1025  &  n_n1004 ) ;
 assign n_n937 = ( n_n305  &  n_n304  &  n_n306 ) ;
 assign n_n477 = ( n_n980  &  n_n1000 ) ;
 assign n_n910 = ( n_n1396  &  n_n935 ) ;
 assign n_n466 = ( n_n979  &  n_n918 ) ;
 assign n_n460 = ( n_n903  &  n_n901 ) ;
 assign n_n453 = ( n_n931  &  n_n885 ) ;
 assign n_n445 = ( n_n888  &  n_n872 ) ;
 assign n_n435 = ( n_n853  &  n_n951 ) ;
 assign n_n430 = ( n_n855  &  n_n845 ) ;
 assign n_n813 = ( n_n860  &  n_n831 ) ;
 assign n_n414 = ( n_n823  &  n_n804 ) ;
 assign n_n785 = ( n_n1398  &  n_n798 ) ;
 assign n_n385 = ( n_n736  &  n_n743 ) ;
 assign n_n378 = ( n_n722  &  n_n718 ) ;
 assign n_n707 = ( (~ n_n373) ) ;
 assign n_n368 = ( (~ n_n725) ) ;
 assign n_n1663 = ( (~ n_n734) ) ;
 assign n_n704 = ( (~ n_n742) ) ;
 assign n_n756 = ( (~ n_n397) ) ;
 assign n_n778 = ( (~ n_n406) ) ;
 assign n_n790 = ( (~ n_n796) ) ;
 assign n_n804 = ( (~ n_n416) ) ;
 assign n_n818 = ( (~ n_n424) ) ;
 assign n_n827 = ( (~ n_n839) ) ;
 assign n_n844 = ( (~ n_n434) ) ;
 assign n_n856 = ( (~ n_n443) ) ;
 assign n_n863 = ( (~ n_n449) ) ;
 assign n_n327 = ( (~ n_n907) ) ;
 assign n_n320 = ( (~ n_n1369) ) ;
 assign n_n905 = ( (~ n_n951) ) ;
 assign n_n703 = ( (~ n_n1000) ) ;
 assign n_n315 = ( (~ n_n1055) ) ;
 assign n_n304 = ( (~ n_n1371) ) ;
 assign n_n943 = ( (~ n_n968) ) ;
 assign n_n970 = ( (~ n_n493) ) ;
 assign n_n981 = ( (~ n_n995) ) ;
 assign n_n994 = ( (~ n_n504) ) ;
 assign n_n1004 = ( (~ n_n513) ) ;
 assign n_n1018 = ( (~ n_n520) ) ;
 assign n_n1030 = ( (~ n_n1042) ) ;
 assign n_n1043 = ( (~ n_n1087) ) ;
 assign n_n285 = ( (~ n_n1068) ) ;
 assign n_n1052 = ( (~ n_n1086) ) ;
 assign n_n274 = ( (~ n_n1129) ) ;
 assign n_n267 = ( (~ n_n1138) ) ;
 assign n_n1100 = ( (~ n_n551) ) ;
 assign n_n251 = ( (~ n_n1128) ) ;
 assign n_n243 = ( (~ n_n1242) ) ;
 assign n_n235 = ( (~ n_n1171) ) ;
 assign n_n227 = ( (~ n_n1155) ) ;
 assign n_n220 = ( (~ n_n1153) ) ;
 assign n_n1125 = ( (~ n_n1194) ) ;
 assign n_n1177 = ( (~ n_n570) ) ;
 assign n_n202 = ( (~ n_n1276) ) ;
 assign n_n191 = ( (~ n_n1275) ) ;
 assign n_n169 = ( (~ n_n1226) ) ;
 assign n_n158 = ( (~ n_n1233) ) ;
 assign n_n1202 = ( (~ n_n1315) ) ;
 assign n_n146 = ( (~ n_n1231) ) ;
 assign n_n135 = ( (~ n_n1257) ) ;
 assign n_n124 = ( (~ n_n1333) ) ;
 assign n_n113 = ( (~ n_n1262) ) ;
 assign n_n102 = ( (~ n_n1341) ) ;
 assign n_n77 = ( (~ n_n1362) ) ;
 assign n_n1308 = ( (~ n_n588) ) ;
 assign n_n64 = ( (~ n_n1449) ) ;
 assign n_n56 = ( (~ n_n1451) ) ;
 assign n_n1380 = ( (~ n_n1426) ) ;
 assign n_n52 = ( (~ n_n1401) ) ;
 assign n_n47 = ( (~ n_n1468) ) ;
 assign n_n19 = ( (~ n_n1501) ) ;
 assign n_n1440 = ( (~ n_n618) ) ;
 assign n_n1459 = ( (~ n_n1542) ) ;
 assign n_n1669 = ( (~ n_n1566) ) ;
 assign n_n1509 = ( (~ n_n633) ) ;
 assign n_n700 = ( (~ n_n1719) ) ;
 assign n_n612 = ( n_n30  &  n_n29  &  n_n31 ) ;
 assign n_n607 = ( n_n39  &  n_n38  &  n_n40 ) ;
 assign n_n594 = ( n_n56  &  n_n58  &  n_n59 ) ;
 assign n_n1305 = ( n_n1384  &  n_n1698 ) ;
 assign n_n1292 = ( n_n1387  &  n_n1699 ) ;
 assign n_n1283 = ( n_n1385  &  n_n1701 ) ;
 assign n_n1261 = ( n_n1383  &  n_n1706 ) ;
 assign n_n1217 = ( n_n1381  &  n_n1713 ) ;
 assign n_n1208 = ( n_n120  &  n_n119  &  n_n122  &  n_n121  &  n_n123  &  n_n116  &  n_n118  &  n_n117 ) ;
 assign n_n1188 = ( n_n1316  &  n_n1626  &  n_n1314  &  n_n1315  &  n_n1313 ) ;
 assign n_n572 = ( n_n209  &  n_n208  &  n_n210 ) ;
 assign n_n1165 = ( n_n583  &  n_n1202  &  n_n1695 ) ;
 assign n_n1156 = ( n_n1242  &  n_n1199  &  n_n1696 ) ;
 assign n_n1143 = ( n_n1460  &  n_n1178 ) ;
 assign n_n1134 = ( n_n1652  &  n_n1185 ) ;
 assign n_n553 = ( n_n253  &  n_n252  &  n_n254 ) ;
 assign n_n1082 = ( n_n558  &  n_n1314  &  n_n1694 ) ;
 assign n_n1072 = ( n_n1106  &  n_n562 ) ;
 assign n_n1057 = ( n_n1394  &  n_n1096 ) ;
 assign n_n535 = ( n_n289  &  n_n288  &  n_n290 ) ;
 assign n_n528 = ( n_n1125  &  n_n1077 ) ;
 assign n_n520 = ( n_n1069  &  n_n1038  &  n_n1072  &  n_n1115 ) ;
 assign n_n511 = ( n_n1018  &  n_n1036  &  n_n1015  &  n_n1070 ) ;
 assign n_n503 = ( n_n1027  &  n_n1005 ) ;
 assign n_n936 = ( n_n308  &  n_n307  &  n_n309 ) ;
 assign n_n478 = ( n_n703  &  n_n319 ) ;
 assign n_n909 = ( n_n1396  &  n_n934 ) ;
 assign n_n467 = ( n_n919  &  n_n995 ) ;
 assign n_n459 = ( n_n900  &  n_n895 ) ;
 assign n_n454 = ( n_n884  &  n_n987 ) ;
 assign n_n444 = ( n_n867  &  n_n952 ) ;
 assign n_n436 = ( n_n887  &  n_n865 ) ;
 assign n_n429 = ( n_n479  &  n_n848 ) ;
 assign n_n421 = ( n_n830  &  n_n839 ) ;
 assign n_n413 = ( n_n802  &  n_n844 ) ;
 assign n_n407 = ( n_n343  &  n_n342  &  n_n344 ) ;
 assign n_n384 = ( n_n740  &  n_n735 ) ;
 assign n_n379 = ( n_n367  &  n_n369  &  n_n368  &  n_n370 ) ;
 assign n_n708 = ( (~ n_n374) ) ;
 assign n_n369 = ( (~ n_n720) ) ;
 assign n_n729 = ( (~ n_n384) ) ;
 assign n_n366 = ( (~ n_n753) ) ;
 assign n_n766 = ( (~ n_n778) ) ;
 assign n_n781 = ( (~ n_n787) ) ;
 assign n_n789 = ( (~ n_n409) ) ;
 assign n_n805 = ( (~ n_n417) ) ;
 assign n_n817 = ( (~ n_n423) ) ;
 assign n_n828 = ( (~ n_n842) ) ;
 assign n_n841 = ( (~ n_n865) ) ;
 assign n_n857 = ( (~ n_n444) ) ;
 assign n_n862 = ( (~ n_n448) ) ;
 assign n_n326 = ( (~ n_n928) ) ;
 assign n_n321 = ( (~ n_n914) ) ;
 assign n_n906 = ( (~ n_n472) ) ;
 assign n_n319 = ( (~ n_n955) ) ;
 assign n_n314 = ( (~ n_n960) ) ;
 assign n_n305 = ( (~ n_n957) ) ;
 assign n_n945 = ( (~ n_n970) ) ;
 assign n_n967 = ( (~ n_n492) ) ;
 assign n_n993 = ( (~ n_n503) ) ;
 assign n_n995 = ( (~ n_n505) ) ;
 assign n_n1002 = ( (~ n_n512) ) ;
 assign n_n1019 = ( (~ n_n1074) ) ;
 assign n_n1029 = ( (~ n_n526) ) ;
 assign n_n1044 = ( (~ n_n1088) ) ;
 assign n_n1048 = ( (~ n_n536) ) ;
 assign n_n1053 = ( (~ n_n540) ) ;
 assign n_n275 = ( (~ n_n1130) ) ;
 assign n_n266 = ( (~ n_n1137) ) ;
 assign n_n260 = ( (~ n_n1416) ) ;
 assign n_n259 = ( (~ n_n1147) ) ;
 assign n_n1108 = ( (~ n_n556) ) ;
 assign n_n236 = ( (~ n_n1165) ) ;
 assign n_n1114 = ( (~ n_n562) ) ;
 assign n_n1117 = ( (~ n_n565) ) ;
 assign n_n1126 = ( (~ n_n1308) ) ;
 assign n_n211 = ( (~ n_n1481) ) ;
 assign n_n201 = ( (~ n_n1273) ) ;
 assign n_n192 = ( (~ n_n1274) ) ;
 assign n_n168 = ( (~ n_n1217) ) ;
 assign n_n159 = ( (~ n_n1241) ) ;
 assign n_n1203 = ( (~ n_n1316) ) ;
 assign n_n147 = ( (~ n_n1325) ) ;
 assign n_n134 = ( (~ n_n1265) ) ;
 assign n_n125 = ( (~ n_n1327) ) ;
 assign n_n112 = ( (~ n_n1322) ) ;
 assign n_n103 = ( (~ n_n1336) ) ;
 assign n_n1237 = ( (~ n_n579) ) ;
 assign n_n71 = ( (~ n_n1433) ) ;
 assign n_n65 = ( (~ n_n1439) ) ;
 assign n_n55 = ( (~ n_n1354) ) ;
 assign n_n1377 = ( (~ n_n1422) ) ;
 assign n_n51 = ( (~ n_n1520) ) ;
 assign n_n48 = ( (~ n_n1480) ) ;
 assign n_n18 = ( (~ n_n1591) ) ;
 assign n_n11 = ( (~ n_n1523) ) ;
 assign n_n1460 = ( (~ n_n1547) ) ;
 assign n_n1479 = ( (~ n_n623) ) ;
 assign n_n1510 = ( (~ n_n634) ) ;
 assign n_n1532 = ( (~ n_n643) ) ;
 assign n_n1545 = ( n_n1611  &  n_n688 ) ;
 assign n_n1433 = ( n_n1690  &  n_n1552  &  n_n1453 ) ;
 assign n_n608 = ( n_n36  &  n_n35  &  n_n37 ) ;
 assign n_n1317 = ( n_n1384  &  n_n1681 ) ;
 assign n_n586 = ( n_n1390  &  n_n1515 ) ;
 assign n_n1291 = ( n_n1388  &  n_n1699 ) ;
 assign n_n1273 = ( n_n1386  &  n_n1703 ) ;
 assign n_n1262 = ( n_n1388  &  n_n1706 ) ;
 assign n_n1220 = ( n_n1388  &  n_n1713 ) ;
 assign n_n1209 = ( n_n112  &  n_n111  &  n_n114  &  n_n113  &  n_n115  &  n_n108  &  n_n110  &  n_n109 ) ;
 assign n_n1187 = ( n_n144  &  n_n159  &  n_n114  &  n_n129  &  n_n160  &  n_n156  &  n_n158  &  n_n157 ) ;
 assign n_n569 = ( n_n1229  &  n_n1237 ) ;
 assign n_n1168 = ( n_n578  &  n_n1311  &  n_n1694 ) ;
 assign n_n1157 = ( n_n1247  &  n_n1200  &  n_n1696 ) ;
 assign n_n565 = ( n_n221  &  n_n222 ) ;
 assign n_n554 = ( n_n250  &  n_n249  &  n_n251 ) ;
 assign n_n1081 = ( n_n554  &  n_n1310  &  n_n1694 ) ;
 assign n_n1068 = ( n_n1110  &  n_n1314  &  n_n1697 ) ;
 assign n_n1060 = ( n_n1394  &  n_n1099 ) ;
 assign n_n536 = ( n_n286  &  n_n287 ) ;
 assign n_n527 = ( n_n1124  &  n_n1078 ) ;
 assign n_n1011 = ( n_n1399  &  n_n1034 ) ;
 assign n_n513 = ( n_n1013  &  n_n1189 ) ;
 assign n_n504 = ( n_n1028  &  n_n1006 ) ;
 assign n_n961 = ( n_n1459  &  n_n979 ) ;
 assign n_n489 = ( n_n1089  &  n_n970 ) ;
 assign n_n908 = ( n_n1396  &  n_n933 ) ;
 assign n_n464 = ( n_n922  &  n_n964 ) ;
 assign n_n462 = ( n_n975  &  n_n902 ) ;
 assign n_n873 = ( n_n1452  &  n_n906 ) ;
 assign n_n860 = ( n_n331  &  n_n332 ) ;
 assign n_n437 = ( n_n871  &  n_n857 ) ;
 assign n_n826 = ( n_n1452  &  n_n844 ) ;
 assign n_n420 = ( n_n819  &  n_n813 ) ;
 assign n_n801 = ( n_n825  &  n_n825 ) ;
 assign n_n408 = ( n_n803  &  n_n793 ) ;
 assign n_n387 = ( n_n738  &  n_n746 ) ;
 assign n_n380 = ( n_n727  &  n_n733 ) ;
 assign n_n709 = ( (~ n_n375) ) ;
 assign n_n716 = ( (~ n_n379) ) ;
 assign n_n727 = ( (~ n_n732) ) ;
 assign n_n738 = ( (~ n_n390) ) ;
 assign n_n355 = ( (~ n_n780) ) ;
 assign n_n347 = ( (~ n_n785) ) ;
 assign n_n340 = ( (~ n_n806) ) ;
 assign n_n807 = ( (~ n_n418) ) ;
 assign n_n820 = ( (~ n_n831) ) ;
 assign n_n825 = ( (~ n_n427) ) ;
 assign n_n840 = ( (~ n_n433) ) ;
 assign n_n872 = ( (~ n_n454) ) ;
 assign n_n884 = ( (~ n_n926) ) ;
 assign n_n322 = ( (~ n_n1060) ) ;
 assign n_n916 = ( (~ n_n962) ) ;
 assign n_n925 = ( (~ n_n480) ) ;
 assign n_n317 = ( (~ n_n959) ) ;
 assign n_n306 = ( (~ n_n1059) ) ;
 assign n_n946 = ( (~ n_n486) ) ;
 assign n_n979 = ( (~ n_n993) ) ;
 assign n_n992 = ( (~ n_n502) ) ;
 assign n_n1020 = ( (~ n_n1077) ) ;
 assign n_n1032 = ( (~ n_n528) ) ;
 assign n_n1037 = ( (~ n_n532) ) ;
 assign n_n286 = ( (~ n_n1071) ) ;
 assign n_n277 = ( (~ n_n1102) ) ;
 assign n_n273 = ( (~ n_n1132) ) ;
 assign n_n268 = ( (~ n_n1135) ) ;
 assign n_n261 = ( (~ n_n1143) ) ;
 assign n_n242 = ( (~ n_n1164) ) ;
 assign n_n1111 = ( (~ n_n559) ) ;
 assign n_n1113 = ( (~ n_n561) ) ;
 assign n_n221 = ( (~ n_n1158) ) ;
 assign n_n216 = ( (~ n_n1175) ) ;
 assign n_n210 = ( (~ n_n1214) ) ;
 assign n_n204 = ( (~ n_n1285) ) ;
 assign n_n193 = ( (~ n_n1277) ) ;
 assign n_n167 = ( (~ n_n1303) ) ;
 assign n_n156 = ( (~ n_n1215) ) ;
 assign n_n1200 = ( (~ n_n1313) ) ;
 assign n_n148 = ( (~ n_n1267) ) ;
 assign n_n133 = ( (~ n_n1319) ) ;
 assign n_n122 = ( (~ n_n1248) ) ;
 assign n_n115 = ( (~ n_n1347) ) ;
 assign n_n104 = ( (~ n_n1330) ) ;
 assign n_n83 = ( (~ n_n1364) ) ;
 assign n_n75 = ( (~ n_n1423) ) ;
 assign n_n1311 = ( (~ n_n591) ) ;
 assign n_n1315 = ( (~ n_n595) ) ;
 assign n_n1382 = ( (~ n_n1506) ) ;
 assign n_n1389 = ( (~ n_n1515) ) ;
 assign n_n49 = ( (~ n_n1562) ) ;
 assign n_n33 = ( (~ n_n1527) ) ;
 assign n_n1431 = ( (~ n_n613) ) ;
 assign n_n1461 = ( (~ n_n1548) ) ;
 assign n_n701 = ( (~ n_n1709) ) ;
 assign n_n1507 = ( (~ n_n631) ) ;
 assign n_n1531 = ( (~ n_n642) ) ;
 assign n_n642 = ( n_n1670  &  n_n685 ) ;
 assign n_n614 = ( n_n24  &  n_n23  &  n_n25 ) ;
 assign n_n609 = ( n_n1492  &  n_n1574 ) ;
 assign n_n596 = ( n_n56  &  n_n53  &  n_n54 ) ;
 assign n_n587 = ( n_n1389  &  n_n1518 ) ;
 assign n_n1281 = ( n_n1381  &  n_n1701 ) ;
 assign n_n1272 = ( n_n1384  &  n_n1704 ) ;
 assign n_n1263 = ( n_n1387  &  n_n1706 ) ;
 assign n_n1219 = ( n_n1387  &  n_n1713 ) ;
 assign n_n1210 = ( n_n104  &  n_n103  &  n_n106  &  n_n105  &  n_n107  &  n_n100  &  n_n102  &  n_n101 ) ;
 assign n_n1186 = ( n_n152  &  n_n164  &  n_n122  &  n_n137  &  n_n165  &  n_n161  &  n_n163  &  n_n162 ) ;
 assign n_n570 = ( n_n212  &  n_n211  &  n_n213 ) ;
 assign n_n1167 = ( n_n575  &  n_n1309  &  n_n1694 ) ;
 assign n_n1158 = ( n_n1260  &  n_n1202  &  n_n1696 ) ;
 assign n_n564 = ( n_n223  &  n_n224 ) ;
 assign n_n555 = ( n_n247  &  n_n246  &  n_n248 ) ;
 assign n_n1080 = ( n_n558  &  n_n1201  &  n_n1695 ) ;
 assign n_n1069 = ( n_n1104  &  n_n561 ) ;
 assign n_n1059 = ( n_n1394  &  n_n1098 ) ;
 assign n_n537 = ( n_n284  &  n_n285 ) ;
 assign n_n526 = ( n_n1123  &  n_n1072 ) ;
 assign n_n519 = ( n_n1038  &  n_n1114  &  n_n1069 ) ;
 assign n_n1003 = ( n_n1017  &  n_n1023 ) ;
 assign n_n505 = ( n_n1029  &  n_n1007 ) ;
 assign n_n960 = ( n_n1459  &  n_n983 ) ;
 assign n_n950 = ( n_n966  &  n_n1673 ) ;
 assign n_n907 = ( n_n969  &  n_n927  &  n_n1673 ) ;
 assign n_n465 = ( n_n925  &  n_n923  &  n_n921  &  n_n1026 ) ;
 assign n_n461 = ( n_n326  &  n_n327 ) ;
 assign n_n874 = ( n_n1396  &  n_n891 ) ;
 assign n_n446 = ( n_n334  &  n_n333  &  n_n335 ) ;
 assign n_n849 = ( n_n877  &  n_n877 ) ;
 assign n_n427 = ( n_n337  &  n_n336  &  n_n338 ) ;
 assign n_n812 = ( n_n1452  &  n_n831 ) ;
 assign n_n799 = ( n_n1452  &  n_n821 ) ;
 assign n_n788 = ( n_n860  &  n_n844  &  n_n796  &  n_n831 ) ;
 assign n_n386 = ( n_n737  &  n_n744 ) ;
 assign n_n719 = ( n_n723  &  n_n642  &  n_n727 ) ;
 assign n_n710 = ( (~ n_n376) ) ;
 assign n_n367 = ( (~ n_n719) ) ;
 assign n_n728 = ( (~ n_n733) ) ;
 assign n_n737 = ( (~ n_n389) ) ;
 assign n_n348 = ( (~ n_n824) ) ;
 assign n_n346 = ( (~ n_n874) ) ;
 assign n_n341 = ( (~ n_n795) ) ;
 assign n_n808 = ( (~ n_n419) ) ;
 assign n_n819 = ( (~ n_n844) ) ;
 assign n_n428 = ( (~ n_n860) ) ;
 assign n_n839 = ( (~ n_n432) ) ;
 assign n_n330 = ( (~ n_n1367) ) ;
 assign n_n883 = ( (~ n_n902) ) ;
 assign n_n885 = ( (~ n_n460) ) ;
 assign n_n918 = ( (~ n_n473) ) ;
 assign n_n479 = ( (~ n_n478) ) ;
 assign n_n316 = ( (~ n_n1033) ) ;
 assign n_n307 = ( (~ n_n1368) ) ;
 assign n_n971 = ( (~ n_n494) ) ;
 assign n_n980 = ( (~ n_n994) ) ;
 assign n_n991 = ( (~ n_n501) ) ;
 assign n_n1021 = ( (~ n_n521) ) ;
 assign n_n1031 = ( (~ n_n527) ) ;
 assign n_n1040 = ( (~ n_n1083) ) ;
 assign n_n287 = ( (~ n_n1067) ) ;
 assign n_n276 = ( (~ n_n1400) ) ;
 assign n_n1093 = ( (~ n_n544) ) ;
 assign n_n1096 = ( (~ n_n547) ) ;
 assign n_n1099 = ( (~ n_n550) ) ;
 assign n_n241 = ( (~ n_n1170) ) ;
 assign n_n234 = ( (~ n_n1260) ) ;
 assign n_n228 = ( (~ n_n1149) ) ;
 assign n_n222 = ( (~ n_n1152) ) ;
 assign n_n215 = ( (~ n_n1462) ) ;
 assign n_n1178 = ( (~ n_n571) ) ;
 assign n_n203 = ( (~ n_n1280) ) ;
 assign n_n194 = ( (~ n_n1281) ) ;
 assign n_n166 = ( (~ n_n1296) ) ;
 assign n_n157 = ( (~ n_n1224) ) ;
 assign n_n1201 = ( (~ n_n1314) ) ;
 assign n_n149 = ( (~ n_n1259) ) ;
 assign n_n132 = ( (~ n_n1326) ) ;
 assign n_n123 = ( (~ n_n1343) ) ;
 assign n_n114 = ( (~ n_n1254) ) ;
 assign n_n105 = ( (~ n_n1323) ) ;
 assign n_n82 = ( (~ n_n1483) ) ;
 assign n_n76 = ( (~ n_n1498) ) ;
 assign n_n1307 = ( (~ n_n587) ) ;
 assign n_n54 = ( (~ n_n1448) ) ;
 assign n_n1381 = ( (~ n_n1505) ) ;
 assign n_n1390 = ( (~ n_n1518) ) ;
 assign n_n1404 = ( (~ n_n600) ) ;
 assign n_n32 = ( (~ n_n1490) ) ;
 assign n_n26 = ( (~ n_n1514) ) ;
 assign n_n1462 = ( (~ n_n1549) ) ;
 assign n_n1484 = ( (~ n_n624) ) ;
 assign n_n1508 = ( (~ n_n632) ) ;
 assign n_n1526 = ( (~ n_n641) ) ;
 assign n_n649 = ( n_n1716  &  n_n1607 ) ;
 assign n_n643 = ( n_n1718  &  n_n1625  &  n_n1719 ) ;
 assign n_n1435 = ( n_n1689  &  n_n1552  &  n_n1453 ) ;
 assign n_n1423 = ( n_n1604  &  n_n1454  &  n_n1707 ) ;
 assign n_n1319 = ( n_n1386  &  n_n1681 ) ;
 assign n_n588 = ( n_n1392  &  n_n1393 ) ;
 assign n_n582 = ( n_n1380  &  n_n1417 ) ;
 assign n_n580 = ( n_n82  &  n_n81  &  n_n83 ) ;
 assign n_n1231 = ( n_n1383  &  n_n1711 ) ;
 assign n_n1185 = ( n_n170  &  n_n169  &  n_n130  &  n_n145  &  n_n171  &  n_n166  &  n_n168  &  n_n167 ) ;
 assign n_n1174 = ( n_n1538  &  n_n1230 ) ;
 assign n_n1148 = ( n_n1222  &  n_n1309  &  n_n1697 ) ;
 assign n_n1137 = ( n_n1716  &  n_n1207 ) ;
 assign n_n567 = ( n_n217  &  n_n218 ) ;
 assign n_n556 = ( n_n244  &  n_n243  &  n_n245 ) ;
 assign n_n1079 = ( n_n554  &  n_n1197  &  n_n1695 ) ;
 assign n_n541 = ( n_n1107  &  n_n1178 ) ;
 assign n_n1054 = ( n_n1394  &  n_n1093 ) ;
 assign n_n1041 = ( n_n1581  &  n_n1048 ) ;
 assign n_n532 = ( n_n1049  &  n_n1074 ) ;
 assign n_n522 = ( n_n1074  &  n_n1039  &  n_n1077  &  n_n1118 ) ;
 assign n_n515 = ( n_n1016  &  n_n1191 ) ;
 assign n_n506 = ( n_n294  &  n_n295 ) ;
 assign n_n959 = ( n_n1459  &  n_n982 ) ;
 assign n_n487 = ( n_n983  &  n_n1088 ) ;
 assign n_n933 = ( n_n317  &  n_n316  &  n_n318 ) ;
 assign n_n473 = ( n_n949  &  n_n948  &  n_n1030 ) ;
 assign n_n889 = ( n_n962  &  n_n894  &  n_n1673 ) ;
 assign n_n875 = ( n_n1396  &  n_n892 ) ;
 assign n_n441 = ( n_n866  &  n_n950 ) ;
 assign n_n433 = ( n_n863  &  n_n852 ) ;
 assign n_n837 = ( n_n1452  &  n_n856 ) ;
 assign n_n424 = ( n_n868  &  n_n840 ) ;
 assign n_n416 = ( n_n822  &  n_n842 ) ;
 assign n_n409 = ( n_n340  &  n_n341 ) ;
 assign n_n724 = ( n_n729  &  n_n642  &  n_n732 ) ;
 assign n_n374 = ( n_n712  &  n_n717 ) ;
 assign n_n705 = ( n_n707  &  n_n707 ) ;
 assign n_n714 = ( (~ n_n717) ) ;
 assign n_n723 = ( (~ n_n729) ) ;
 assign n_n736 = ( (~ n_n748) ) ;
 assign n_n343 = ( (~ n_n1212) ) ;
 assign n_n339 = ( (~ n_n811) ) ;
 assign n_n798 = ( (~ n_n414) ) ;
 assign n_n814 = ( (~ n_n421) ) ;
 assign n_n337 = ( (~ n_n838) ) ;
 assign n_n834 = ( (~ n_n859) ) ;
 assign n_n887 = ( (~ n_n930) ) ;
 assign n_n897 = ( (~ n_n466) ) ;
 assign n_n922 = ( (~ n_n942) ) ;
 assign n_n932 = ( (~ n_n482) ) ;
 assign n_n308 = ( (~ n_n958) ) ;
 assign n_n996 = ( (~ n_n506) ) ;
 assign n_n1009 = ( (~ n_n517) ) ;
 assign n_n1035 = ( (~ n_n530) ) ;
 assign n_n1047 = ( (~ n_n535) ) ;
 assign n_n256 = ( (~ n_n1144) ) ;
 assign n_n248 = ( (~ n_n1162) ) ;
 assign n_n1116 = ( (~ n_n564) ) ;
 assign n_n214 = ( (~ n_n1413) ) ;
 assign n_n187 = ( (~ n_n1287) ) ;
 assign n_n176 = ( (~ n_n1227) ) ;
 assign n_n131 = ( (~ n_n1338) ) ;
 assign n_n120 = ( (~ n_n1263) ) ;
 assign n_n98 = ( (~ n_n1324) ) ;
 assign n_n1229 = ( (~ n_n576) ) ;
 assign n_n53 = ( (~ n_n1353) ) ;
 assign n_n1384 = ( (~ n_n1508) ) ;
 assign n_n1392 = ( (~ n_n598) ) ;
 assign n_n44 = ( (~ n_n1503) ) ;
 assign n_n38 = ( (~ n_n1485) ) ;
 assign n_n1465 = ( (~ n_n1551) ) ;
 assign n_n1492 = ( (~ n_n626) ) ;
 assign n_n1515 = ( (~ n_n637) ) ;
 assign n_n1537 = ( (~ n_n645) ) ;
 assign n_n1656 = ( (~ n_n1711) ) ;
 assign n_n1546 = ( n_n1611  &  n_n1649 ) ;
 assign n_n1533 = ( n_n1617  &  n_n1719 ) ;
 assign n_n615 = ( n_n21  &  n_n20  &  n_n22 ) ;
 assign n_n1424 = ( n_n1463  &  n_n693 ) ;
 assign n_n1318 = ( n_n1385  &  n_n1681 ) ;
 assign n_n589 = ( n_n64  &  n_n70  &  n_n71 ) ;
 assign n_n1252 = ( n_n1381  &  n_n1708 ) ;
 assign n_n1243 = ( n_n1383  &  n_n1709 ) ;
 assign n_n1221 = ( n_n1383  &  n_n1713 ) ;
 assign n_n1184 = ( n_n176  &  n_n175  &  n_n138  &  n_n153  &  n_n177  &  n_n172  &  n_n174  &  n_n173 ) ;
 assign n_n1175 = ( n_n1460  &  n_n1308 ) ;
 assign n_n1147 = ( n_n1555  &  n_n1176 ) ;
 assign n_n1138 = ( n_n1652  &  n_n1183 ) ;
 assign n_n566 = ( n_n219  &  n_n220 ) ;
 assign n_n557 = ( n_n241  &  n_n240  &  n_n242 ) ;
 assign n_n1078 = ( n_n1112  &  n_n566 ) ;
 assign n_n1067 = ( n_n1105  &  n_n1310  &  n_n1697 ) ;
 assign n_n540 = ( n_n1090  &  n_n1091 ) ;
 assign n_n1042 = ( n_n1583  &  n_n1049 ) ;
 assign n_n531 = ( n_n1048  &  n_n1069 ) ;
 assign n_n523 = ( n_n1120  &  n_n1069 ) ;
 assign n_n514 = ( n_n1019  &  n_n1190 ) ;
 assign n_n507 = ( n_n1031  &  n_n1009 ) ;
 assign n_n958 = ( n_n1455  &  n_n978 ) ;
 assign n_n488 = ( n_n998  &  n_n1088  &  n_n970 ) ;
 assign n_n482 = ( n_n943  &  n_n1673 ) ;
 assign n_n474 = ( n_n981  &  n_n941 ) ;
 assign n_n463 = ( n_n953  &  n_n926 ) ;
 assign n_n876 = ( n_n1398  &  n_n906 ) ;
 assign n_n440 = ( n_n864  &  n_n992 ) ;
 assign n_n842 = ( n_n478  &  n_n858 ) ;
 assign n_n836 = ( n_n1452  &  n_n858 ) ;
 assign n_n425 = ( n_n846  &  n_n832 ) ;
 assign n_n415 = ( n_n428  &  n_n820 ) ;
 assign n_n410 = ( n_n797  &  n_n809 ) ;
 assign n_n382 = ( n_n728  &  n_n732 ) ;
 assign n_n375 = ( n_n711  &  n_n721 ) ;
 assign n_n371 = ( n_n706  &  n_n706 ) ;
 assign n_n713 = ( (~ n_n377) ) ;
 assign n_n726 = ( (~ n_n383) ) ;
 assign n_n735 = ( (~ n_n388) ) ;
 assign n_n342 = ( (~ n_n792) ) ;
 assign n_n794 = ( (~ n_n805) ) ;
 assign n_n800 = ( (~ n_n825) ) ;
 assign n_n811 = ( (~ n_n821) ) ;
 assign n_n336 = ( (~ n_n911) ) ;
 assign n_n833 = ( (~ n_n848) ) ;
 assign n_n888 = ( (~ n_n463) ) ;
 assign n_n896 = ( (~ n_n465) ) ;
 assign n_n901 = ( (~ n_n469) ) ;
 assign n_n318 = ( (~ n_n1054) ) ;
 assign n_n309 = ( (~ n_n1061) ) ;
 assign n_n997 = ( (~ n_n507) ) ;
 assign n_n1007 = ( (~ n_n516) ) ;
 assign n_n1036 = ( (~ n_n531) ) ;
 assign n_n288 = ( (~ n_n1424) ) ;
 assign n_n255 = ( (~ n_n1402) ) ;
 assign n_n1105 = ( (~ n_n554) ) ;
 assign n_n229 = ( (~ n_n1154) ) ;
 assign n_n209 = ( (~ n_n1477) ) ;
 assign n_n186 = ( (~ n_n1282) ) ;
 assign n_n177 = ( (~ n_n1284) ) ;
 assign n_n130 = ( (~ n_n1243) ) ;
 assign n_n121 = ( (~ n_n1255) ) ;
 assign n_n97 = ( (~ n_n1331) ) ;
 assign n_n1222 = ( (~ n_n575) ) ;
 assign n_n1316 = ( (~ n_n596) ) ;
 assign n_n1383 = ( (~ n_n1507) ) ;
 assign n_n45 = ( (~ n_n1472) ) ;
 assign n_n1407 = ( (~ n_n602) ) ;
 assign n_n39 = ( (~ n_n1500) ) ;
 assign n_n1467 = ( (~ n_n620) ) ;
 assign n_n1489 = ( (~ n_n625) ) ;
 assign n_n1518 = ( (~ n_n638) ) ;
 assign n_n1536 = ( (~ n_n1602) ) ;
 assign n_n651 = ( n_n1652  &  n_n1607 ) ;
 assign n_n644 = ( n_n6  &  n_n700 ) ;
 assign n_n1437 = ( n_n1688  &  n_n1552  &  n_n1453 ) ;
 assign n_n1425 = ( n_n1462  &  n_n1576 ) ;
 assign n_n590 = ( n_n64  &  n_n68  &  n_n69 ) ;
 assign n_n1251 = ( n_n1382  &  n_n1708 ) ;
 assign n_n1233 = ( n_n1381  &  n_n1711 ) ;
 assign n_n575 = ( n_n90  &  n_n89  &  n_n91 ) ;
 assign n_n1164 = ( n_n581  &  n_n1200  &  n_n1695 ) ;
 assign n_n1153 = ( n_n1269  &  n_n1316  &  n_n1697 ) ;
 assign n_n1146 = ( n_n1465  &  n_n1180 ) ;
 assign n_n1135 = ( n_n1716  &  n_n1208 ) ;
 assign n_n1128 = ( n_n1536  &  n_n1179 ) ;
 assign n_n558 = ( n_n238  &  n_n237  &  n_n239 ) ;
 assign n_n1077 = ( n_n1111  &  n_n565 ) ;
 assign n_n1063 = ( n_n1460  &  n_n1101 ) ;
 assign n_n1056 = ( n_n1394  &  n_n1095 ) ;
 assign n_n533 = ( n_n1053  &  n_n1053 ) ;
 assign n_n530 = ( n_n1046  &  n_n1066 ) ;
 assign n_n521 = ( n_n1039  &  n_n1117  &  n_n1074 ) ;
 assign n_n1008 = ( n_n1583  &  n_n1023 ) ;
 assign n_n508 = ( n_n1032  &  n_n1010 ) ;
 assign n_n957 = ( n_n1455  &  n_n981 ) ;
 assign n_n944 = ( n_n998  &  n_n970  &  n_n997 ) ;
 assign n_n935 = ( n_n311  &  n_n310  &  n_n312 ) ;
 assign n_n475 = ( n_n995  &  n_n1085  &  n_n964 ) ;
 assign n_n912 = ( n_n1396  &  n_n937 ) ;
 assign n_n468 = ( n_n940  &  n_n942 ) ;
 assign n_n443 = ( n_n886  &  n_n870 ) ;
 assign n_n843 = ( n_n851  &  n_n1673 ) ;
 assign n_n835 = ( n_n859  &  n_n859 ) ;
 assign n_n422 = ( n_n833  &  n_n478 ) ;
 assign n_n806 = ( n_n478  &  n_n847  &  n_n821  &  n_n858 ) ;
 assign n_n792 = ( n_n1456  &  n_n807 ) ;
 assign n_n383 = ( n_n730  &  n_n748 ) ;
 assign n_n376 = ( n_n717  &  n_n715 ) ;
 assign n_n1662 = ( (~ n_n371) ) ;
 assign n_n370 = ( (~ n_n724) ) ;
 assign n_n721 = ( (~ n_n381) ) ;
 assign n_n733 = ( (~ n_n387) ) ;
 assign n_n345 = ( (~ n_n790) ) ;
 assign n_n793 = ( (~ n_n411) ) ;
 assign n_n802 = ( (~ n_n813) ) ;
 assign n_n816 = ( (~ n_n422) ) ;
 assign n_n823 = ( (~ n_n426) ) ;
 assign n_n832 = ( (~ n_n431) ) ;
 assign n_n1664 = ( (~ n_n461) ) ;
 assign n_n895 = ( (~ n_n464) ) ;
 assign n_n902 = ( (~ n_n470) ) ;
 assign n_n924 = ( (~ n_n477) ) ;
 assign n_n310 = ( (~ n_n1092) ) ;
 assign n_n295 = ( (~ n_n1084) ) ;
 assign n_n1006 = ( (~ n_n515) ) ;
 assign n_n1015 = ( (~ n_n519) ) ;
 assign n_n1028 = ( (~ n_n525) ) ;
 assign n_n258 = ( (~ n_n1466) ) ;
 assign n_n249 = ( (~ n_n1405) ) ;
 assign n_n1110 = ( (~ n_n558) ) ;
 assign n_n200 = ( (~ n_n1271) ) ;
 assign n_n189 = ( (~ n_n1300) ) ;
 assign n_n178 = ( (~ n_n1283) ) ;
 assign n_n111 = ( (~ n_n1329) ) ;
 assign n_n100 = ( (~ n_n1348) ) ;
 assign n_n89 = ( (~ n_n1403) ) ;
 assign n_n1370 = ( (~ n_n1404) ) ;
 assign n_n50 = ( (~ n_n1446) ) ;
 assign n_n46 = ( (~ n_n1563) ) ;
 assign n_n702 = ( (~ n_n1713) ) ;
 assign n_n1499 = ( (~ n_n628) ) ;
 assign n_n1511 = ( (~ n_n635) ) ;
 assign n_n1534 = ( (~ n_n644) ) ;
 assign n_n650 = ( n_n697  &  n_n1716 ) ;
 assign n_n1535 = ( n_n1718  &  n_n1612  &  n_n1719 ) ;
 assign n_n616 = ( n_n18  &  n_n17  &  n_n19 ) ;
 assign n_n610 = ( n_n1495  &  n_n1499 ) ;
 assign n_n1320 = ( n_n1381  &  n_n1681 ) ;
 assign n_n1241 = ( n_n1382  &  n_n1710 ) ;
 assign n_n1232 = ( n_n1388  &  n_n1711 ) ;
 assign n_n1223 = ( n_n1383  &  n_n1712 ) ;
 assign n_n1163 = ( n_n580  &  n_n1199  &  n_n1695 ) ;
 assign n_n1154 = ( n_n1222  &  n_n1196  &  n_n1696 ) ;
 assign n_n568 = ( n_n215  &  n_n214  &  n_n216 ) ;
 assign n_n1136 = ( n_n1652  &  n_n1184 ) ;
 assign n_n1127 = ( n_n1536  &  n_n1177 ) ;
 assign n_n559 = ( n_n235  &  n_n234  &  n_n236 ) ;
 assign n_n1076 = ( n_n1110  &  n_n1201  &  n_n1696 ) ;
 assign n_n1064 = ( n_n276  &  n_n277 ) ;
 assign n_n1055 = ( n_n1394  &  n_n1094 ) ;
 assign n_n1045 = ( n_n1460  &  n_n1064 ) ;
 assign n_n529 = ( n_n292  &  n_n291  &  n_n293 ) ;
 assign n_n1023 = ( n_n1078  &  n_n1039  &  n_n1077  &  n_n1074 ) ;
 assign n_n516 = ( n_n1014  &  n_n1192 ) ;
 assign n_n509 = ( n_n1043  &  n_n1039 ) ;
 assign n_n956 = ( n_n1455  &  n_n980 ) ;
 assign n_n486 = ( n_n703  &  n_n994 ) ;
 assign n_n934 = ( n_n314  &  n_n313  &  n_n315 ) ;
 assign n_n476 = ( n_n1086  &  n_n964 ) ;
 assign n_n911 = ( n_n1396  &  n_n938 ) ;
 assign n_n469 = ( n_n927  &  n_n970 ) ;
 assign n_n442 = ( n_n905  &  n_n881 ) ;
 assign n_n434 = ( n_n869  &  n_n854 ) ;
 assign n_n431 = ( n_n841  &  n_n930 ) ;
 assign n_n423 = ( n_n827  &  n_n843 ) ;
 assign n_n417 = ( n_n829  &  n_n816 ) ;
 assign n_n411 = ( n_n810  &  n_n860 ) ;
 assign n_n725 = ( n_n729  &  n_n1531  &  n_n727 ) ;
 assign n_n377 = ( n_n714  &  n_n716 ) ;
 assign n_n706 = ( (~ n_n372) ) ;
 assign n_n715 = ( (~ n_n378) ) ;
 assign n_n722 = ( (~ n_n382) ) ;
 assign n_n732 = ( (~ n_n386) ) ;
 assign n_n344 = ( (~ n_n1174) ) ;
 assign n_n791 = ( (~ n_n410) ) ;
 assign n_n803 = ( (~ n_n415) ) ;
 assign n_n815 = ( (~ n_n840) ) ;
 assign n_n338 = ( (~ n_n837) ) ;
 assign n_n831 = ( (~ n_n430) ) ;
 assign n_n886 = ( (~ n_n462) ) ;
 assign n_n894 = ( (~ n_n939) ) ;
 assign n_n903 = ( (~ n_n471) ) ;
 assign n_n923 = ( (~ n_n476) ) ;
 assign n_n931 = ( (~ n_n952) ) ;
 assign n_n294 = ( (~ n_n1008) ) ;
 assign n_n1005 = ( (~ n_n514) ) ;
 assign n_n1016 = ( (~ n_n1073) ) ;
 assign n_n1027 = ( (~ n_n524) ) ;
 assign n_n257 = ( (~ n_n1146) ) ;
 assign n_n250 = ( (~ n_n1474) ) ;
 assign n_n244 = ( (~ n_n1169) ) ;
 assign n_n190 = ( (~ n_n1220) ) ;
 assign n_n188 = ( (~ n_n1293) ) ;
 assign n_n179 = ( (~ n_n1288) ) ;
 assign n_n110 = ( (~ n_n1335) ) ;
 assign n_n101 = ( (~ n_n1345) ) ;
 assign n_n99 = ( (~ n_n1352) ) ;
 assign n_n1385 = ( (~ n_n1509) ) ;
 assign n_n1391 = ( (~ n_n597) ) ;
 assign n_n1406 = ( (~ n_n601) ) ;
 assign n_n7 = ( (~ n_n1534) ) ;
 assign n_n1495 = ( (~ n_n627) ) ;
 assign n_n1512 = ( (~ n_n636) ) ;
 assign n_n6 = ( (~ n_n1605) ) ;
 assign n_n685 = ( n_n1  &  n_n2 ) ;
 assign n_n640 = ( n_n1600  &  n_n1592 ) ;
 assign n_n1514 = ( n_n1550  &  n_n1690 ) ;
 assign n_n1503 = ( n_n1543  &  n_n1699 ) ;
 assign n_n626 = ( n_n1658  &  n_n1708 ) ;
 assign n_n1481 = ( n_n1543  &  n_n1710 ) ;
 assign n_n1416 = ( n_n1463  &  n_n1657 ) ;
 assign n_n1405 = ( n_n1603  &  n_n1454  &  n_n1712 ) ;
 assign n_n598 = ( n_n1447  &  n_n1522 ) ;
 assign n_n1365 = ( n_n1536  &  n_n1406 ) ;
 assign n_n1354 = ( n_n1440  &  n_n1535 ) ;
 assign n_n1343 = ( n_n1384  &  n_n1677 ) ;
 assign n_n1332 = ( n_n1384  &  n_n1679 ) ;
 assign n_n1321 = ( n_n1382  &  n_n1681 ) ;
 assign n_n1290 = ( n_n1384  &  n_n1700 ) ;
 assign n_n1279 = ( n_n1384  &  n_n1702 ) ;
 assign n_n584 = ( n_n1376  &  n_n1426 ) ;
 assign n_n1257 = ( n_n1382  &  n_n1707 ) ;
 assign n_n1246 = ( n_n1382  &  n_n1709 ) ;
 assign n_n1235 = ( n_n1387  &  n_n1711 ) ;
 assign n_n1224 = ( n_n1386  &  n_n1712 ) ;
 assign n_n1152 = ( n_n1260  &  n_n1315  &  n_n1697 ) ;
 assign n_n1141 = ( n_n1716  &  n_n1205 ) ;
 assign n_n1130 = ( n_n1652  &  n_n1187 ) ;
 assign n_n560 = ( n_n232  &  n_n231  &  n_n233 ) ;
 assign n_n548 = ( n_n266  &  n_n267 ) ;
 assign n_n1086 = ( n_n1583  &  n_n1114 ) ;
 assign n_n1000 = ( n_n1583  &  n_n1002 ) ;
 assign n_n498 = ( n_n990  &  n_n1087 ) ;
 assign n_n966 = ( n_n994  &  n_n995  &  n_n996 ) ;
 assign n_n782 = ( n_n428  &  n_n345 ) ;
 assign n_n770 = ( n_n1398  &  n_n776 ) ;
 assign n_n755 = ( n_n761  &  n_n1644 ) ;
 assign n_n391 = ( n_n754  &  n_n755 ) ;
 assign n_n743 = ( (~ n_n392) ) ;
 assign n_n760 = ( (~ n_n773) ) ;
 assign n_n768 = ( (~ n_n401) ) ;
 assign n_n776 = ( (~ n_n404) ) ;
 assign n_n847 = ( (~ n_n437) ) ;
 assign n_n335 = ( (~ n_n873) ) ;
 assign n_n866 = ( (~ n_n882) ) ;
 assign n_n878 = ( (~ n_n456) ) ;
 assign n_n323 = ( (~ n_n1062) ) ;
 assign n_n947 = ( (~ n_n487) ) ;
 assign n_n297 = ( (~ n_n1089) ) ;
 assign n_n984 = ( (~ n_n498) ) ;
 assign n_n1666 = ( (~ n_n510) ) ;
 assign n_n1014 = ( (~ n_n1072) ) ;
 assign n_n272 = ( (~ n_n1131) ) ;
 assign n_n265 = ( (~ n_n1140) ) ;
 assign n_n253 = ( (~ n_n1167) ) ;
 assign n_n1107 = ( (~ n_n1176) ) ;
 assign n_n237 = ( (~ n_n1418) ) ;
 assign n_n199 = ( (~ n_n1272) ) ;
 assign n_n183 = ( (~ n_n1228) ) ;
 assign n_n172 = ( (~ n_n1289) ) ;
 assign n_n161 = ( (~ n_n1304) ) ;
 assign n_n1199 = ( (~ n_n1312) ) ;
 assign n_n94 = ( (~ n_n1346) ) ;
 assign n_n86 = ( (~ n_n1365) ) ;
 assign n_n78 = ( (~ n_n1415) ) ;
 assign n_n1269 = ( (~ n_n585) ) ;
 assign n_n66 = ( (~ n_n1358) ) ;
 assign n_n43 = ( (~ n_n1567) ) ;
 assign n_n35 = ( (~ n_n1476) ) ;
 assign n_n29 = ( (~ n_n1513) ) ;
 assign n_n21 = ( (~ n_n1589) ) ;
 assign n_n13 = ( (~ n_n1529) ) ;
 assign n_n1453 = ( (~ n_n1535) ) ;
 assign n_n693 = ( (~ n_n1706) ) ;
 assign n_n686 = ( n_n1718  &  n_n1719 ) ;
 assign n_n1524 = ( n_n1550  &  n_n1684 ) ;
 assign n_n637 = ( n_n1586  &  n_n1588 ) ;
 assign n_n1502 = ( n_n7  &  n_n693 ) ;
 assign n_n1493 = ( n_n699  &  n_n1708 ) ;
 assign n_n1471 = ( n_n1543  &  n_n1712 ) ;
 assign n_n1415 = ( n_n1604  &  n_n1454  &  n_n1709 ) ;
 assign n_n601 = ( n_n48  &  n_n47  &  n_n49 ) ;
 assign n_n597 = ( n_n51  &  n_n50  &  n_n52 ) ;
 assign n_n1366 = ( n_n1536  &  n_n1407 ) ;
 assign n_n1353 = ( n_n1443  &  n_n1535 ) ;
 assign n_n1344 = ( n_n1385  &  n_n1677 ) ;
 assign n_n1331 = ( n_n1388  &  n_n1680 ) ;
 assign n_n1322 = ( n_n1387  &  n_n1681 ) ;
 assign n_n1300 = ( n_n1387  &  n_n1698 ) ;
 assign n_n1278 = ( n_n1385  &  n_n1702 ) ;
 assign n_n585 = ( n_n73  &  n_n72  &  n_n74 ) ;
 assign n_n1256 = ( n_n1387  &  n_n1707 ) ;
 assign n_n581 = ( n_n79  &  n_n78  &  n_n80 ) ;
 assign n_n1234 = ( n_n1382  &  n_n1711 ) ;
 assign n_n1225 = ( n_n1381  &  n_n1712 ) ;
 assign n_n1151 = ( n_n1247  &  n_n1313  &  n_n1697 ) ;
 assign n_n1142 = ( n_n1652  &  n_n1181 ) ;
 assign n_n1129 = ( n_n1716  &  n_n1211 ) ;
 assign n_n561 = ( n_n229  &  n_n230 ) ;
 assign n_n547 = ( n_n268  &  n_n269 ) ;
 assign n_n1087 = ( n_n1110  &  n_n1582 ) ;
 assign n_n517 = ( n_n1022  &  n_n1193 ) ;
 assign n_n497 = ( n_n989  &  n_n1083 ) ;
 assign n_n492 = ( n_n1085  &  n_n995 ) ;
 assign n_n780 = ( n_n1398  &  n_n791 ) ;
 assign n_n771 = ( n_n1644  &  n_n773 ) ;
 assign n_n753 = ( n_n399  &  n_n685  &  n_n403 ) ;
 assign n_n742 = ( n_n750  &  n_n762 ) ;
 assign n_n744 = ( (~ n_n393) ) ;
 assign n_n758 = ( (~ n_n398) ) ;
 assign n_n359 = ( (~ n_n799) ) ;
 assign n_n352 = ( (~ n_n788) ) ;
 assign n_n848 = ( (~ n_n858) ) ;
 assign n_n858 = ( (~ n_n445) ) ;
 assign n_n867 = ( (~ n_n885) ) ;
 assign n_n877 = ( (~ n_n455) ) ;
 assign n_n900 = ( (~ n_n468) ) ;
 assign n_n300 = ( (~ n_n963) ) ;
 assign n_n296 = ( (~ n_n985) ) ;
 assign n_n983 = ( (~ n_n998) ) ;
 assign n_n1001 = ( (~ n_n511) ) ;
 assign n_n1013 = ( (~ n_n1069) ) ;
 assign n_n1094 = ( (~ n_n545) ) ;
 assign n_n1097 = ( (~ n_n548) ) ;
 assign n_n252 = ( (~ n_n1222) ) ;
 assign n_n1106 = ( (~ n_n555) ) ;
 assign n_n230 = ( (~ n_n1148) ) ;
 assign n_n208 = ( (~ n_n1504) ) ;
 assign n_n182 = ( (~ n_n1219) ) ;
 assign n_n173 = ( (~ n_n1295) ) ;
 assign n_n160 = ( (~ n_n1305) ) ;
 assign n_n1198 = ( (~ n_n1311) ) ;
 assign n_n93 = ( (~ n_n1349) ) ;
 assign n_n1230 = ( (~ n_n577) ) ;
 assign n_n1247 = ( (~ n_n581) ) ;
 assign n_n72 = ( (~ n_n1428) ) ;
 assign n_n59 = ( (~ n_n1444) ) ;
 assign n_n42 = ( (~ n_n1486) ) ;
 assign n_n36 = ( (~ n_n1491) ) ;
 assign n_n1430 = ( (~ n_n612) ) ;
 assign n_n22 = ( (~ n_n1497) ) ;
 assign n_n12 = ( (~ n_n1596) ) ;
 assign n_n1452 = ( (~ n_n1533) ) ;
 assign n_n1658 = ( (~ n_n1707) ) ;
 assign n_n677 = ( n_n1713  &  n_n1690 ) ;
 assign n_n1614 = ( n_n1654  &  n_n700 ) ;
 assign n_n1523 = ( n_n1550  &  n_n1685 ) ;
 assign n_n636 = ( n_n1546  &  n_n1627 ) ;
 assign n_n629 = ( n_n1579  &  n_n676 ) ;
 assign n_n1494 = ( n_n7  &  n_n1657 ) ;
 assign n_n1454 = ( n_n1534  &  n_n1602 ) ;
 assign n_n1414 = ( n_n1462  &  n_n1569 ) ;
 assign n_n1403 = ( n_n1603  &  n_n1454  &  n_n1713 ) ;
 assign n_n1395 = ( n_n1719  &  n_n1539 ) ;
 assign n_n1367 = ( n_n1398  &  n_n1556 ) ;
 assign n_n1352 = ( n_n1384  &  n_n1674 ) ;
 assign n_n1341 = ( n_n1381  &  n_n1678 ) ;
 assign n_n1334 = ( n_n1386  &  n_n1679 ) ;
 assign n_n1323 = ( n_n1388  &  n_n1681 ) ;
 assign n_n1299 = ( n_n1388  &  n_n1698 ) ;
 assign n_n1288 = ( n_n1386  &  n_n1700 ) ;
 assign n_n1270 = ( n_n1384  &  n_n1705 ) ;
 assign n_n1255 = ( n_n1388  &  n_n1707 ) ;
 assign n_n1244 = ( n_n1388  &  n_n1709 ) ;
 assign n_n579 = ( n_n1370  &  n_n1410 ) ;
 assign n_n1226 = ( n_n1382  &  n_n1712 ) ;
 assign n_n1212 = ( n_n1458  &  n_n1378 ) ;
 assign n_n1194 = ( n_n1260  &  n_n1582 ) ;
 assign n_n1150 = ( n_n1242  &  n_n1312  &  n_n1697 ) ;
 assign n_n1139 = ( n_n1716  &  n_n1206 ) ;
 assign n_n1132 = ( n_n1652  &  n_n1186 ) ;
 assign n_n562 = ( n_n227  &  n_n228 ) ;
 assign n_n550 = ( n_n262  &  n_n263 ) ;
 assign n_n1088 = ( n_n1583  &  n_n1118 ) ;
 assign n_n524 = ( n_n1121  &  n_n1074 ) ;
 assign n_n986 = ( n_n996  &  n_n1673 ) ;
 assign n_n968 = ( n_n997  &  n_n997 ) ;
 assign n_n779 = ( n_n1398  &  n_n789 ) ;
 assign n_n401 = ( n_n361  &  n_n360  &  n_n362 ) ;
 assign n_n398 = ( n_n766  &  n_n772 ) ;
 assign n_n392 = ( n_n749  &  n_n758 ) ;
 assign n_n381 = ( n_n726  &  n_n731 ) ;
 assign n_n745 = ( (~ n_n768) ) ;
 assign n_n364 = ( (~ n_n770) ) ;
 assign n_n361 = ( (~ n_n774) ) ;
 assign n_n353 = ( (~ n_n782) ) ;
 assign n_n786 = ( (~ n_n407) ) ;
 assign n_n797 = ( (~ n_n413) ) ;
 assign n_n850 = ( (~ n_n438) ) ;
 assign n_n333 = ( (~ n_n908) ) ;
 assign n_n864 = ( (~ n_n896) ) ;
 assign n_n328 = ( (~ n_n1379) ) ;
 assign n_n325 = ( (~ n_n1056) ) ;
 assign n_n899 = ( (~ n_n918) ) ;
 assign n_n939 = ( (~ n_n483) ) ;
 assign n_n949 = ( (~ n_n489) ) ;
 assign n_n982 = ( (~ n_n997) ) ;
 assign n_n998 = ( (~ n_n508) ) ;
 assign n_n1012 = ( (~ n_n1035) ) ;
 assign n_n281 = ( (~ n_n1105) ) ;
 assign n_n1066 = ( (~ n_n541) ) ;
 assign n_n1103 = ( (~ n_n552) ) ;
 assign n_n246 = ( (~ n_n1236) ) ;
 assign n_n223 = ( (~ n_n1157) ) ;
 assign n_n1145 = ( (~ n_n568) ) ;
 assign n_n185 = ( (~ n_n1278) ) ;
 assign n_n174 = ( (~ n_n1302) ) ;
 assign n_n151 = ( (~ n_n1246) ) ;
 assign n_n140 = ( (~ n_n1318) ) ;
 assign n_n96 = ( (~ n_n1337) ) ;
 assign n_n87 = ( (~ n_n1560) ) ;
 assign n_n1253 = ( (~ n_n582) ) ;
 assign n_n1310 = ( (~ n_n590) ) ;
 assign n_n1313 = ( (~ n_n593) ) ;
 assign n_n1408 = ( (~ n_n603) ) ;
 assign n_n37 = ( (~ n_n1573) ) ;
 assign n_n28 = ( (~ n_n1487) ) ;
 assign n_n1434 = ( (~ n_n615) ) ;
 assign n_n14 = ( (~ n_n1521) ) ;
 assign n_n1447 = ( (~ n_n1526) ) ;
 assign n_n1657 = ( (~ n_n1708) ) ;
 assign n_n676 = ( n_n3  &  n_n5 ) ;
 assign n_n1615 = ( n_n1714  &  n_n700 ) ;
 assign n_n639 = ( n_n1595  &  n_n1597 ) ;
 assign n_n1513 = ( n_n1550  &  n_n1691 ) ;
 assign n_n1504 = ( n_n1543  &  n_n1698 ) ;
 assign n_n627 = ( n_n1577  &  n_n1658 ) ;
 assign n_n618 = ( n_n12  &  n_n11  &  n_n13 ) ;
 assign n_n1413 = ( n_n1463  &  n_n701 ) ;
 assign n_n600 = ( n_n1467  &  n_n1559 ) ;
 assign n_n599 = ( n_n1442  &  n_n1526 ) ;
 assign n_n1368 = ( n_n1397  &  n_n702 ) ;
 assign n_n1351 = ( n_n1385  &  n_n1675 ) ;
 assign n_n1342 = ( n_n1382  &  n_n1678 ) ;
 assign n_n1333 = ( n_n1385  &  n_n1679 ) ;
 assign n_n1324 = ( n_n1383  &  n_n1681 ) ;
 assign n_n1298 = ( n_n1383  &  n_n1698 ) ;
 assign n_n1289 = ( n_n1385  &  n_n1700 ) ;
 assign n_n1280 = ( n_n1382  &  n_n1701 ) ;
 assign n_n1254 = ( n_n1383  &  n_n1707 ) ;
 assign n_n1245 = ( n_n1387  &  n_n1709 ) ;
 assign n_n578 = ( n_n85  &  n_n84  &  n_n86 ) ;
 assign n_n1227 = ( n_n1387  &  n_n1712 ) ;
 assign n_n1211 = ( n_n96  &  n_n95  &  n_n98  &  n_n97  &  n_n99  &  n_n92  &  n_n94  &  n_n93 ) ;
 assign n_n573 = ( n_n1306  &  n_n1307 ) ;
 assign n_n1149 = ( n_n1236  &  n_n1311  &  n_n1697 ) ;
 assign n_n1140 = ( n_n1652  &  n_n1182 ) ;
 assign n_n1131 = ( n_n1716  &  n_n1210 ) ;
 assign n_n563 = ( n_n225  &  n_n226 ) ;
 assign n_n549 = ( n_n264  &  n_n265 ) ;
 assign n_n1089 = ( n_n1583  &  n_n1117 ) ;
 assign n_n1038 = ( n_n1050  &  n_n536 ) ;
 assign n_n985 = ( n_n1088  &  n_n998 ) ;
 assign n_n969 = ( n_n998  &  n_n997 ) ;
 assign n_n406 = ( n_n347  &  n_n346  &  n_n348 ) ;
 assign n_n769 = ( n_n773  &  n_n773 ) ;
 assign n_n397 = ( n_n764  &  n_n859 ) ;
 assign n_n393 = ( n_n800  &  n_n768 ) ;
 assign n_n373 = ( n_n713  &  n_n708 ) ;
 assign n_n746 = ( (~ n_n394) ) ;
 assign n_n365 = ( (~ n_n783) ) ;
 assign n_n360 = ( (~ n_n912) ) ;
 assign n_n773 = ( (~ n_n403) ) ;
 assign n_n787 = ( (~ n_n408) ) ;
 assign n_n796 = ( (~ n_n412) ) ;
 assign n_n851 = ( (~ n_n439) ) ;
 assign n_n334 = ( (~ n_n876) ) ;
 assign n_n865 = ( (~ n_n450) ) ;
 assign n_n329 = ( (~ n_n890) ) ;
 assign n_n324 = ( (~ n_n915) ) ;
 assign n_n898 = ( (~ n_n467) ) ;
 assign n_n940 = ( (~ n_n964) ) ;
 assign n_n948 = ( (~ n_n488) ) ;
 assign n_n973 = ( (~ n_n495) ) ;
 assign n_n999 = ( (~ n_n509) ) ;
 assign n_n1010 = ( (~ n_n518) ) ;
 assign n_n1050 = ( (~ n_n538) ) ;
 assign n_n1065 = ( (~ n_n1178) ) ;
 assign n_n254 = ( (~ n_n1161) ) ;
 assign n_n247 = ( (~ n_n1168) ) ;
 assign n_n1119 = ( (~ n_n567) ) ;
 assign n_n1120 = ( (~ n_n1189) ) ;
 assign n_n184 = ( (~ n_n1279) ) ;
 assign n_n175 = ( (~ n_n1218) ) ;
 assign n_n150 = ( (~ n_n1252) ) ;
 assign n_n141 = ( (~ n_n1266) ) ;
 assign n_n95 = ( (~ n_n1342) ) ;
 assign n_n88 = ( (~ n_n1373) ) ;
 assign n_n1306 = ( (~ n_n586) ) ;
 assign n_n67 = ( (~ n_n1437) ) ;
 assign n_n60 = ( (~ n_n1356) ) ;
 assign n_n1410 = ( (~ n_n604) ) ;
 assign n_n1420 = ( (~ n_n607) ) ;
 assign n_n27 = ( (~ n_n1585) ) ;
 assign n_n20 = ( (~ n_n1517) ) ;
 assign n_n1438 = ( (~ n_n617) ) ;
 assign n_n1443 = ( (~ n_n619) ) ;
 assign n_n692 = ( (~ n_n1710) ) ;
 assign n_n1600 = ( n_n1641  &  n_n1639  &  n_n1640  &  n_n1636 ) ;
 assign n_n1589 = ( n_n1613  &  n_n1689 ) ;
 assign n_n1521 = ( n_n1550  &  n_n1686 ) ;
 assign n_n1485 = ( n_n1543  &  n_n1709 ) ;
 assign n_n1474 = ( n_n7  &  n_n1655 ) ;
 assign n_n1457 = ( n_n1608  &  n_n1541 ) ;
 assign n_n1441 = ( n_n1686  &  n_n1553  &  n_n1453 ) ;
 assign n_n1412 = ( n_n1603  &  n_n1454  &  n_n1710 ) ;
 assign n_n1401 = ( n_n1458  &  n_n1556 ) ;
 assign n_n1374 = ( n_n1397  &  n_n692 ) ;
 assign n_n1361 = ( n_n1536  &  n_n1427 ) ;
 assign n_n1358 = ( n_n1432  &  n_n1535 ) ;
 assign n_n1347 = ( n_n1384  &  n_n1676 ) ;
 assign n_n1336 = ( n_n1382  &  n_n1679 ) ;
 assign n_n1325 = ( n_n1384  &  n_n1680 ) ;
 assign n_n591 = ( n_n64  &  n_n66  &  n_n67 ) ;
 assign n_n1297 = ( n_n1384  &  n_n1699 ) ;
 assign n_n1286 = ( n_n1382  &  n_n1700 ) ;
 assign n_n1275 = ( n_n1384  &  n_n1703 ) ;
 assign n_n1264 = ( n_n1382  &  n_n1706 ) ;
 assign n_n1250 = ( n_n1387  &  n_n1708 ) ;
 assign n_n1239 = ( n_n1388  &  n_n1710 ) ;
 assign n_n1228 = ( n_n1388  &  n_n1712 ) ;
 assign n_n1214 = ( n_n5  &  n_n1372 ) ;
 assign n_n574 = ( n_n1391  &  n_n1391 ) ;
 assign n_n1193 = ( n_n1269  &  n_n1582 ) ;
 assign n_n1182 = ( n_n189  &  n_n188  &  n_n154  &  n_n190  &  n_n191  &  n_n185  &  n_n187  &  n_n186 ) ;
 assign n_n1170 = ( n_n581  &  n_n1313  &  n_n1694 ) ;
 assign n_n1159 = ( n_n1269  &  n_n1203  &  n_n1696 ) ;
 assign n_n1101 = ( n_n258  &  n_n259 ) ;
 assign n_n542 = ( n_n1126  &  n_n1195 ) ;
 assign n_n538 = ( n_n282  &  n_n281  &  n_n283 ) ;
 assign n_n500 = ( n_n1002  &  n_n1017 ) ;
 assign n_n493 = ( n_n999  &  n_n984 ) ;
 assign n_n405 = ( n_n350  &  n_n349  &  n_n351 ) ;
 assign n_n765 = ( n_n777  &  n_n777 ) ;
 assign n_n750 = ( n_n399  &  n_n401  &  n_n403  &  n_n427 ) ;
 assign n_n388 = ( n_n741  &  n_n771 ) ;
 assign n_n711 = ( (~ n_n715) ) ;
 assign n_n747 = ( (~ n_n761) ) ;
 assign n_n761 = ( (~ n_n399) ) ;
 assign n_n772 = ( (~ n_n402) ) ;
 assign n_n777 = ( (~ n_n405) ) ;
 assign n_n809 = ( (~ n_n420) ) ;
 assign n_n822 = ( (~ n_n847) ) ;
 assign n_n852 = ( (~ n_n440) ) ;
 assign n_n332 = ( (~ n_n889) ) ;
 assign n_n870 = ( (~ n_n452) ) ;
 assign n_n882 = ( (~ n_n459) ) ;
 assign n_n919 = ( (~ n_n941) ) ;
 assign n_n927 = ( (~ n_n974) ) ;
 assign n_n311 = ( (~ n_n961) ) ;
 assign n_n299 = ( (~ n_n1085) ) ;
 assign n_n954 = ( (~ n_n490) ) ;
 assign n_n977 = ( (~ n_n497) ) ;
 assign n_n990 = ( (~ n_n1039) ) ;
 assign n_n1022 = ( (~ n_n1078) ) ;
 assign n_n292 = ( (~ n_n1425) ) ;
 assign n_n290 = ( (~ n_n1063) ) ;
 assign n_n282 = ( (~ n_n1081) ) ;
 assign n_n280 = ( (~ n_n1080) ) ;
 assign n_n1075 = ( (~ n_n1116) ) ;
 assign n_n1095 = ( (~ n_n546) ) ;
 assign n_n262 = ( (~ n_n1141) ) ;
 assign n_n240 = ( (~ n_n1247) ) ;
 assign n_n232 = ( (~ n_n1172) ) ;
 assign n_n1115 = ( (~ n_n563) ) ;
 assign n_n217 = ( (~ n_n1160) ) ;
 assign n_n1121 = ( (~ n_n1190) ) ;
 assign n_n1176 = ( (~ n_n569) ) ;
 assign n_n206 = ( (~ n_n1298) ) ;
 assign n_n195 = ( (~ n_n1286) ) ;
 assign n_n165 = ( (~ n_n1297) ) ;
 assign n_n1668 = ( (~ n_n574) ) ;
 assign n_n153 = ( (~ n_n1232) ) ;
 assign n_n142 = ( (~ n_n1258) ) ;
 assign n_n139 = ( (~ n_n1332) ) ;
 assign n_n128 = ( (~ n_n1256) ) ;
 assign n_n117 = ( (~ n_n1334) ) ;
 assign n_n106 = ( (~ n_n1261) ) ;
 assign n_n90 = ( (~ n_n1469) ) ;
 assign n_n81 = ( (~ n_n1412) ) ;
 assign n_n1268 = ( (~ n_n584) ) ;
 assign n_n69 = ( (~ n_n1435) ) ;
 assign n_n61 = ( (~ n_n1450) ) ;
 assign n_n1372 = ( (~ n_n1408) ) ;
 assign n_n1387 = ( (~ n_n1511) ) ;
 assign n_n1398 = ( (~ n_n1539) ) ;
 assign n_n1417 = ( (~ n_n606) ) ;
 assign n_n34 = ( (~ n_n1578) ) ;
 assign n_n1427 = ( (~ n_n611) ) ;
 assign n_n24 = ( (~ n_n1587) ) ;
 assign n_n16 = ( (~ n_n1528) ) ;
 assign n_n8 = ( (~ n_n1524) ) ;
 assign n_n1505 = ( (~ n_n629) ) ;
 assign n_n1525 = ( (~ n_n640) ) ;
 assign n_n695 = ( (~ n_n1684) ) ;
 assign n_n665 = ( n_n1642  &  n_n1684 ) ;
 assign n_n661 = ( n_n1635  &  n_n1688 ) ;
 assign n_n635 = ( n_n1545  &  n_n1627 ) ;
 assign n_n624 = ( n_n1570  &  n_n701 ) ;
 assign n_n622 = ( n_n1565  &  n_n1656 ) ;
 assign n_n1456 = ( n_n1541  &  n_n1606 ) ;
 assign n_n619 = ( n_n9  &  n_n8  &  n_n10 ) ;
 assign n_n605 = ( n_n42  &  n_n41  &  n_n43 ) ;
 assign n_n1402 = ( n_n1464  &  n_n702 ) ;
 assign n_n1373 = ( n_n1710  &  n_n1557  &  n_n1408 ) ;
 assign n_n1362 = ( n_n1536  &  n_n1420 ) ;
 assign n_n1357 = ( n_n1434  &  n_n1535 ) ;
 assign n_n1348 = ( n_n1385  &  n_n1676 ) ;
 assign n_n1335 = ( n_n1381  &  n_n1679 ) ;
 assign n_n1326 = ( n_n1385  &  n_n1680 ) ;
 assign n_n1301 = ( n_n1382  &  n_n1698 ) ;
 assign n_n1296 = ( n_n1385  &  n_n1699 ) ;
 assign n_n1287 = ( n_n1381  &  n_n1700 ) ;
 assign n_n1274 = ( n_n1385  &  n_n1703 ) ;
 assign n_n1265 = ( n_n1381  &  n_n1706 ) ;
 assign n_n583 = ( n_n76  &  n_n75  &  n_n77 ) ;
 assign n_n1238 = ( n_n1383  &  n_n1710 ) ;
 assign n_n576 = ( n_n1375  &  n_n1404 ) ;
 assign n_n1213 = ( n_n5  &  n_n1377 ) ;
 assign n_n1204 = ( n_n152  &  n_n151  &  n_n154  &  n_n153  &  n_n155  &  n_n148  &  n_n150  &  n_n149 ) ;
 assign n_n1192 = ( n_n1236  &  n_n1582 ) ;
 assign n_n1183 = ( n_n182  &  n_n181  &  n_n146  &  n_n183  &  n_n184  &  n_n178  &  n_n180  &  n_n179 ) ;
 assign n_n1169 = ( n_n580  &  n_n1312  &  n_n1694 ) ;
 assign n_n1160 = ( n_n1203  &  n_n1696  &  n_n1201  &  n_n1202  &  n_n1200 ) ;
 assign n_n551 = ( n_n215  &  n_n260  &  n_n261 ) ;
 assign n_n543 = ( n_n1173  &  n_n1308 ) ;
 assign n_n1061 = ( n_n1394  &  n_n1103 ) ;
 assign n_n987 = ( n_n997  &  n_n1673 ) ;
 assign n_n494 = ( n_n994  &  n_n1000  &  n_n995 ) ;
 assign n_n404 = ( n_n352  &  n_n353 ) ;
 assign n_n767 = ( n_n778  &  n_n778 ) ;
 assign n_n396 = ( n_n757  &  n_n778 ) ;
 assign n_n389 = ( n_n745  &  n_n825 ) ;
 assign n_n717 = ( (~ n_n721) ) ;
 assign n_n748 = ( (~ n_n395) ) ;
 assign n_n363 = ( (~ n_n913) ) ;
 assign n_n356 = ( (~ n_n826) ) ;
 assign n_n349 = ( (~ n_n909) ) ;
 assign n_n810 = ( (~ n_n820) ) ;
 assign n_n821 = ( (~ n_n425) ) ;
 assign n_n853 = ( (~ n_n881) ) ;
 assign n_n859 = ( (~ n_n446) ) ;
 assign n_n871 = ( (~ n_n453) ) ;
 assign n_n881 = ( (~ n_n458) ) ;
 assign n_n920 = ( (~ n_n474) ) ;
 assign n_n926 = ( (~ n_n481) ) ;
 assign n_n301 = ( (~ n_n1374) ) ;
 assign n_n298 = ( (~ n_n972) ) ;
 assign n_n953 = ( (~ n_n987) ) ;
 assign n_n978 = ( (~ n_n992) ) ;
 assign n_n989 = ( (~ n_n1038) ) ;
 assign n_n1024 = ( (~ n_n522) ) ;
 assign n_n293 = ( (~ n_n1045) ) ;
 assign n_n289 = ( (~ n_n1414) ) ;
 assign n_n283 = ( (~ n_n1079) ) ;
 assign n_n279 = ( (~ n_n1082) ) ;
 assign n_n1070 = ( (~ n_n1113) ) ;
 assign n_n269 = ( (~ n_n1136) ) ;
 assign n_n263 = ( (~ n_n1142) ) ;
 assign n_n1109 = ( (~ n_n557) ) ;
 assign n_n233 = ( (~ n_n1166) ) ;
 assign n_n224 = ( (~ n_n1151) ) ;
 assign n_n218 = ( (~ n_n1188) ) ;
 assign n_n1122 = ( (~ n_n1191) ) ;
 assign n_n1173 = ( (~ n_n1195) ) ;
 assign n_n205 = ( (~ n_n1291) ) ;
 assign n_n196 = ( (~ n_n1292) ) ;
 assign n_n164 = ( (~ n_n1234) ) ;
 assign n_n1195 = ( (~ n_n573) ) ;
 assign n_n152 = ( (~ n_n1240) ) ;
 assign n_n143 = ( (~ n_n1251) ) ;
 assign n_n138 = ( (~ n_n1238) ) ;
 assign n_n129 = ( (~ n_n1249) ) ;
 assign n_n116 = ( (~ n_n1339) ) ;
 assign n_n107 = ( (~ n_n1350) ) ;
 assign n_n1236 = ( (~ n_n578) ) ;
 assign n_n1242 = ( (~ n_n580) ) ;
 assign n_n1260 = ( (~ n_n583) ) ;
 assign n_n68 = ( (~ n_n1359) ) ;
 assign n_n62 = ( (~ n_n1441) ) ;
 assign n_n58 = ( (~ n_n1355) ) ;
 assign n_n1388 = ( (~ n_n1512) ) ;
 assign n_n1394 = ( (~ n_n1532) ) ;
 assign n_n40 = ( (~ n_n1572) ) ;
 assign n_n1426 = ( (~ n_n610) ) ;
 assign n_n1429 = ( (~ n_n1583) ) ;
 assign n_n25 = ( (~ n_n1493) ) ;
 assign n_n15 = ( (~ n_n1594) ) ;
 assign n_n9 = ( (~ n_n1598) ) ;
 assign n_n1506 = ( (~ n_n630) ) ;
 assign n_n1522 = ( (~ n_n639) ) ;
 assign n_n696 = ( (~ n_n1685) ) ;
 assign n_n1579 = ( n_n1650  &  n_n1694 ) ;
 assign n_n1562 = ( n_n5  &  n_n1656 ) ;
 assign n_n1501 = ( n_n699  &  n_n1706 ) ;
 assign n_n1483 = ( n_n7  &  n_n692 ) ;
 assign n_n1472 = ( n_n1544  &  n_n1712 ) ;
 assign n_n1464 = ( n_n1548  &  n_n1551 ) ;
 assign n_n1444 = ( n_n1685  &  n_n1554  &  n_n1453 ) ;
 assign n_n604 = ( n_n1475  &  n_n1479 ) ;
 assign n_n1399 = ( n_n1542  &  n_n1532 ) ;
 assign n_n1379 = ( n_n1395  &  n_n1575 ) ;
 assign n_n1363 = ( n_n1536  &  n_n1421 ) ;
 assign n_n1356 = ( n_n1436  &  n_n1535 ) ;
 assign n_n1345 = ( n_n1386  &  n_n1677 ) ;
 assign n_n1338 = ( n_n1384  &  n_n1678 ) ;
 assign n_n1327 = ( n_n1386  &  n_n1680 ) ;
 assign n_n593 = ( n_n61  &  n_n60  &  n_n62 ) ;
 assign n_n1302 = ( n_n1381  &  n_n1698 ) ;
 assign n_n1295 = ( n_n1386  &  n_n1699 ) ;
 assign n_n1284 = ( n_n1384  &  n_n1701 ) ;
 assign n_n1277 = ( n_n1386  &  n_n1702 ) ;
 assign n_n1266 = ( n_n1386  &  n_n1706 ) ;
 assign n_n1259 = ( n_n1386  &  n_n1707 ) ;
 assign n_n1248 = ( n_n1383  &  n_n1708 ) ;
 assign n_n577 = ( n_n87  &  n_n88 ) ;
 assign n_n1216 = ( n_n1386  &  n_n1713 ) ;
 assign n_n1205 = ( n_n144  &  n_n143  &  n_n146  &  n_n145  &  n_n147  &  n_n140  &  n_n142  &  n_n141 ) ;
 assign n_n1191 = ( n_n1242  &  n_n1582 ) ;
 assign n_n1180 = ( n_n204  &  n_n203  &  n_n206  &  n_n205  &  n_n207  &  n_n200  &  n_n202  &  n_n201 ) ;
 assign n_n1172 = ( n_n585  &  n_n1316  &  n_n1694 ) ;
 assign n_n1161 = ( n_n575  &  n_n1196  &  n_n1695 ) ;
 assign n_n552 = ( n_n256  &  n_n255  &  n_n257 ) ;
 assign n_n1092 = ( n_n1399  &  n_n1145 ) ;
 assign n_n1073 = ( n_n1108  &  n_n563 ) ;
 assign n_n775 = ( n_n786  &  n_n786 ) ;
 assign n_n762 = ( n_n402  &  n_n405  &  n_n406  &  n_n446 ) ;
 assign n_n752 = ( n_n761  &  n_n761 ) ;
 assign n_n390 = ( n_n747  &  n_n773 ) ;
 assign n_n730 = ( (~ n_n743) ) ;
 assign n_n749 = ( (~ n_n396) ) ;
 assign n_n764 = ( (~ n_n777) ) ;
 assign n_n358 = ( (~ n_n779) ) ;
 assign n_n350 = ( (~ n_n784) ) ;
 assign n_n829 = ( (~ n_n429) ) ;
 assign n_n846 = ( (~ n_n436) ) ;
 assign n_n854 = ( (~ n_n441) ) ;
 assign n_n861 = ( (~ n_n447) ) ;
 assign n_n868 = ( (~ n_n904) ) ;
 assign n_n880 = ( (~ n_n917) ) ;
 assign n_n921 = ( (~ n_n475) ) ;
 assign n_n313 = ( (~ n_n1011) ) ;
 assign n_n302 = ( (~ n_n956) ) ;
 assign n_n941 = ( (~ n_n484) ) ;
 assign n_n964 = ( (~ n_n491) ) ;
 assign n_n974 = ( (~ n_n496) ) ;
 assign n_n988 = ( (~ n_n500) ) ;
 assign n_n1025 = ( (~ n_n523) ) ;
 assign n_n1034 = ( (~ n_n529) ) ;
 assign n_n1667 = ( (~ n_n533) ) ;
 assign n_n1049 = ( (~ n_n537) ) ;
 assign n_n278 = ( (~ n_n1110) ) ;
 assign n_n1091 = ( (~ n_n543) ) ;
 assign n_n271 = ( (~ n_n1134) ) ;
 assign n_n1098 = ( (~ n_n549) ) ;
 assign n_n1104 = ( (~ n_n553) ) ;
 assign n_n239 = ( (~ n_n1127) ) ;
 assign n_n1112 = ( (~ n_n560) ) ;
 assign n_n226 = ( (~ n_n1150) ) ;
 assign n_n1118 = ( (~ n_n566) ) ;
 assign n_n1123 = ( (~ n_n1192) ) ;
 assign n_n212 = ( (~ n_n1496) ) ;
 assign n_n1179 = ( (~ n_n572) ) ;
 assign n_n197 = ( (~ n_n1299) ) ;
 assign n_n181 = ( (~ n_n1301) ) ;
 assign n_n170 = ( (~ n_n1235) ) ;
 assign n_n163 = ( (~ n_n1225) ) ;
 assign n_n1197 = ( (~ n_n1310) ) ;
 assign n_n155 = ( (~ n_n1317) ) ;
 assign n_n144 = ( (~ n_n1245) ) ;
 assign n_n137 = ( (~ n_n1244) ) ;
 assign n_n126 = ( (~ n_n1320) ) ;
 assign n_n119 = ( (~ n_n1321) ) ;
 assign n_n108 = ( (~ n_n1344) ) ;
 assign n_n92 = ( (~ n_n1351) ) ;
 assign n_n84 = ( (~ n_n1409) ) ;
 assign n_n80 = ( (~ n_n1363) ) ;
 assign n_n73 = ( (~ n_n1502) ) ;
 assign n_n70 = ( (~ n_n1360) ) ;
 assign n_n1312 = ( (~ n_n592) ) ;
 assign n_n1314 = ( (~ n_n594) ) ;
 assign n_n1376 = ( (~ n_n1417) ) ;
 assign n_n1393 = ( (~ n_n599) ) ;
 assign n_n41 = ( (~ n_n1471) ) ;
 assign n_n1422 = ( (~ n_n609) ) ;
 assign n_n31 = ( (~ n_n1482) ) ;
 assign n_n1432 = ( (~ n_n614) ) ;
 assign n_n17 = ( (~ n_n1519) ) ;
 assign n_n10 = ( (~ n_n1530) ) ;
 assign n_n1455 = ( (~ n_n1537) ) ;
 assign n_n1475 = ( (~ n_n622) ) ;
 assign n_n1660 = ( (~ n_n1693) ) ;
 assign n_n1578 = ( n_n5  &  n_n1706 ) ;
 assign n_n1563 = ( n_n5  &  n_n1620 ) ;
 assign n_n1491 = ( n_n1544  &  n_n1708 ) ;
 assign n_n1482 = ( n_n699  &  n_n1710 ) ;
 assign n_n621 = ( n_n1656  &  n_n1712 ) ;
 assign n_n1463 = ( n_n1549  &  n_n1547 ) ;
 assign n_n1445 = ( n_n1684  &  n_n1554  &  n_n1453 ) ;
 assign n_n1409 = ( n_n1603  &  n_n1454  &  n_n1711 ) ;
 assign n_n1400 = ( n_n691  &  n_n1470 ) ;
 assign n_n1378 = ( n_n1422  &  n_n1706 ) ;
 assign n_n1364 = ( n_n1536  &  n_n1411 ) ;
 assign n_n1355 = ( n_n1438  &  n_n1535 ) ;
 assign n_n1346 = ( n_n1381  &  n_n1677 ) ;
 assign n_n1337 = ( n_n1387  &  n_n1679 ) ;
 assign n_n1328 = ( n_n1381  &  n_n1680 ) ;
 assign n_n592 = ( n_n64  &  n_n63  &  n_n65 ) ;
 assign n_n1303 = ( n_n1386  &  n_n1698 ) ;
 assign n_n1294 = ( n_n1381  &  n_n1699 ) ;
 assign n_n1285 = ( n_n1387  &  n_n1700 ) ;
 assign n_n1276 = ( n_n1381  &  n_n1702 ) ;
 assign n_n1267 = ( n_n1385  &  n_n1706 ) ;
 assign n_n1258 = ( n_n1381  &  n_n1707 ) ;
 assign n_n1249 = ( n_n1388  &  n_n1708 ) ;
 assign n_n1240 = ( n_n1387  &  n_n1710 ) ;
 assign n_n1215 = ( n_n1385  &  n_n1713 ) ;
 assign n_n1206 = ( n_n136  &  n_n135  &  n_n138  &  n_n137  &  n_n139  &  n_n132  &  n_n134  &  n_n133 ) ;
 assign n_n1190 = ( n_n1247  &  n_n1582 ) ;
 assign n_n1181 = ( n_n196  &  n_n195  &  n_n198  &  n_n197  &  n_n199  &  n_n192  &  n_n194  &  n_n193 ) ;
 assign n_n1171 = ( n_n583  &  n_n1315  &  n_n1694 ) ;
 assign n_n1162 = ( n_n578  &  n_n1198  &  n_n1695 ) ;
 assign n_n1102 = ( n_n1555  &  n_n1173 ) ;
 assign n_n544 = ( n_n274  &  n_n275 ) ;
 assign n_n1084 = ( n_n1429  &  n_n1119 ) ;
 assign n_n774 = ( n_n1398  &  n_n781 ) ;
 assign n_n400 = ( n_n834  &  n_n777 ) ;
 assign n_n751 = ( n_n768  &  n_n768 ) ;
 assign n_n739 = ( n_n704  &  n_n366 ) ;
 assign n_n740 = ( (~ n_n391) ) ;
 assign n_n754 = ( (~ n_n771) ) ;
 assign n_n763 = ( (~ n_n400) ) ;
 assign n_n357 = ( (~ n_n910) ) ;
 assign n_n351 = ( (~ n_n836) ) ;
 assign n_n830 = ( (~ n_n843) ) ;
 assign n_n845 = ( (~ n_n435) ) ;
 assign n_n855 = ( (~ n_n442) ) ;
 assign n_n331 = ( (~ n_n893) ) ;
 assign n_n869 = ( (~ n_n451) ) ;
 assign n_n879 = ( (~ n_n457) ) ;
 assign n_n929 = ( (~ n_n950) ) ;
 assign n_n312 = ( (~ n_n1057) ) ;
 assign n_n303 = ( (~ n_n1058) ) ;
 assign n_n942 = ( (~ n_n485) ) ;
 assign n_n1665 = ( (~ n_n976) ) ;
 assign n_n975 = ( (~ n_n986) ) ;
 assign n_n499 = ( (~ n_n1001) ) ;
 assign n_n1026 = ( (~ n_n1041) ) ;
 assign n_n291 = ( (~ n_n1419) ) ;
 assign n_n1046 = ( (~ n_n534) ) ;
 assign n_n284 = ( (~ n_n1076) ) ;
 assign n_n1051 = ( (~ n_n539) ) ;
 assign n_n1090 = ( (~ n_n542) ) ;
 assign n_n270 = ( (~ n_n1133) ) ;
 assign n_n264 = ( (~ n_n1139) ) ;
 assign n_n245 = ( (~ n_n1163) ) ;
 assign n_n238 = ( (~ n_n1494) ) ;
 assign n_n231 = ( (~ n_n1269) ) ;
 assign n_n225 = ( (~ n_n1156) ) ;
 assign n_n219 = ( (~ n_n1159) ) ;
 assign n_n1124 = ( (~ n_n1193) ) ;
 assign n_n213 = ( (~ n_n1213) ) ;
 assign n_n207 = ( (~ n_n1270) ) ;
 assign n_n198 = ( (~ n_n1221) ) ;
 assign n_n180 = ( (~ n_n1294) ) ;
 assign n_n171 = ( (~ n_n1290) ) ;
 assign n_n162 = ( (~ n_n1216) ) ;
 assign n_n1196 = ( (~ n_n1309) ) ;
 assign n_n154 = ( (~ n_n1223) ) ;
 assign n_n145 = ( (~ n_n1239) ) ;
 assign n_n136 = ( (~ n_n1250) ) ;
 assign n_n127 = ( (~ n_n1264) ) ;
 assign n_n118 = ( (~ n_n1328) ) ;
 assign n_n109 = ( (~ n_n1340) ) ;
 assign n_n91 = ( (~ n_n1366) ) ;
 assign n_n85 = ( (~ n_n1478) ) ;
 assign n_n79 = ( (~ n_n1488) ) ;
 assign n_n74 = ( (~ n_n1361) ) ;
 assign n_n1309 = ( (~ n_n589) ) ;
 assign n_n63 = ( (~ n_n1357) ) ;
 assign n_n57 = ( (~ n_n1445) ) ;
 assign n_n1375 = ( (~ n_n1410) ) ;
 assign n_n1386 = ( (~ n_n1510) ) ;
 assign n_n1411 = ( (~ n_n605) ) ;
 assign n_n1421 = ( (~ n_n608) ) ;
 assign n_n30 = ( (~ n_n1584) ) ;
 assign n_n23 = ( (~ n_n1516) ) ;
 assign n_n1436 = ( (~ n_n616) ) ;
 assign n_n1442 = ( (~ n_n1522) ) ;
 assign n_n1458 = ( (~ n_n1541) ) ;
 assign n_n1473 = ( (~ n_n621) ) ;
 assign n_n1659 = ( (~ n_n1694) ) ;
 assign n_n690 = ( n_n691  &  n_n697 ) ;
 assign n_n682 = ( n_n1708  &  n_n1685 ) ;
 assign n_n673 = ( n_n1710  &  n_n1711 ) ;
 assign n_n668 = ( n_n700  &  n_n699 ) ;
 assign n_n662 = ( n_n1633  &  n_n1687 ) ;
 assign n_n658 = ( n_n1693  &  n_n1609 ) ;
 assign n_n654 = ( n_n1655  &  n_n1711 ) ;
 assign n_n1500 = ( n_n1544  &  n_n1706 ) ;
 assign n_n625 = ( n_n1568  &  n_n1657 ) ;
 assign n_n1478 = ( n_n7  &  n_n1656 ) ;
 assign n_n620 = ( n_n1558  &  n_n1713 ) ;
 assign n_n1446 = ( n_n1457  &  n_n1525 ) ;
 assign n_n1340 = ( n_n1386  &  n_n1678 ) ;
 assign n_n1329 = ( n_n1382  &  n_n1680 ) ;
 assign n_n1544 = ( (~ n_n1610) ) ;
 assign n_n1559 = ( (~ n_n653) ) ;
 assign n_n1577 = ( (~ n_n693) ) ;
 assign n_n5 = ( (~ n_n698) ) ;
 assign n_n1613 = ( (~ n_n1653) ) ;
 assign n_n694 = ( n_n695  &  n_n696 ) ;
 assign n_n1638 = ( n_n1661  &  n_n1686 ) ;
 assign n_n674 = ( n_n1658  &  n_n1657 ) ;
 assign n_n667 = ( n_n700  &  n_n5 ) ;
 assign n_n1594 = ( n_n1613  &  n_n1687 ) ;
 assign n_n1580 = ( n_n1650  &  n_n1659 ) ;
 assign n_n655 = ( n_n1619  &  n_n692 ) ;
 assign n_n634 = ( n_n1580  &  n_n1627 ) ;
 assign n_n1488 = ( n_n7  &  n_n701 ) ;
 assign n_n623 = ( n_n1561  &  n_n692 ) ;
 assign n_n1466 = ( n_n691  &  n_n1556 ) ;
 assign n_n1448 = ( n_n1683  &  n_n1554  &  n_n1453 ) ;
 assign n_n1339 = ( n_n1385  &  n_n1678 ) ;
 assign n_n1330 = ( n_n1387  &  n_n1680 ) ;
 assign n_n1542 = ( (~ n_n648) ) ;
 assign n_n1561 = ( (~ n_n1656) ) ;
 assign n_n1576 = ( (~ n_n1575) ) ;
 assign n_n1603 = ( (~ n_n667) ) ;
 assign n_n1612 = ( (~ n_n1651) ) ;
 assign n_n1651 = ( n_n1715  &  n_n1716 ) ;
 assign n_n684 = ( n_n1706  &  n_n1683 ) ;
 assign n_n1623 = ( n_n1657  &  n_n1658  &  n_n701 ) ;
 assign n_n1602 = ( n_n1646  &  n_n1645 ) ;
 assign n_n1591 = ( n_n1613  &  n_n1688 ) ;
 assign n_n1584 = ( n_n1613  &  n_n1692 ) ;
 assign n_n1567 = ( n_n5  &  n_n1710 ) ;
 assign n_n1520 = ( n_n1540  &  n_n1638 ) ;
 assign n_n1487 = ( n_n699  &  n_n1709 ) ;
 assign n_n1476 = ( n_n1543  &  n_n1711 ) ;
 assign n_n1469 = ( n_n7  &  n_n702 ) ;
 assign n_n1449 = ( n_n1682  &  n_n1614  &  n_n1453 ) ;
 assign n_n1360 = ( n_n1430  &  n_n1535 ) ;
 assign n_n1349 = ( n_n1386  &  n_n1676 ) ;
 assign n_n1541 = ( (~ n_n647) ) ;
 assign n_n1564 = ( (~ n_n654) ) ;
 assign n_n1583 = ( (~ n_n1582) ) ;
 assign n_n1599 = ( (~ n_n665) ) ;
 assign n_n1611 = ( (~ n_n1650) ) ;
 assign n_n689 = ( n_n1652  &  n_n0 ) ;
 assign n_n683 = ( n_n1707  &  n_n1684 ) ;
 assign n_n675 = ( n_n4  &  n_n5 ) ;
 assign n_n666 = ( n_n695  &  n_n1683 ) ;
 assign n_n1592 = ( n_n1634  &  n_n1630  &  n_n1632  &  n_n1628 ) ;
 assign n_n1582 = ( n_n1693  &  n_n1672  &  n_n1609 ) ;
 assign n_n656 = ( n_n1622  &  n_n1709 ) ;
 assign n_n1530 = ( n_n699  &  n_n1679 ) ;
 assign n_n1486 = ( n_n1544  &  n_n1709 ) ;
 assign n_n1477 = ( n_n1544  &  n_n1711 ) ;
 assign n_n1468 = ( n_n1543  &  n_n1713 ) ;
 assign n_n1450 = ( n_n1682  &  n_n1615  &  n_n1453 ) ;
 assign n_n1359 = ( n_n1431  &  n_n1535 ) ;
 assign n_n1350 = ( n_n1384  &  n_n1675 ) ;
 assign n_n1540 = ( (~ n_n1608) ) ;
 assign n_n1565 = ( (~ n_n692) ) ;
 assign n_n1581 = ( (~ n_n658) ) ;
 assign n_n1601 = ( (~ n_n666) ) ;
 assign n_n1610 = ( (~ n_n670) ) ;
 assign n_n1661 = ( (~ n_n694) ) ;
 assign n_n688 = ( n_n1694  &  n_n1717 ) ;
 assign n_n679 = ( n_n1711  &  n_n1688 ) ;
 assign n_n1616 = ( n_n1714  &  n_n697  &  n_n700 ) ;
 assign n_n670 = ( n_n698  &  n_n699 ) ;
 assign n_n664 = ( n_n1637  &  n_n1685 ) ;
 assign n_n659 = ( n_n1631  &  n_n1690 ) ;
 assign n_n1572 = ( n_n5  &  n_n1658 ) ;
 assign n_n1529 = ( n_n699  &  n_n1680 ) ;
 assign n_n638 = ( n_n1590  &  n_n1593 ) ;
 assign n_n631 = ( n_n1545  &  n_n676 ) ;
 assign n_n1496 = ( n_n1544  &  n_n1707 ) ;
 assign n_n1451 = ( n_n1682  &  n_n1616  &  n_n1453 ) ;
 assign n_n1397 = ( n_n1537  &  n_n1532 ) ;
 assign n_n1369 = ( n_n1397  &  n_n1655 ) ;
 assign n_n495 = ( n_n1044  &  n_n998 ) ;
 assign n_n962 = ( n_n1017  &  n_n996 ) ;
 assign n_n399 = ( n_n364  &  n_n363  &  n_n365 ) ;
 assign n_n394 = ( n_n760  &  n_n761 ) ;
 assign n_n354 = ( (~ n_n875) ) ;
 assign n_n1539 = ( (~ n_n646) ) ;
 assign n_n4 = ( (~ n_n1697) ) ;
 assign n_n1634 = ( (~ n_n680) ) ;
 assign n_n1644 = ( (~ n_n685) ) ;
 assign n_n1655 = ( (~ n_n1712) ) ;
 assign n_n1650 = ( n_n1696  &  n_n1717 ) ;
 assign n_n678 = ( n_n1712  &  n_n1689 ) ;
 assign n_n671 = ( n_n698  &  n_n1714  &  n_n1718 ) ;
 assign n_n1609 = ( n_n1718  &  n_n698  &  n_n700 ) ;
 assign n_n1598 = ( n_n1613  &  n_n1685 ) ;
 assign n_n1585 = ( n_n1613  &  n_n1691 ) ;
 assign n_n1573 = ( n_n5  &  n_n1624 ) ;
 assign n_n1528 = ( n_n699  &  n_n1681 ) ;
 assign n_n1519 = ( n_n1550  &  n_n1687 ) ;
 assign n_n630 = ( n_n1580  &  n_n676 ) ;
 assign n_n1497 = ( n_n699  &  n_n1707 ) ;
 assign n_n1470 = ( n_n1712  &  n_n1621  &  n_n702  &  n_n1575 ) ;
 assign n_n1396 = ( n_n1539  &  n_n1533 ) ;
 assign n_n1371 = ( n_n1397  &  n_n1656 ) ;
 assign n_n972 = ( n_n994  &  n_n1000 ) ;
 assign n_n963 = ( n_n1017  &  n_n1000 ) ;
 assign n_n759 = ( n_n772  &  n_n772 ) ;
 assign n_n395 = ( n_n756  &  n_n763 ) ;
 assign n_n362 = ( (~ n_n812) ) ;
 assign n_n1538 = ( (~ n_n1606) ) ;
 assign n_n1625 = ( (~ n_n675) ) ;
 assign n_n1633 = ( (~ n_n1688) ) ;
 assign n_n1645 = ( (~ n_n686) ) ;
 assign n_n691 = ( (~ n_n1714) ) ;
 assign n_n687 = ( n_n1717  &  n_n1716  &  n_n1719 ) ;
 assign n_n681 = ( n_n1709  &  n_n1686 ) ;
 assign n_n672 = ( n_n1656  &  n_n1655 ) ;
 assign n_n1607 = ( n_n1648  &  n_n1717  &  n_n1719 ) ;
 assign n_n663 = ( n_n696  &  n_n1686 ) ;
 assign n_n660 = ( n_n1629  &  n_n1689 ) ;
 assign n_n657 = ( n_n1657  &  n_n1707 ) ;
 assign n_n1527 = ( n_n1544  &  n_n1681 ) ;
 assign n_n1516 = ( n_n1550  &  n_n1689 ) ;
 assign n_n633 = ( n_n1579  &  n_n1627 ) ;
 assign n_n1498 = ( n_n7  &  n_n1658 ) ;
 assign n_n1480 = ( n_n1544  &  n_n1710 ) ;
 assign n_n1418 = ( n_n1604  &  n_n1454  &  n_n1708 ) ;
 assign n_n602 = ( n_n45  &  n_n44  &  n_n46 ) ;
 assign n_n546 = ( n_n270  &  n_n271 ) ;
 assign n_n976 = ( n_n499  &  n_n988 ) ;
 assign n_n491 = ( n_n991  &  n_n977 ) ;
 assign n_n784 = ( n_n1398  &  n_n794 ) ;
 assign n_n402 = ( n_n358  &  n_n357  &  n_n359 ) ;
 assign n_n757 = ( (~ n_n772) ) ;
 assign n_n1626 = ( (~ n_n1696) ) ;
 assign n_n1636 = ( (~ n_n681) ) ;
 assign n_n2 = ( (~ n_n1660) ) ;
 assign n_n1654 = ( (~ n_n690) ) ;
 assign n_n1647 = ( n_n1717  &  n_n1718 ) ;
 assign n_n680 = ( n_n1710  &  n_n1687 ) ;
 assign n_n1619 = ( n_n1655  &  n_n1656  &  n_n702 ) ;
 assign n_n669 = ( n_n1648  &  n_n1719 ) ;
 assign n_n1596 = ( n_n1613  &  n_n1686 ) ;
 assign n_n1587 = ( n_n1613  &  n_n1690 ) ;
 assign n_n1575 = ( n_n1623  &  n_n693 ) ;
 assign n_n641 = ( n_n1599  &  n_n1601 ) ;
 assign n_n1517 = ( n_n1550  &  n_n1688 ) ;
 assign n_n632 = ( n_n1546  &  n_n676 ) ;
 assign n_n628 = ( n_n1571  &  n_n693 ) ;
 assign n_n1490 = ( n_n1543  &  n_n1708 ) ;
 assign n_n606 = ( n_n1484  &  n_n1489 ) ;
 assign n_n603 = ( n_n1473  &  n_n1564 ) ;
 assign n_n1085 = ( n_n1583  &  n_n1115 ) ;
 assign n_n496 = ( n_n296  &  n_n297 ) ;
 assign n_n965 = ( n_n994  &  n_n996 ) ;
 assign n_n783 = ( n_n1452  &  n_n796 ) ;
 assign n_n403 = ( n_n355  &  n_n354  &  n_n356 ) ;
 assign n_n741 = ( (~ n_n755) ) ;
 assign n_n3 = ( (~ n_n1695) ) ;
 assign n_n1635 = ( (~ n_n1687) ) ;
 assign n_n1 = ( (~ n_n1672) ) ;
 assign n_n697 = ( (~ n_n1715) ) ;
 assign n_n652 = ( n_n697  &  n_n1652 ) ;
 assign n_n645 = ( n_n1652  &  n_n1648 ) ;
 assign n_n1439 = ( n_n1687  &  n_n1552  &  n_n1453 ) ;
 assign n_n611 = ( n_n33  &  n_n32  &  n_n34 ) ;
 assign n_n1074 = ( n_n1109  &  n_n564 ) ;
 assign n_n955 = ( n_n996  &  n_n703  &  n_n1673 ) ;
 assign n_n484 = ( n_n298  &  n_n299 ) ;
 assign n_n481 = ( n_n947  &  n_n973 ) ;
 assign n_n913 = ( n_n1396  &  n_n936 ) ;
 assign n_n419 = ( n_n815  &  n_n904 ) ;
 assign n_n795 = ( n_n479  &  n_n339 ) ;
 assign n_n731 = ( (~ n_n385) ) ;
 assign n_n1586 = ( (~ n_n659) ) ;
 assign n_n1604 = ( (~ n_n668) ) ;
 assign n_n1620 = ( (~ n_n1619) ) ;
 assign n_n1630 = ( (~ n_n678) ) ;
 assign n_n1642 = ( (~ n_n1683) ) ;
 assign n_n1653 = ( (~ n_n689) ) ;
 assign n_n1550 = ( n_n1653  &  n_n1652 ) ;
 assign n_n646 = ( n_n697  &  n_n1648  &  n_n1717  &  n_n1719 ) ;
 assign n_n617 = ( n_n15  &  n_n14  &  n_n16 ) ;
 assign n_n1428 = ( n_n1604  &  n_n1454  &  n_n1706 ) ;
 assign n_n1062 = ( n_n1399  &  n_n1100 ) ;
 assign n_n490 = ( n_n1643  &  n_n968 ) ;
 assign n_n485 = ( n_n967  &  n_n971  &  n_n1052 ) ;
 assign n_n480 = ( n_n1000  &  n_n995  &  n_n994  &  n_n964 ) ;
 assign n_n914 = ( n_n1455  &  n_n940 ) ;
 assign n_n418 = ( n_n814  &  n_n817 ) ;
 assign n_n412 = ( n_n818  &  n_n808 ) ;
 assign n_n718 = ( (~ n_n380) ) ;
 assign n_n1588 = ( (~ n_n660) ) ;
 assign n_n699 = ( (~ n_n1652) ) ;
 assign n_n1621 = ( (~ n_n673) ) ;
 assign n_n1629 = ( (~ n_n1690) ) ;
 assign n_n1643 = ( (~ n_n1673) ) ;
 assign n_n0 = ( (~ n_n1671) ) ;
 assign n_n653 = ( n_n702  &  n_n1655 ) ;
 assign n_n647 = ( n_n1718  &  n_n1717  &  n_n1719 ) ;
 assign n_n539 = ( n_n279  &  n_n278  &  n_n280 ) ;
 assign n_n952 = ( n_n969  &  n_n1673 ) ;
 assign n_n938 = ( n_n302  &  n_n301  &  n_n303 ) ;
 assign n_n930 = ( n_n944  &  n_n1673 ) ;
 assign n_n915 = ( n_n1459  &  n_n945 ) ;
 assign n_n432 = ( n_n861  &  n_n850 ) ;
 assign n_n426 = ( n_n828  &  n_n847 ) ;
 assign n_n712 = ( (~ n_n716) ) ;
 assign n_n1552 = ( (~ n_n1614) ) ;
 assign n_n1568 = ( (~ n_n701) ) ;
 assign n_n1622 = ( (~ n_n674) ) ;
 assign n_n1632 = ( (~ n_n679) ) ;
 assign n_n1640 = ( (~ n_n683) ) ;
 assign n_n1652 = ( (~ n_n1716) ) ;
 assign n_n1556 = ( n_n1618  &  n_n1713 ) ;
 assign n_n648 = ( n_n698  &  n_n1652  &  n_n1648 ) ;
 assign n_n1039 = ( n_n1051  &  n_n537 ) ;
 assign n_n951 = ( n_n965  &  n_n1673 ) ;
 assign n_n483 = ( n_n300  &  n_n499 ) ;
 assign n_n928 = ( n_n974  &  n_n974 ) ;
 assign n_n917 = ( n_n994  &  n_n964  &  n_n995  &  n_n996 ) ;
 assign n_n838 = ( n_n1398  &  n_n856 ) ;
 assign n_n824 = ( n_n1452  &  n_n847 ) ;
 assign n_n372 = ( n_n709  &  n_n710 ) ;
 assign n_n1553 = ( (~ n_n1615) ) ;
 assign n_n1566 = ( (~ n_n655) ) ;
 assign n_n1624 = ( (~ n_n1623) ) ;
 assign n_n1631 = ( (~ n_n1689) ) ;
 assign n_n1641 = ( (~ n_n684) ) ;
 assign n_n1649 = ( (~ n_n688) ) ;
 assign n_n1543 = ( n_n1610  &  n_n698 ) ;
 assign n_n525 = ( n_n1122  &  n_n1073 ) ;
 assign n_n472 = ( n_n932  &  n_n954 ) ;
 assign n_n892 = ( n_n321  &  n_n320  &  n_n322 ) ;
 assign n_n456 = ( n_n916  &  n_n917 ) ;
 assign n_n449 = ( n_n978  &  n_n896 ) ;
 assign n_n448 = ( n_n880  &  n_n962 ) ;
 assign n_n438 = ( n_n864  &  n_n939 ) ;
 assign n_n720 = ( n_n723  &  n_n1531  &  n_n732 ) ;
 assign n_n1551 = ( (~ n_n652) ) ;
 assign n_n1554 = ( (~ n_n1616) ) ;
 assign n_n1570 = ( (~ n_n1657) ) ;
 assign n_n1595 = ( (~ n_n663) ) ;
 assign n_n698 = ( (~ n_n1717) ) ;
 assign n_n1637 = ( (~ n_n1686) ) ;
 assign n_n1648 = ( (~ n_n1718) ) ;
 assign n_n1560 = ( n_n702  &  n_n1711 ) ;
 assign n_n518 = ( n_n1020  &  n_n1194 ) ;
 assign n_n904 = ( n_n917  &  n_n1673 ) ;
 assign n_n893 = ( n_n939  &  n_n939 ) ;
 assign n_n455 = ( n_n329  &  n_n328  &  n_n330 ) ;
 assign n_n450 = ( n_n897  &  n_n879 ) ;
 assign n_n447 = ( n_n894  &  n_n896 ) ;
 assign n_n439 = ( n_n862  &  n_n878 ) ;
 assign n_n734 = ( n_n739  &  n_n1693 ) ;
 assign n_n1549 = ( (~ n_n651) ) ;
 assign n_n1555 = ( (~ n_n691) ) ;
 assign n_n1569 = ( (~ n_n656) ) ;
 assign n_n1597 = ( (~ n_n664) ) ;
 assign n_n1608 = ( (~ n_n1607) ) ;
 assign n_n1639 = ( (~ n_n682) ) ;
 assign n_n1646 = ( (~ n_n687) ) ;
 assign n_n510 = ( n_n1012  &  n_n1012 ) ;
 assign n_n471 = ( n_n945  &  n_n974 ) ;
 assign n_n890 = ( n_n700  &  n_n479 ) ;
 assign n_n458 = ( n_n920  &  n_n898 ) ;
 assign n_n451 = ( n_n929  &  n_n882 ) ;
 assign n_n1548 = ( (~ n_n650) ) ;
 assign n_n1557 = ( (~ n_n702) ) ;
 assign n_n1574 = ( (~ n_n657) ) ;
 assign n_n1590 = ( (~ n_n661) ) ;
 assign n_n1606 = ( (~ n_n669) ) ;
 assign n_n1617 = ( (~ n_n671) ) ;
 assign n_n1628 = ( (~ n_n677) ) ;
 assign n_n501 = ( n_n1040  &  n_n1038 ) ;
 assign n_n470 = ( n_n924  &  n_n946 ) ;
 assign n_n891 = ( n_n324  &  n_n323  &  n_n325 ) ;
 assign n_n457 = ( n_n899  &  n_n993 ) ;
 assign n_n452 = ( n_n883  &  n_n986 ) ;
 assign n_n1547 = ( (~ n_n649) ) ;
 assign n_n1558 = ( (~ n_n1655) ) ;
 assign n_n1571 = ( (~ n_n1658) ) ;
 assign n_n1593 = ( (~ n_n662) ) ;
 assign n_n1605 = ( (~ n_n1647) ) ;
 assign n_n1618 = ( (~ n_n672) ) ;
 assign n_n1627 = ( (~ n_n676) ) ;


endmodule

