module cps (
	i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, 
	i_8_, i_9_, i_10_, i_11_, i_12_, i_13_, i_14_, i_15_, i_16_, i_17_, 
	i_18_, i_19_, i_20_, i_21_, i_22_, i_23_, o_0_, o_1_, o_2_, o_3_, 
	o_4_, o_5_, o_6_, o_7_, o_8_, o_9_, o_10_, o_11_, o_12_, o_13_, 
	o_14_, o_15_, o_16_, o_17_, o_18_, o_19_, o_20_, o_21_, o_22_, o_23_, 
	o_24_, o_25_, o_26_, o_27_, o_28_, o_29_, o_30_, o_31_, o_32_, o_33_, 
	o_34_, o_35_, o_36_, o_37_, o_38_, o_39_, o_40_, o_41_, o_42_, o_43_, 
	o_44_, o_45_, o_46_, o_47_, o_48_, o_49_, o_50_, o_51_, o_52_, o_53_, 
	o_54_, o_55_, o_56_, o_57_, o_58_, o_59_, o_60_, o_61_, o_62_, o_63_, 
	o_64_, o_65_, o_66_, o_67_, o_68_, o_69_, o_70_, o_71_, o_72_, o_73_, 
	o_74_, o_75_, o_76_, o_77_, o_78_, o_79_, o_80_, o_81_, o_82_, o_83_, 
	o_84_, o_85_, o_86_, o_87_, o_88_, o_89_, o_90_, o_91_, o_92_, o_93_, 
	o_94_, o_95_, o_96_, o_97_, o_98_, o_99_, o_100_, o_101_, o_102_, o_103_, 
	o_104_, o_105_, o_106_, o_107_, o_108_);

input i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, i_8_, i_9_, i_10_, i_11_, i_12_, i_13_, i_14_, i_15_, i_16_, i_17_, i_18_, i_19_, i_20_, i_21_, i_22_, i_23_;

output o_0_, o_1_, o_2_, o_3_, o_4_, o_5_, o_6_, o_7_, o_8_, o_9_, o_10_, o_11_, o_12_, o_13_, o_14_, o_15_, o_16_, o_17_, o_18_, o_19_, o_20_, o_21_, o_22_, o_23_, o_24_, o_25_, o_26_, o_27_, o_28_, o_29_, o_30_, o_31_, o_32_, o_33_, o_34_, o_35_, o_36_, o_37_, o_38_, o_39_, o_40_, o_41_, o_42_, o_43_, o_44_, o_45_, o_46_, o_47_, o_48_, o_49_, o_50_, o_51_, o_52_, o_53_, o_54_, o_55_, o_56_, o_57_, o_58_, o_59_, o_60_, o_61_, o_62_, o_63_, o_64_, o_65_, o_66_, o_67_, o_68_, o_69_, o_70_, o_71_, o_72_, o_73_, o_74_, o_75_, o_76_, o_77_, o_78_, o_79_, o_80_, o_81_, o_82_, o_83_, o_84_, o_85_, o_86_, o_87_, o_88_, o_89_, o_90_, o_91_, o_92_, o_93_, o_94_, o_95_, o_96_, o_97_, o_98_, o_99_, o_100_, o_101_, o_102_, o_103_, o_104_, o_105_, o_106_, o_107_, o_108_;

wire n11, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n24, n25, n23, n26, n27, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n42, n44, n45, n46, n47, n43, n49, n50, n51, n52, n48, n54, n53, n55, n56, n58, n59, n60, n57, n62, n63, n65, n66, n67, n68, n64, n69, n71, n72, n73, n74, n70, n75, n77, n78, n76, n81, n82, n80, n83, n85, n87, n88, n86, n91, n94, n90, n95, n96, n97, n98, n99, n100, n101, n104, n105, n108, n102, n111, n113, n115, n116, n109, n117, n119, n122, n123, n124, n125, n118, n128, n130, n131, n132, n135, n134, n136, n137, n138, n140, n139, n141, n142, n144, n145, n147, n148, n152, n153, n154, n155, n156, n151, n157, n158, n159, n160, n161, n167, n168, n166, n171, n173, n177, n178, n179, n180, n182, n183, n184, n185, n186, n188, n189, n191, n192, n194, n195, n196, n197, n199, n201, n203, n204, n205, n206, n209, n207, n211, n210, n214, n219, n220, n221, n222, n225, n227, n228, n229, n230, n231, n232, n233, n234, n236, n237, n239, n240, n241, n243, n245, n246, n244, n249, n248, n247, n251, n252, n250, n254, n255, n256, n257, n258, n259, n253, n262, n261, n260, n263, n267, n268, n269, n270, n273, n275, n276, n277, n278, n280, n281, n279, n283, n282, n288, n286, n285, n289, n290, n291, n293, n295, n297, n299, n300, n305, n303, n306, n308, n309, n310, n311, n313, n314, n318, n319, n320, n322, n323, n326, n325, n324, n328, n327, n330, n331, n335, n337, n339, n340, n338, n343, n341, n345, n346, n347, n349, n350, n353, n351, n355, n354, n357, n356, n360, n359, n364, n367, n371, n372, n374, n375, n373, n377, n376, n380, n379, n378, n382, n384, n385, n386, n387, n381, n389, n390, n388, n392, n391, n396, n395, n393, n397, n399, n398, n401, n403, n400, n404, n407, n406, n414, n417, n418, n421, n423, n422, n425, n427, n428, n429, n430, n431, n426, n433, n434, n435, n438, n437, n436, n440, n439, n441, n443, n442, n444, n445, n447, n448, n449, n451, n453, n452, n457, n456, n459, n460, n463, n461, n465, n466, n468, n467, n471, n472, n470, n474, n475, n476, n478, n473, n480, n479, n484, n482, n486, n487, n485, n489, n488, n493, n490, n496, n494, n497, n498, n502, n506, n505, n508, n507, n510, n511, n509, n512, n514, n513, n518, n519, n523, n524, n522, n526, n527, n528, n529, n525, n530, n531, n532, n533, n534, n536, n537, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n553, n554, n555, n556, n557, n558, n559, n560, n561, n563, n564, n565, n566, n567, n568, n570, n571, n572, n573, n574, n575, n576, n577, n579, n580, n581, n583, n584, n585, n587, n588, n589, n590, n591, n593, n594, n595, n596, n597, n598, n600, n601, n604, n606, n605, n607, n609, n611, n612, n613, n615, n617, n620, n621, n622, n624, n623, n627, n626, n630, n631, n634, n637, n636, n635, n638, n639, n641, n643, n644, n645, n646, n647, n648, n650, n652, n651, n653, n655, n657, n658, n659, n661;

assign o_0_ = ( (~ n525) ) ;
 assign o_1_ = ( o_99_ ) | ( n157 ) | ( n158 ) | ( n159 ) | ( n160 ) | ( n161 ) | ( (~ n482) ) | ( (~ n648) ) ;
 assign o_2_ = ( (~ n151) ) ;
 assign o_3_ = ( i_9_  &  (~ n168)  &  n191 ) ;
 assign o_4_ = ( (~ n168)  &  n189 ) ;
 assign o_5_ = ( (~ n587) ) ;
 assign o_6_ = ( (~ i_12_)  &  n186  &  n188 ) ;
 assign o_7_ = ( n185  &  (~ n195)  &  n514 ) ;
 assign o_8_ = ( n173  &  n185  &  (~ n293) ) ;
 assign o_9_ = ( n185  &  n182 ) ;
 assign o_10_ = ( n180  &  n185  &  (~ n293) ) ;
 assign o_11_ = ( n184  &  n185 ) ;
 assign o_12_ = ( n514  &  n177 ) ;
 assign o_13_ = ( (~ n195)  &  (~ n197)  &  (~ n222) ) ;
 assign o_14_ = ( n514  &  n183 ) ;
 assign o_15_ = ( n183  &  n180 ) ;
 assign o_16_ = ( (~ n590) ) ;
 assign o_17_ = ( n179  &  (~ n508) ) ;
 assign o_18_ = ( n514  &  n179 ) ;
 assign o_19_ = ( (~ n195)  &  n514  &  (~ n549) ) ;
 assign o_20_ = ( n182  &  (~ n549) ) ;
 assign o_21_ = ( n179  &  n180 ) ;
 assign o_22_ = ( n184  &  (~ n549) ) ;
 assign o_23_ = ( (~ n509) ) ;
 assign o_24_ = ( (~ n46) ) | ( n144 ) | ( n145 ) | ( n147 ) | ( n148 ) | ( (~ n482) ) | ( (~ n645) ) ;
 assign o_25_ = ( (~ n595) ) ;
 assign o_26_ = ( (~ n594) ) ;
 assign o_27_ = ( i_5_  &  n142 ) | ( i_5_  &  (~ n635) ) ;
 assign o_28_ = ( (~ n141) ) ;
 assign o_29_ = ( (~ n139) ) ;
 assign o_30_ = ( (~ n11) ) ;
 assign o_31_ = ( (~ n138) ) ;
 assign o_32_ = ( (~ n604) ) ;
 assign o_33_ = ( (~ n137) ) ;
 assign o_34_ = ( o_14_ ) | ( (~ n433) ) ;
 assign o_35_ = ( (~ n136) ) ;
 assign o_36_ = ( (~ n134) ) ;
 assign o_37_ = ( (~ n426) ) ;
 assign o_38_ = ( n128 ) | ( n130 ) | ( n131 ) | ( n132 ) | ( (~ n398) ) | ( (~ n417) ) | ( (~ n621) ) | ( (~ n622) ) ;
 assign o_39_ = ( (~ n381) ) ;
 assign o_40_ = ( (~ n118) ) ;
 assign o_41_ = ( (~ n117) ) ;
 assign o_42_ = ( (~ n109) ) ;
 assign o_43_ = ( (~ n32) ) ;
 assign o_44_ = ( (~ n102) ) ;
 assign o_45_ = ( (~ n101) ) ;
 assign o_46_ = ( (~ n13) ) ;
 assign o_47_ = ( n97 ) | ( n98 ) | ( n99 ) | ( n100 ) ;
 assign o_48_ = ( n178  &  i_22_ ) ;
 assign o_49_ = ( i_20_  &  (~ i_22_)  &  n177 ) ;
 assign o_50_ = ( (~ n96) ) ;
 assign o_51_ = ( (~ n14) ) ;
 assign o_52_ = ( o_7_ ) | ( o_47_ ) ;
 assign o_53_ = ( n95 ) | ( (~ n96) ) ;
 assign o_54_ = ( (~ n90) ) ;
 assign o_55_ = ( (~ n86) ) ;
 assign o_56_ = ( n62 ) | ( n63 ) | ( n83 ) | ( n85 ) | ( (~ n88) ) ;
 assign o_57_ = ( (~ n80) ) ;
 assign o_58_ = ( (~ n540)  &  (~ n547) ) ;
 assign o_59_ = ( (~ n76) ) ;
 assign o_60_ = ( (~ n15) ) ;
 assign o_61_ = ( (~ n16) ) ;
 assign o_62_ = ( n173  &  (~ n293)  &  (~ n299) ) ;
 assign o_63_ = ( (~ n17) ) ;
 assign o_64_ = ( (~ n18) ) ;
 assign o_65_ = ( (~ n75) ) ;
 assign o_66_ = ( (~ n279) ) ;
 assign o_67_ = ( (~ n19) ) ;
 assign o_68_ = ( o_12_ ) | ( n20 ) ;
 assign o_69_ = ( (~ n21) ) ;
 assign o_70_ = ( (~ n70) ) ;
 assign o_71_ = ( i_21_  &  n171  &  (~ n268) ) ;
 assign o_72_ = ( (~ n69) ) ;
 assign o_73_ = ( (~ n253) ) ;
 assign o_74_ = ( (~ n64) ) ;
 assign o_75_ = ( n62 ) | ( n63 ) | ( (~ n73) ) | ( (~ n210) ) | ( (~ n276) ) ;
 assign o_76_ = ( n171  &  n227  &  (~ n300) ) ;
 assign o_77_ = ( (~ n57) ) ;
 assign o_78_ = ( o_76_ ) | ( (~ n42) ) | ( n55 ) | ( n56 ) ;
 assign o_79_ = ( (~ n53) ) ;
 assign o_80_ = ( o_17_ ) | ( (~ n53) ) ;
 assign o_81_ = ( (~ n48) ) ;
 assign o_82_ = ( (~ n43) ) ;
 assign o_83_ = ( (~ n42) ) ;
 assign o_84_ = ( o_13_ ) | ( n39 ) | ( (~ n210) ) | ( (~ n273) ) ;
 assign o_85_ = ( (~ i_9_)  &  n209  &  n541 ) ;
 assign o_86_ = ( n36 ) | ( n37 ) | ( n38 ) ;
 assign o_87_ = ( (~ n32) ) | ( n34 ) | ( n35 ) | ( (~ n587) ) ;
 assign o_88_ = ( (~ n33) ) ;
 assign o_89_ = ( (~ i_1_) ) | ( n30 ) | ( n31 ) | ( (~ n209) ) ;
 assign o_90_ = ( (~ n22) ) ;
 assign o_91_ = ( (~ n201)  &  (~ n540) ) ;
 assign o_92_ = ( n209  &  n188 ) ;
 assign o_93_ = ( (~ n23) ) ;
 assign o_95_ = ( (~ n276) ) ;
 assign o_96_ = ( i_12_  &  n311  &  n209 ) ;
 assign o_97_ = ( (~ n166) ) ;
 assign o_98_ = ( (~ n26) ) ;
 assign o_99_ = ( i_9_  &  (~ i_10_)  &  n186  &  n245 ) ;
 assign o_100_ = ( (~ n27) ) ;
 assign o_101_ = ( (~ n195)  &  (~ n540)  &  (~ n553) ) ;
 assign o_102_ =((~ i_0_) & i_0_);
 assign o_103_ =((~ i_0_) & i_0_);
 assign o_104_ =((~ i_0_) & i_0_);
 assign o_105_ =((~ i_0_) & i_0_);
 assign o_106_ =((~ i_0_) & i_0_);
 assign o_107_ =((~ i_0_) & i_0_);
 assign o_108_ =((~ i_0_) & i_0_);
 assign n11 = ( (~ o_92_)  &  (~ n189)  &  n451 ) | ( (~ o_92_)  &  n237  &  n451 ) ;
 assign n13 = ( n167  &  (~ n173) ) | ( n167  &  (~ n183) ) | ( (~ n173)  &  n237 ) | ( (~ n183)  &  n237 ) ;
 assign n14 = ( i_11_  &  n314 ) | ( n270  &  n314 ) | ( i_11_  &  (~ n519) ) | ( n270  &  (~ n519) ) ;
 assign n15 = ( i_21_  &  (~ n182) ) | ( n73  &  (~ n182) ) | ( i_21_  &  n299 ) | ( n73  &  n299 ) ;
 assign n16 = ( i_21_  &  n297 ) | ( (~ n178)  &  n297 ) ;
 assign n17 = ( (~ i_21_)  &  n295 ) | ( n73  &  n295 ) ;
 assign n18 = ( (~ n227)  &  n277 ) | ( n275  &  n277 ) | ( n277  &  n293 ) ;
 assign n19 = ( (~ i_22_)  &  n73 ) | ( n73  &  n195 ) | ( n73  &  n275 ) ;
 assign n20 = ( n186  &  n311 ) ;
 assign n21 = ( (~ o_22_)  &  n211  &  n273 ) | ( (~ o_22_)  &  n273  &  (~ n360) ) ;
 assign n22 = ( n67  &  n195 ) | ( n67  &  n196 ) | ( n67  &  n197 ) ;
 assign n24 = ( (~ i_9_) ) | ( (~ n245) ) | ( n305 ) ;
 assign n25 = ( i_9_ ) | ( (~ n186) ) | ( n303 ) ;
 assign n23 = ( n24  &  n25 ) ;
 assign n26 = ( i_12_  &  n192 ) | ( n192  &  n194 ) | ( i_12_  &  (~ n313) ) | ( n194  &  (~ n313) ) ;
 assign n27 = ( (~ i_11_)  &  n314 ) | ( n91  &  n314 ) | ( (~ i_11_)  &  (~ n439) ) | ( n91  &  (~ n439) ) ;
 assign n30 = ( i_11_  &  i_10_ ) ;
 assign n31 = ( i_10_  &  i_9_ ) ;
 assign n32 = ( (~ n184)  &  n199 ) | ( n196  &  n199 ) ;
 assign n33 = ( (~ i_20_)  &  n32 ) | ( i_21_  &  n32 ) | ( n32  &  n201 ) ;
 assign n34 = ( n203  &  n204  &  (~ n300) ) ;
 assign n35 = ( (~ n201)  &  n205 ) ;
 assign n36 = ( i_20_  &  (~ i_22_)  &  (~ n201) ) ;
 assign n37 = ( n204  &  n206  &  (~ n300) ) ;
 assign n38 = ( n189  &  n209 ) | ( n209  &  n207 ) | ( n209  &  (~ n597) ) ;
 assign n39 = ( i_22_  &  (~ n547) ) ;
 assign n42 = ( (~ o_19_)  &  n54  &  (~ n206) ) | ( (~ o_19_)  &  n54  &  n214 ) ;
 assign n44 = ( n221 ) | ( n222 ) | ( (~ n506) ) | ( (~ n598) ) ;
 assign n45 = ( n168  &  n225 ) ;
 assign n46 = ( i_9_ ) | ( n192 ) ;
 assign n47 = ( n219 ) | ( n220 ) | ( (~ n283) ) | ( (~ n288) ) | ( (~ n328) ) ;
 assign n43 = ( n44  &  n45  &  n46  &  n47 ) ;
 assign n49 = ( (~ i_21_) ) | ( n195 ) | ( (~ n414) ) ;
 assign n50 = ( n225 ) | ( i_10_ ) ;
 assign n51 = ( i_9_ ) | ( n168 ) ;
 assign n52 = ( i_22_ ) | ( n214 ) ;
 assign n48 = ( n49  &  n50  &  n51  &  n52 ) ;
 assign n54 = ( n225  &  n51  &  n49 ) ;
 assign n53 = ( n52  &  n54 ) ;
 assign n55 = ( (~ n195)  &  (~ n222)  &  n227 ) ;
 assign n56 = ( n179  &  (~ n540) ) ;
 assign n58 = ( n232 ) | ( n233 ) ;
 assign n59 = ( i_22_ ) | ( n228 ) | ( n229 ) | ( (~ n540) ) ;
 assign n60 = ( i_21_ ) | ( n230 ) | ( n231 ) | ( (~ n283) ) ;
 assign n57 = ( n58  &  n45  &  n59  &  n60 ) ;
 assign n62 = ( i_21_  &  (~ n547) ) ;
 assign n63 = ( (~ i_20_)  &  i_21_  &  n177 ) ;
 assign n65 = ( (~ n227) ) | ( n234 ) | ( n236 ) ;
 assign n66 = ( (~ n188) ) | ( n237 ) ;
 assign n67 = ( i_12_ ) | ( (~ n209) ) | ( (~ n311) ) ;
 assign n68 = ( (~ n204) ) | ( (~ n227) ) | ( n231 ) | ( n457 ) ;
 assign n64 = ( n65  &  n66  &  n67  &  n68 ) ;
 assign n69 = ( (~ i_10_)  &  (~ n263)  &  n267 ) | ( n94  &  (~ n263)  &  n267 ) ;
 assign n71 = ( (~ i_22_) ) | ( n268 ) | ( n269 ) ;
 assign n72 = ( (~ i_9_) ) | ( n270 ) ;
 assign n73 = ( i_20_ ) | ( n547 ) ;
 assign n74 = ( (~ i_20_) ) | ( n195 ) | ( n476 ) ;
 assign n70 = ( n71  &  n72  &  n73  &  n74 ) ;
 assign n75 = ( (~ o_96_)  &  n78  &  n291 ) | ( (~ o_96_)  &  n78  &  (~ n607) ) ;
 assign n77 = ( i_22_ ) | ( (~ n286) ) | ( n300 ) ;
 assign n78 = ( n289  &  n25  &  n290 ) ;
 assign n76 = ( (~ o_10_)  &  n74  &  n77  &  n78 ) ;
 assign n81 = ( n276  &  n277  &  n88  &  n278 ) ;
 assign n82 = ( (~ n178)  &  n273 ) ;
 assign n80 = ( n81  &  n82 ) ;
 assign n83 = ( (~ i_18_)  &  (~ i_19_)  &  n227  &  (~ n268) ) ;
 assign n85 = ( i_17_  &  (~ i_18_)  &  (~ n195)  &  n227 ) ;
 assign n87 = ( n276 ) | ( i_12_ ) ;
 assign n88 = ( n195 ) | ( n540 ) | ( n299 ) ;
 assign n86 = ( n82  &  n87  &  n88  &  (~ n661) ) ;
 assign n91 = ( i_9_ ) | ( n314 ) ;
 assign n94 = ( n561  &  n270 ) ;
 assign n90 = ( (~ o_7_)  &  n82  &  n91  &  n94  &  (~ n95) ) ;
 assign n95 = ( (~ i_10_)  &  n313  &  n493 ) ;
 assign n96 = ( (~ o_96_)  &  n94  &  n123  &  n308  &  n309 ) ;
 assign n97 = ( (~ i_10_)  &  n262  &  n313 ) ;
 assign n98 = ( i_1_  &  (~ n23) ) ;
 assign n99 = ( n360  &  n559 ) ;
 assign n100 = ( (~ i_8_)  &  i_12_  &  n310  &  n311 ) ;
 assign n101 = ( (~ o_75_)  &  n195 ) | ( (~ o_75_)  &  (~ n206) ) | ( (~ o_75_)  &  n269 ) ;
 assign n104 = ( n115  &  (~ n173)  &  n243 ) | ( n115  &  n239  &  n243 ) ;
 assign n105 = ( (~ n95)  &  n254  &  n255  &  n305  &  n322  &  n323 ) ;
 assign n108 = ( n240 ) | ( n247 ) | ( n252 ) ;
 assign n102 = ( (~ o_85_)  &  (~ o_96_)  &  n104  &  n105  &  n108  &  (~ n324) ) ;
 assign n111 = ( n240 ) | ( (~ n283) ) | ( (~ n328) ) ;
 assign n113 = ( i_10_ ) | ( (~ i_11_) ) | ( n330 ) ;
 assign n115 = ( n197  &  n240 ) | ( n239  &  n240 ) | ( n197  &  n241 ) | ( n239  &  n241 ) ;
 assign n116 = ( n240  &  n542 ) | ( n240  &  (~ n564) ) | ( n542  &  n565 ) | ( (~ n564)  &  n565 ) ;
 assign n109 = ( (~ o_92_)  &  n105  &  n111  &  n113  &  n115  &  n116  &  (~ n326)  &  (~ n331) ) ;
 assign n117 = ( n339  &  n340  &  n241 ) | ( n339  &  n340  &  n338 ) ;
 assign n119 = ( (~ i_21_) ) | ( n233 ) | ( (~ n380) ) ;
 assign n122 = ( (~ i_3_)  &  i_4_ ) | ( (~ i_3_)  &  n351 ) | ( i_4_  &  n577 ) | ( n351  &  n577 ) ;
 assign n123 = ( (~ n262)  &  n305 ) | ( n305  &  n303 ) ;
 assign n124 = ( (~ o_99_)  &  n345  &  n346  &  n347  &  n349  &  n350 ) ;
 assign n125 = ( (~ i_11_) ) | ( (~ n262) ) ;
 assign n118 = ( n94  &  n119  &  n122  &  n123  &  n124  &  n125  &  (~ n364)  &  (~ n367) ) ;
 assign n128 = ( i_10_  &  (~ n391) ) | ( i_10_  &  i_11_  &  n209 ) ;
 assign n130 = ( (~ n406)  &  (~ n524) ) | ( (~ n404)  &  (~ n524)  &  (~ n581) ) ;
 assign n131 = ( n227  &  (~ n400) ) | ( n227  &  n414  &  (~ n579) ) ;
 assign n132 = ( (~ i_4_)  &  (~ i_8_)  &  n311 ) ;
 assign n135 = ( (~ n206) ) | ( n457 ) | ( n486 ) ;
 assign n134 = ( n64  &  n135 ) ;
 assign n136 = ( (~ o_18_)  &  n13  &  n49  &  n433  &  n434  &  n435 ) ;
 assign n137 = ( n339  &  n440  &  n439 ) | ( n339  &  n440  &  n46 ) ;
 assign n138 = ( n448  &  n449  &  n442 ) | ( n448  &  n449  &  n300 ) ;
 assign n140 = ( (~ i_12_) ) | ( (~ n209) ) | ( (~ n246) ) ;
 assign n139 = ( (~ o_85_)  &  (~ o_96_)  &  n24  &  n140 ) ;
 assign n141 = ( (~ n262)  &  n471  &  n472 ) | ( n471  &  n472  &  n470 ) ;
 assign n142 = ( (~ i_4_)  &  (~ n473) ) | ( (~ i_4_)  &  (~ i_8_)  &  n188 ) ;
 assign n144 = ( n498  &  n502 ) | ( (~ n203)  &  n414  &  n502 ) ;
 assign n145 = ( (~ n484)  &  n497 ) | ( n407  &  (~ n484)  &  (~ n553) ) ;
 assign n147 = ( i_18_  &  n206  &  n283  &  (~ n591) ) ;
 assign n148 = ( (~ i_11_)  &  n506 ) | ( (~ n485)  &  n506 ) | ( n506  &  n505 ) ;
 assign n152 = ( (~ n371)  &  n427 ) ;
 assign n153 = ( (~ n209)  &  n347 ) | ( n347  &  n459 ) ;
 assign n154 = ( i_3_  &  n460 ) | ( n570  &  n460 ) | ( i_3_  &  n457 ) | ( n570  &  n457 ) ;
 assign n155 = ( (~ i_12_)  &  n231 ) | ( n231  &  (~ n262) ) | ( (~ i_12_)  &  n456 ) | ( (~ n262)  &  n456 ) ;
 assign n156 = ( (~ o_99_)  &  n330  &  n461  &  n465  &  n466  &  (~ n467)  &  n571  &  n572 ) ;
 assign n151 = ( n94  &  n152  &  n153  &  n154  &  n155  &  n156 ) ;
 assign n157 = ( (~ n444)  &  n502 ) | ( n502  &  n513 ) | ( n502  &  (~ n596) ) ;
 assign n158 = ( (~ n484)  &  n512 ) | ( (~ n484)  &  n514  &  (~ n553) ) ;
 assign n159 = ( (~ n356)  &  (~ n591) ) | ( (~ n591)  &  (~ n646) ) ;
 assign n160 = ( (~ i_4_)  &  (~ n647) ) | ( (~ i_4_)  &  n518  &  n519 ) ;
 assign n161 = ( n209  &  (~ n311) ) ;
 assign n167 = ( (~ i_11_) ) | ( (~ n246) ) ;
 assign n168 = ( i_12_ ) | ( (~ n506) ) ;
 assign n166 = ( n167 ) | ( n168 ) ;
 assign n171 = ( (~ i_18_)  &  (~ i_19_)  &  i_20_ ) ;
 assign n173 = ( (~ i_20_)  &  n203 ) ;
 assign n177 = ( (~ n293)  &  (~ n553) ) ;
 assign n178 = ( i_20_  &  (~ n195)  &  (~ n553) ) ;
 assign n179 = ( (~ n293)  &  (~ n549) ) ;
 assign n180 = ( (~ i_20_)  &  n206 ) ;
 assign n182 = ( n173  &  (~ n195) ) ;
 assign n183 = ( (~ n222)  &  (~ n293) ) ;
 assign n184 = ( n180  &  (~ n195) ) ;
 assign n185 = ( i_17_  &  i_18_  &  (~ i_19_) ) ;
 assign n186 = ( (~ i_8_)  &  n493 ) ;
 assign n188 = ( (~ i_9_)  &  n30 ) ;
 assign n189 = ( i_9_  &  n541 ) ;
 assign n191 = ( i_10_  &  (~ i_11_) ) ;
 assign n192 = ( (~ i_10_) ) | ( (~ n506) ) ;
 assign n194 = ( (~ n311) ) | ( (~ n506) ) ;
 assign n195 = ( n534 ) | ( n475 ) | ( n474 ) ;
 assign n196 = ( i_19_ ) | ( n536 ) ;
 assign n197 = ( (~ i_22_) ) | ( n540 ) ;
 assign n199 = ( i_12_  &  (~ o_85_) ) | ( (~ o_85_)  &  (~ n209) ) | ( (~ o_85_)  &  (~ n246) ) ;
 assign n201 = ( n293 ) | ( n196 ) ;
 assign n203 = ( (~ i_21_)  &  i_22_ ) ;
 assign n204 = ( i_18_  &  (~ i_19_)  &  i_20_ ) ;
 assign n205 = ( i_22_  &  i_20_ ) ;
 assign n206 = ( (~ i_21_)  &  (~ i_22_) ) ;
 assign n209 = ( (~ i_8_)  &  n532 ) ;
 assign n207 = ( (~ i_9_)  &  n191 ) ;
 assign n211 = ( i_18_ ) | ( (~ i_22_) ) | ( n268 ) ;
 assign n210 = ( i_20_  &  (~ n83) ) | ( (~ n83)  &  n211 ) ;
 assign n214 = ( n300 ) | ( (~ n453) ) ;
 assign n219 = ( (~ i_8_) ) | ( (~ n30) ) ;
 assign n220 = ( i_15_ ) | ( n487 ) ;
 assign n221 = ( i_13_ ) | ( (~ n30) ) ;
 assign n222 = ( (~ i_19_) ) | ( n536 ) ;
 assign n225 = ( i_9_ ) | ( i_11_ ) | ( (~ n506) ) ;
 assign n227 = ( i_22_  &  i_21_ ) ;
 assign n228 = ( (~ i_19_) ) | ( n194 ) | ( n220 ) ;
 assign n229 = ( i_16_ ) | ( n536 ) ;
 assign n230 = ( (~ i_18_) ) | ( n233 ) ;
 assign n231 = ( i_17_ ) | ( n531 ) ;
 assign n232 = ( (~ i_21_) ) | ( n234 ) ;
 assign n233 = ( (~ i_11_) ) | ( n487 ) | ( n534 ) ;
 assign n234 = ( n231 ) | ( (~ n453) ) ;
 assign n236 = ( (~ n310) ) | ( n437 ) ;
 assign n237 = ( (~ i_12_) ) | ( (~ n506) ) ;
 assign n239 = ( n549 ) | ( n558 ) ;
 assign n240 = ( n534 ) | ( n220 ) ;
 assign n241 = ( (~ i_21_) ) | ( n229 ) | ( (~ n360) ) ;
 assign n243 = ( (~ o_99_)  &  (~ n180) ) | ( (~ o_99_)  &  n229 ) | ( (~ o_99_)  &  n240 ) ;
 assign n245 = ( i_12_  &  i_11_ ) ;
 assign n246 = ( (~ i_9_)  &  (~ i_10_) ) ;
 assign n244 = ( n167  &  n245 ) | ( n167  &  n246 ) ;
 assign n249 = ( i_21_ ) | ( n248 ) ;
 assign n248 = ( i_19_ ) | ( i_20_ ) ;
 assign n247 = ( n249  &  i_22_ ) | ( n249  &  n248 ) ;
 assign n251 = ( i_16_ ) | ( n548 ) ;
 assign n252 = ( i_16_ ) | ( (~ i_17_) ) | ( (~ i_18_) ) ;
 assign n250 = ( n247  &  n252 ) | ( n251  &  n252 ) | ( n247  &  n249 ) | ( n251  &  n249 ) ;
 assign n254 = ( n554 ) | ( n555 ) ;
 assign n255 = ( n508 ) | ( n240 ) | ( i_19_ ) | ( n229 ) ;
 assign n256 = ( (~ n206)  &  n600 ) | ( n222  &  n600 ) | ( n558  &  n600 ) ;
 assign n257 = ( (~ i_12_) ) | ( n167 ) | ( (~ n186) ) ;
 assign n258 = ( (~ n325) ) | ( n459 ) ;
 assign n259 = ( n239  &  n601 ) | ( (~ n514)  &  n601 ) ;
 assign n253 = ( n254  &  n255  &  n111  &  n256  &  n257  &  n104  &  n258  &  n259 ) ;
 assign n262 = ( (~ i_9_)  &  n493 ) ;
 assign n261 = ( n245  &  i_10_ ) ;
 assign n260 = ( n262  &  n261 ) | ( (~ i_12_)  &  n191  &  n262 ) ;
 assign n263 = ( i_21_  &  n99 ) | ( i_21_  &  (~ n195)  &  (~ n476) ) ;
 assign n267 = ( (~ n260)  &  (~ n379)  &  n604 ) | ( (~ n260)  &  (~ n559)  &  n604 ) ;
 assign n268 = ( n544 ) | ( n545 ) ;
 assign n269 = ( i_18_ ) | ( n248 ) ;
 assign n270 = ( i_12_ ) | ( n314 ) ;
 assign n273 = ( i_22_ ) | ( n268 ) | ( (~ n286) ) ;
 assign n275 = ( i_20_ ) | ( n299 ) ;
 assign n276 = ( (~ i_9_) ) | ( (~ i_10_) ) | ( (~ n186) ) ;
 assign n277 = ( (~ n227) ) | ( n293 ) | ( n546 ) ;
 assign n278 = ( (~ i_22_)  &  (~ n661) ) | ( n275  &  (~ n661) ) | ( n293  &  (~ n661) ) ;
 assign n280 = ( n195  &  (~ n380) ) | ( (~ n286)  &  (~ n380) ) | ( n195  &  n544 ) | ( (~ n286)  &  n544 ) ;
 assign n281 = ( (~ o_10_)  &  (~ n186)  &  n605 ) | ( (~ o_10_)  &  n303  &  n605 ) ;
 assign n279 = ( n280  &  n81  &  n281 ) ;
 assign n283 = ( i_20_  &  i_19_ ) ;
 assign n282 = ( i_22_  &  n283  &  (~ n560) ) ;
 assign n288 = ( (~ i_1_)  &  n532 ) ;
 assign n286 = ( (~ i_18_)  &  n283 ) ;
 assign n285 = ( n282  &  n288 ) | ( (~ n231)  &  n288  &  n286 ) ;
 assign n289 = ( (~ i_9_) ) | ( n561 ) ;
 assign n290 = ( (~ i_9_)  &  (~ i_12_) ) | ( (~ i_9_)  &  n427 ) | ( (~ i_12_)  &  n606 ) | ( n427  &  n606 ) ;
 assign n291 = ( (~ i_12_) ) | ( n487 ) ;
 assign n293 = ( n475 ) | ( n539 ) ;
 assign n295 = ( n195 ) | ( (~ n227) ) | ( n275 ) ;
 assign n297 = ( (~ n206) ) | ( n268 ) | ( (~ n286) ) ;
 assign n299 = ( (~ i_17_) ) | ( i_18_ ) ;
 assign n300 = ( n544 ) | ( n231 ) ;
 assign n305 = ( i_10_ ) | ( n314 ) ;
 assign n303 = ( (~ i_10_) ) | ( (~ i_12_) ) ;
 assign n306 = ( i_16_  &  (~ i_19_) ) | ( i_16_  &  n251 ) | ( (~ i_19_)  &  (~ n286) ) | ( n251  &  (~ n286) ) ;
 assign n308 = ( (~ n288) ) | ( n291 ) | ( (~ n311) ) | ( n486 ) ;
 assign n309 = ( i_22_ ) | ( n220 ) | ( (~ n261) ) | ( n306 ) | ( (~ n563) ) ;
 assign n310 = ( n532  &  i_1_ ) ;
 assign n311 = ( i_9_  &  n30 ) ;
 assign n313 = ( (~ i_11_)  &  i_12_ ) ;
 assign n314 = ( (~ i_8_) ) | ( (~ n493) ) ;
 assign n318 = ( i_12_  &  i_11_ ) | ( i_12_  &  n246 ) ;
 assign n319 = ( i_17_  &  (~ n286) ) | ( (~ i_19_)  &  (~ n286) ) | ( (~ n286)  &  (~ n540) ) ;
 assign n320 = ( i_17_  &  i_22_ ) | ( i_17_  &  n319 ) | ( i_22_  &  (~ n423) ) | ( n319  &  (~ n423) ) ;
 assign n322 = ( (~ i_12_)  &  n320 ) | ( (~ n262)  &  n320 ) | ( (~ i_12_)  &  n558 ) | ( (~ n262)  &  n558 ) ;
 assign n323 = ( i_4_  &  n593 ) | ( (~ i_8_)  &  n593 ) | ( n318  &  n593 ) ;
 assign n326 = ( n191  &  n563 ) ;
 assign n325 = ( (~ i_9_)  &  n532 ) ;
 assign n324 = ( (~ i_12_)  &  n326 ) | ( (~ i_10_)  &  (~ i_12_)  &  n325 ) ;
 assign n328 = ( (~ i_21_)  &  (~ n229) ) ;
 assign n327 = ( i_19_  &  (~ i_20_)  &  n328 ) ;
 assign n330 = ( i_4_ ) | ( (~ i_8_) ) | ( i_9_ ) ;
 assign n331 = ( n327  &  (~ n555) ) | ( (~ n249)  &  (~ n251)  &  (~ n555) ) ;
 assign n335 = ( n231 ) | ( n236 ) | ( n269 ) | ( (~ n407) ) ;
 assign n337 = ( (~ n506) ) | ( (~ n519) ) ;
 assign n339 = ( n68  &  n135  &  n67  &  n571  &  n572  &  n335  &  n337 ) ;
 assign n340 = ( n46  &  n589 ) | ( n46  &  n570 ) ;
 assign n338 = ( n220 ) | ( (~ n261) ) | ( (~ n506) ) ;
 assign n343 = ( i_19_ ) | ( n545 ) ;
 assign n341 = ( (~ n180)  &  n343 ) | ( n231  &  n343 ) | ( (~ n180)  &  (~ n514) ) | ( n231  &  (~ n514) ) ;
 assign n345 = ( i_4_ ) | ( (~ n439) ) | ( n533 ) ;
 assign n346 = ( i_0_ ) | ( (~ i_1_) ) | ( (~ i_20_) ) | ( (~ n407) ) | ( n475 ) | ( n548 ) | ( n574 ) ;
 assign n347 = ( i_10_ ) | ( (~ n468) ) ;
 assign n349 = ( n230  &  n330 ) | ( n330  &  n341 ) | ( n230  &  (~ n541) ) | ( n341  &  (~ n541) ) ;
 assign n350 = ( n613  &  n228 ) | ( n613  &  n523 ) ;
 assign n353 = ( (~ i_8_)  &  n612 ) | ( n459  &  n543  &  n612 ) ;
 assign n351 = ( (~ n313)  &  n353 ) | ( n353  &  (~ n518) ) ;
 assign n355 = ( (~ i_11_) ) | ( n487 ) | ( n537 ) ;
 assign n354 = ( (~ i_20_)  &  n269 ) | ( n230  &  n269 ) | ( (~ i_20_)  &  n355 ) | ( n230  &  n355 ) ;
 assign n357 = ( (~ i_18_) ) | ( (~ i_20_) ) ;
 assign n356 = ( i_21_  &  (~ n206) ) | ( (~ n204)  &  (~ n206) ) | ( i_21_  &  n357 ) | ( (~ n204)  &  n357 ) ;
 assign n360 = ( i_19_  &  (~ i_20_) ) ;
 assign n359 = ( (~ n355)  &  (~ n356) ) | ( (~ i_22_)  &  (~ n355)  &  n360 ) ;
 assign n364 = ( (~ n231)  &  (~ n609) ) | ( n203  &  (~ n231)  &  (~ n354) ) ;
 assign n367 = ( n209  &  (~ n611) ) | ( (~ i_10_)  &  n209  &  (~ n245) ) ;
 assign n371 = ( n191  &  n262 ) | ( (~ i_10_)  &  i_11_  &  n262 ) ;
 assign n372 = ( (~ i_19_)  &  i_21_ ) | ( i_21_  &  (~ n206) ) | ( (~ i_19_)  &  n269 ) | ( (~ n206)  &  n269 ) ;
 assign n374 = ( (~ n204) ) | ( n233 ) | ( (~ n407) ) ;
 assign n375 = ( (~ n203) ) | ( n230 ) | ( (~ n283) ) ;
 assign n373 = ( n374  &  n375  &  n372 ) | ( n374  &  n375  &  n355 ) ;
 assign n377 = ( (~ i_9_) ) | ( i_11_ ) ;
 assign n376 = ( i_9_  &  (~ n313)  &  n377 ) | ( n303  &  (~ n313)  &  n377 ) ;
 assign n380 = ( (~ i_22_)  &  n283  &  (~ n560) ) ;
 assign n379 = ( i_19_  &  n407 ) ;
 assign n378 = ( (~ n355)  &  n380 ) | ( (~ n355)  &  n379  &  (~ n560) ) ;
 assign n382 = ( n508 ) | ( n228 ) | ( i_16_ ) | ( i_18_ ) ;
 assign n384 = ( n615  &  i_2_ ) | ( n615  &  n577  &  n617 ) ;
 assign n385 = ( n231  &  (~ n313) ) | ( (~ n313)  &  n373 ) | ( n231  &  (~ n563) ) | ( n373  &  (~ n563) ) ;
 assign n386 = ( (~ n209)  &  n459 ) | ( n376  &  n459 ) | ( (~ n209)  &  (~ n532) ) | ( n376  &  (~ n532) ) ;
 assign n387 = ( n124  &  n152  &  (~ n262) ) | ( n124  &  n152  &  (~ n439) ) ;
 assign n381 = ( (~ n20)  &  n27  &  n289  &  n382  &  n384  &  n385  &  n386  &  n387 ) ;
 assign n389 = ( i_2_ ) | ( (~ i_3_) ) | ( n567 ) ;
 assign n390 = ( (~ n206) ) | ( n536 ) ;
 assign n388 = ( n389  &  n390  &  i_21_ ) | ( n389  &  n390  &  n196 ) ;
 assign n392 = ( n475 ) | ( n197 ) | ( n549 ) ;
 assign n391 = ( i_0_ ) | ( (~ i_1_) ) | ( i_3_ ) | ( i_13_ ) | ( n237 ) | ( n392 ) ;
 assign n396 = ( n620  &  i_20_ ) | ( n620  &  n523 ) | ( n620  &  n581 ) ;
 assign n395 = ( (~ n288) ) | ( n580 ) ;
 assign n393 = ( (~ n205)  &  n396 ) | ( n229  &  n396 ) | ( n396  &  n395 ) ;
 assign n397 = ( i_9_  &  (~ n519) ) | ( i_11_  &  (~ n519) ) | ( i_12_  &  (~ n519) ) ;
 assign n399 = ( i_6_ ) | ( n542 ) | ( (~ n564) ) ;
 assign n398 = ( n24  &  (~ n209)  &  n399 ) | ( n24  &  n397  &  n399 ) ;
 assign n401 = ( (~ n171) ) | ( n231 ) | ( n291 ) ;
 assign n403 = ( i_4_ ) | ( n566 ) ;
 assign n400 = ( (~ i_1_) ) | ( (~ i_2_) ) | ( n401 ) | ( n403 ) ;
 assign n404 = ( i_22_  &  (~ n379) ) | ( (~ n283)  &  (~ n379) ) ;
 assign n407 = ( i_21_  &  (~ i_22_) ) ;
 assign n406 = ( (~ n283) ) | ( n395 ) | ( n407 ) ;
 assign n414 = ( (~ i_20_)  &  (~ n222) ) ;
 assign n417 = ( n395 ) | ( n241 ) ;
 assign n418 = ( (~ i_1_)  &  (~ n575) ) | ( (~ i_3_)  &  (~ n575) ) ;
 assign n421 = ( i_18_  &  (~ n180) ) | ( i_22_  &  (~ n180) ) ;
 assign n423 = ( (~ i_18_)  &  n514 ) ;
 assign n422 = ( (~ i_17_)  &  n423 ) | ( (~ i_17_)  &  i_18_  &  n180 ) ;
 assign n425 = ( (~ n195)  &  n422 ) | ( (~ n195)  &  n286  &  n407 ) ;
 assign n427 = ( (~ n189) ) | ( (~ n493) ) ;
 assign n428 = ( (~ i_19_)  &  n623 ) | ( n300  &  n623 ) | ( n421  &  n623 ) ;
 assign n429 = ( (~ i_6_)  &  (~ n262) ) | ( (~ i_6_)  &  n480 ) | ( (~ n262)  &  n587 ) | ( n480  &  n587 ) ;
 assign n430 = ( i_10_  &  (~ n425) ) | ( n245  &  (~ n425) ) | ( n330  &  (~ n425) ) ;
 assign n431 = ( (~ n173) ) | ( (~ n179) ) ;
 assign n426 = ( (~ o_7_)  &  (~ o_99_)  &  n94  &  n427  &  n428  &  n429  &  n430  &  n431 ) ;
 assign n433 = ( i_1_ ) | ( n588 ) ;
 assign n434 = ( n214  &  n588 ) | ( (~ n407)  &  n588 ) | ( n214  &  n589 ) | ( (~ n407)  &  n589 ) ;
 assign n435 = ( n245 ) | ( n46 ) ;
 assign n438 = ( n541 ) | ( n330 ) ;
 assign n437 = ( n291 ) | ( n219 ) ;
 assign n436 = ( n438  &  i_4_ ) | ( n438  &  n232 ) | ( n438  &  n437 ) ;
 assign n440 = ( n626  &  i_22_ ) | ( n626  &  n241 ) | ( n626  &  n338 ) ;
 assign n439 = ( i_11_  &  (~ i_12_) ) ;
 assign n441 = ( (~ i_19_)  &  (~ n514) ) | ( i_22_  &  (~ n514) ) ;
 assign n443 = ( (~ i_22_)  &  (~ n206) ) | ( (~ i_22_)  &  (~ n283) ) | ( (~ n206)  &  (~ n360) ) | ( (~ n283)  &  (~ n360) ) ;
 assign n442 = ( i_21_  &  n443 ) | ( (~ n204)  &  n443 ) ;
 assign n444 = ( (~ i_20_)  &  n390 ) | ( n196  &  n390 ) ;
 assign n445 = ( i_17_  &  n444 ) | ( (~ i_19_)  &  n444 ) | ( n444  &  (~ n508) ) ;
 assign n447 = ( n186  &  n207 ) | ( (~ i_12_)  &  n186  &  n189 ) ;
 assign n448 = ( (~ n179)  &  n441 ) | ( (~ n203)  &  n441 ) | ( (~ n179)  &  (~ n559) ) | ( (~ n203)  &  (~ n559) ) ;
 assign n449 = ( n25  &  n195  &  (~ n447) ) | ( n25  &  n445  &  (~ n447) ) ;
 assign n451 = ( n556 ) | ( n459 ) ;
 assign n453 = ( i_18_  &  n360 ) ;
 assign n452 = ( (~ n236)  &  (~ n631) ) | ( (~ i_21_)  &  (~ n236)  &  n453 ) ;
 assign n457 = ( (~ n288) ) | ( n437 ) ;
 assign n456 = ( (~ i_21_)  &  (~ n452) ) | ( (~ n204)  &  (~ n452) ) | ( (~ n452)  &  n457 ) ;
 assign n459 = ( i_10_ ) | ( (~ n439) ) ;
 assign n460 = ( (~ i_18_)  &  n232  &  (~ n380) ) | ( n232  &  n341  &  (~ n380) ) ;
 assign n463 = ( n220 ) | ( n554 ) ;
 assign n461 = ( (~ i_1_) ) | ( (~ n261) ) | ( n463 ) | ( (~ n506) ) | ( (~ n630) ) ;
 assign n465 = ( n251 ) | ( n441 ) | ( n338 ) ;
 assign n466 = ( i_4_ ) | ( i_9_ ) | ( (~ n313) ) ;
 assign n468 = ( i_9_  &  n209 ) ;
 assign n467 = ( (~ i_12_)  &  n468 ) | ( i_6_  &  (~ i_11_)  &  n468 ) ;
 assign n471 = ( n245  &  n634 ) | ( (~ n468)  &  n634 ) ;
 assign n472 = ( n94  &  n153  &  n313 ) | ( n94  &  n153  &  n330 ) ;
 assign n470 = ( (~ i_10_) ) | ( (~ n439) ) ;
 assign n474 = ( i_13_ ) | ( (~ n245) ) ;
 assign n475 = ( i_14_ ) | ( n531 ) ;
 assign n476 = ( (~ i_19_) ) | ( n548 ) ;
 assign n478 = ( (~ i_10_) ) | ( n533 ) ;
 assign n473 = ( (~ i_7_) ) | ( i_22_ ) | ( n474 ) | ( n475 ) | ( n476 ) | ( n478 ) ;
 assign n480 = ( (~ i_12_)  &  n541 ) ;
 assign n479 = ( i_9_  &  (~ n189) ) | ( (~ n189)  &  n480 ) ;
 assign n484 = ( (~ i_8_) ) | ( (~ n310) ) | ( n557 ) ;
 assign n482 = ( (~ n20)  &  n407 ) | ( (~ n20)  &  (~ n414) ) | ( (~ n20)  &  n484 ) ;
 assign n486 = ( (~ n286) ) | ( n545 ) ;
 assign n487 = ( i_14_ ) | ( i_13_ ) ;
 assign n485 = ( (~ i_10_) ) | ( i_22_ ) | ( n486 ) | ( n487 ) ;
 assign n489 = ( i_19_ ) | ( (~ n203) ) | ( n566 ) | ( n583 ) ;
 assign n488 = ( (~ i_8_)  &  (~ n188)  &  n489 ) | ( i_11_  &  (~ n188)  &  n489 ) ;
 assign n493 = ( (~ i_4_)  &  (~ i_7_) ) ;
 assign n490 = ( (~ n479)  &  n493 ) | ( n493  &  (~ n643) ) ;
 assign n496 = ( n220  &  n644 ) | ( n403  &  n644 ) | ( (~ n641)  &  n644 ) ;
 assign n494 = ( i_4_  &  (~ n490)  &  n496 ) | ( n488  &  (~ n490)  &  n496 ) ;
 assign n497 = ( n180  &  (~ n549) ) | ( (~ n508)  &  (~ n549) ) ;
 assign n498 = ( i_20_  &  (~ n638) ) | ( i_20_  &  (~ n222)  &  (~ n407) ) ;
 assign n502 = ( i_8_  &  n288  &  (~ n557) ) ;
 assign n506 = ( n532  &  i_8_ ) ;
 assign n505 = ( (~ i_9_)  &  i_12_ ) | ( i_9_  &  (~ i_12_) ) ;
 assign n508 = ( i_22_ ) | ( n540 ) ;
 assign n507 = ( i_1_ ) | ( (~ i_10_) ) | ( n196 ) | ( n474 ) | ( n475 ) | ( n508 ) ;
 assign n510 = ( (~ i_8_)  &  (~ n30) ) | ( i_8_  &  (~ n507) ) | ( (~ n30)  &  (~ n507) ) ;
 assign n511 = ( (~ i_10_)  &  n532 ) | ( n532  &  n543 ) ;
 assign n509 = ( n510  &  n397  &  n511 ) ;
 assign n512 = ( (~ n540)  &  (~ n549) ) | ( (~ i_20_)  &  (~ n227)  &  (~ n549) ) ;
 assign n514 = ( (~ i_20_)  &  n407 ) ;
 assign n513 = ( n514  &  n185 ) ;
 assign n518 = ( (~ i_8_)  &  (~ i_10_) ) ;
 assign n519 = ( (~ i_9_)  &  n245 ) ;
 assign n523 = ( i_22_ ) | ( n251 ) ;
 assign n524 = ( i_16_ ) | ( n299 ) ;
 assign n522 = ( n249  &  n404 ) | ( n523  &  n404 ) | ( n249  &  n524 ) | ( n523  &  n524 ) ;
 assign n526 = ( n522 ) | ( n555 ) ;
 assign n527 = ( n537 ) | ( n576 ) | ( n658 ) | ( n659 ) ;
 assign n528 = ( (~ n209)  &  n398 ) | ( (~ n261)  &  n398 ) ;
 assign n529 = ( (~ i_22_)  &  n245 ) | ( (~ i_22_)  &  n556 ) | ( n245  &  n593 ) | ( n556  &  n593 ) ;
 assign n525 = ( (~ o_92_)  &  (~ n20)  &  n526  &  n527  &  n528  &  n529 ) ;
 assign n530 = ( i_1_  &  i_2_ ) | ( (~ i_1_)  &  (~ i_2_) ) ;
 assign n531 = ( i_16_ ) | ( i_15_ ) ;
 assign n532 = ( (~ i_4_)  &  i_7_ ) ;
 assign n533 = ( (~ i_8_) ) | ( (~ i_9_) ) ;
 assign n534 = ( (~ n288) ) | ( n478 ) ;
 assign n536 = ( i_17_ ) | ( (~ i_18_) ) ;
 assign n537 = ( (~ n310) ) | ( n478 ) ;
 assign n539 = ( n474 ) | ( n537 ) ;
 assign n540 = ( (~ i_20_) ) | ( (~ i_21_) ) ;
 assign n541 = ( (~ i_10_)  &  (~ i_11_) ) ;
 assign n542 = ( (~ i_10_) ) | ( (~ n209) ) ;
 assign n543 = ( (~ i_9_) ) | ( (~ n313) ) ;
 assign n544 = ( n194 ) | ( n291 ) ;
 assign n545 = ( (~ i_17_) ) | ( n531 ) ;
 assign n546 = ( i_19_ ) | ( n299 ) ;
 assign n547 = ( n195 ) | ( n546 ) ;
 assign n548 = ( i_17_ ) | ( i_18_ ) ;
 assign n549 = ( i_19_ ) | ( n548 ) ;
 assign n553 = ( (~ i_19_) ) | ( n299 ) ;
 assign n554 = ( i_19_ ) | ( n540 ) | ( n251 ) ;
 assign n555 = ( n537 ) | ( n220 ) ;
 assign n556 = ( (~ i_9_) ) | ( (~ n506) ) ;
 assign n557 = ( (~ i_10_) ) | ( i_13_ ) | ( n475 ) ;
 assign n558 = ( n556 ) | ( n557 ) ;
 assign n559 = ( (~ i_18_)  &  (~ n300) ) ;
 assign n560 = ( i_18_ ) | ( n531 ) ;
 assign n561 = ( i_11_ ) | ( n314 ) ;
 assign n563 = ( n532  &  i_9_ ) ;
 assign n564 = ( i_12_  &  i_9_ ) ;
 assign n565 = ( i_19_ ) | ( n252 ) | ( (~ n514) ) ;
 assign n566 = ( (~ i_7_) ) | ( (~ i_8_) ) | ( (~ i_10_) ) ;
 assign n567 = ( i_1_ ) | ( i_17_ ) | ( i_19_ ) | ( (~ n227) ) ;
 assign n568 = ( n474 ) | ( n403 ) ;
 assign n570 = ( (~ i_2_) ) | ( n392 ) | ( n568 ) ;
 assign n571 = ( (~ i_2_) ) | ( (~ i_20_) ) | ( n475 ) | ( n567 ) | ( n568 ) ;
 assign n572 = ( (~ i_22_) ) | ( n234 ) | ( n236 ) ;
 assign n573 = ( (~ i_7_) ) | ( n533 ) ;
 assign n574 = ( i_4_ ) | ( n221 ) | ( n573 ) ;
 assign n575 = ( i_1_  &  i_0_ ) ;
 assign n576 = ( (~ i_22_) ) | ( n463 ) ;
 assign n577 = ( n194 ) | ( (~ n575) ) | ( n576 ) ;
 assign n579 = ( n237 ) | ( n557 ) ;
 assign n580 = ( (~ i_8_) ) | ( n220 ) | ( n303 ) ;
 assign n581 = ( (~ n310) ) | ( n580 ) ;
 assign n583 = ( (~ i_1_) ) | ( n220 ) | ( n251 ) ;
 assign n584 = ( i_4_ ) | ( (~ n261) ) | ( n573 ) ;
 assign n585 = ( n194 ) | ( (~ n227) ) | ( n401 ) ;
 assign n587 = ( n542 ) | ( n543 ) ;
 assign n588 = ( (~ i_2_) ) | ( n576 ) | ( n584 ) ;
 assign n589 = ( i_3_  &  i_0_ ) ;
 assign n590 = ( n539 ) | ( n392 ) ;
 assign n591 = ( n192 ) | ( n487 ) | ( n231 ) ;
 assign n593 = ( n240 ) | ( (~ n283) ) | ( n524 ) ;
 assign n594 = ( i_3_  &  n653 ) | ( (~ n575)  &  n653 ) | ( n585  &  n653 ) ;
 assign n595 = ( i_2_  &  n655 ) | ( (~ n589)  &  n655 ) | ( n590  &  n655 ) ;
 assign n596 = ( (~ i_21_)  &  n657 ) | ( (~ n414)  &  n657 ) ;
 assign n597 = ( (~ i_12_)  &  n543 ) | ( n167  &  n543 ) ;
 assign n598 = ( n206  &  (~ n475) ) | ( (~ i_20_)  &  (~ n203)  &  (~ n475) ) ;
 assign n600 = ( n227 ) | ( n229 ) | ( (~ n360) ) | ( n555 ) ;
 assign n601 = ( n240  &  n244 ) | ( n244  &  n250 ) | ( n240  &  (~ n506) ) | ( n250  &  (~ n506) ) ;
 assign n604 = ( i_22_ ) | ( (~ n178) ) ;
 assign n606 = ( n305  &  n270 ) ;
 assign n605 = ( (~ i_9_)  &  (~ n493) ) | ( (~ i_9_)  &  n543 ) | ( (~ n493)  &  n606 ) | ( n543  &  n606 ) ;
 assign n607 = ( n311  &  n285 ) | ( n311  &  n380  &  n310 ) ;
 assign n609 = ( i_22_  &  (~ n359) ) | ( (~ n204)  &  (~ n359) ) | ( n233  &  (~ n359) ) ;
 assign n611 = ( i_11_  &  (~ n261) ) | ( (~ i_6_)  &  (~ n261)  &  n564 ) ;
 assign n612 = ( n392 ) | ( n573 ) | ( n530 ) | ( n221 ) ;
 assign n613 = ( n231 ) | ( n233 ) | ( (~ n423) ) ;
 assign n615 = ( (~ i_22_)  &  (~ n378) ) | ( n233  &  (~ n378) ) | ( (~ n378)  &  n486 ) ;
 assign n617 = ( (~ i_3_) ) | ( n392 ) | ( n574 ) ;
 assign n620 = ( i_18_ ) | ( n231 ) | ( n291 ) | ( n403 ) | ( (~ n407) ) | ( (~ n575) ) ;
 assign n621 = ( (~ i_20_)  &  n46 ) | ( n46  &  n388 ) | ( n46  &  n579 ) ;
 assign n622 = ( i_11_  &  i_19_ ) | ( n556  &  i_19_ ) | ( i_11_  &  n393 ) | ( n556  &  n393 ) ;
 assign n624 = ( n583 ) | ( n584 ) | ( i_0_ ) | ( n508 ) ;
 assign n623 = ( n624  &  i_2_ ) | ( n624  &  n418 ) | ( n624  &  n585 ) ;
 assign n627 = ( (~ n407) ) | ( n475 ) | ( n549 ) | ( n568 ) | ( (~ n575) ) ;
 assign n626 = ( (~ i_0_)  &  n627 ) | ( (~ i_7_)  &  n627 ) | ( n436  &  n627 ) ;
 assign n630 = ( (~ i_0_)  &  i_3_ ) | ( (~ i_2_)  &  i_3_ ) | ( (~ i_0_)  &  n575 ) | ( (~ i_2_)  &  n575 ) ;
 assign n631 = ( i_18_  &  (~ n203) ) | ( i_18_  &  n269 ) | ( (~ n203)  &  (~ n407) ) | ( n269  &  (~ n407) ) ;
 assign n634 = ( i_10_ ) | ( (~ i_12_) ) | ( (~ n186) ) ;
 assign n637 = ( n220 ) | ( n584 ) | ( n650 ) | ( n651 ) ;
 assign n636 = ( (~ i_8_)  &  (~ n245) ) | ( (~ i_8_)  &  (~ n518) ) | ( n245  &  (~ n518) ) ;
 assign n635 = ( (~ n493)  &  n637 ) | ( n479  &  n637  &  n636 ) ;
 assign n638 = ( (~ n227)  &  n553 ) | ( n536  &  n553 ) ;
 assign n639 = ( (~ i_19_)  &  n565 ) | ( n251  &  n565 ) ;
 assign n641 = ( (~ i_1_)  &  (~ n639) ) | ( (~ i_1_)  &  n180  &  (~ n229) ) ;
 assign n643 = ( (~ i_8_)  &  (~ i_12_) ) | ( (~ i_8_)  &  (~ n518) ) | ( (~ i_12_)  &  n564 ) | ( (~ n518)  &  n564 ) ;
 assign n644 = ( n205 ) | ( n476 ) | ( (~ n506) ) | ( n557 ) ;
 assign n645 = ( i_5_  &  n470 ) | ( n470  &  n494 ) | ( i_5_  &  (~ n563) ) | ( n494  &  (~ n563) ) ;
 assign n646 = ( (~ n171)  &  n269 ) | ( (~ n227)  &  n269 ) | ( (~ n171)  &  (~ n407) ) | ( (~ n227)  &  (~ n407) ) ;
 assign n647 = ( (~ i_7_)  &  i_8_ ) | ( i_8_  &  i_12_ ) | ( (~ i_7_)  &  n470 ) | ( i_12_  &  n470 ) ;
 assign n648 = ( i_11_  &  (~ n325) ) | ( i_11_  &  n541 ) | ( (~ n325)  &  (~ n563) ) | ( n541  &  (~ n563) ) ;
 assign n650 = ( i_1_  &  (~ i_22_) ) | ( i_1_  &  n249 ) | ( i_1_  &  n251 ) ;
 assign n652 = ( i_22_ ) | ( n229 ) | ( n249 ) ;
 assign n651 = ( (~ i_1_)  &  n565  &  n652 ) ;
 assign n653 = ( (~ i_3_) ) | ( n575 ) | ( n576 ) | ( n584 ) ;
 assign n655 = ( (~ i_2_) ) | ( i_3_ ) | ( n575 ) | ( n585 ) ;
 assign n657 = ( (~ i_20_) ) | ( i_21_ ) | ( n536 ) ;
 assign n658 = ( i_2_  &  (~ n589) ) ;
 assign n659 = ( i_0_  &  (~ i_2_) ) | ( (~ i_2_)  &  i_3_ ) ;
 assign n661 = ( n407  &  n177 ) ;
 assign o_94_ = ( i_23_ ) ;


endmodule

