module C880 (
	_1gat_0_, _85gat_17_, _135gat_32_, _152gat_37_, _210gat_49_, _259gat_55_, _36gat_6_, _55gat_9_, 
	_75gat_15_, _159gat_40_, _237gat_52_, _138gat_33_, _8gat_1_, _219gat_50_, _26gat_4_, _74gat_14_, _153gat_38_, _59gat_10_, 
	_207gat_48_, _261gat_57_, _88gat_20_, _183gat_44_, _149gat_36_, _260gat_56_, _13gat_2_, _73gat_13_, _116gat_28_, _130gat_31_, 
	_246gat_53_, _89gat_21_, _111gat_27_, _189gat_45_, _68gat_11_, _72gat_12_, _268gat_59_, _90gat_22_, _143gat_34_, _201gat_47_, 
	_267gat_58_, _101gat_25_, _171gat_42_, _29gat_5_, _228gat_51_, _91gat_23_, _146gat_35_, _51gat_8_, _80gat_16_, _87gat_19_, 
	_165gat_41_, _255gat_54_, _156gat_39_, _177gat_43_, _42gat_7_, _86gat_18_, _17gat_3_, _96gat_24_, _106gat_26_, _121gat_29_, 
	_195gat_46_, _126gat_30_, _768gat_334_, _388gat_133_, _420gat_158_, _423gat_155_, _419gat_164_, _850gat_404_, _389gat_132_, _767gat_349_, 
	_874gat_433_, _418gat_168_, _421gat_162_, _422gat_161_, _878gat_442_, _450gat_173_, _447gat_182_, _879gat_441_, _449gat_176_, _863gat_424_, 
	_446gat_183_, _866gat_426_, _880gat_440_, _391gat_124_, _448gat_179_, _865gat_422_, _390gat_131_, _864gat_423_);

input _1gat_0_, _85gat_17_, _135gat_32_, _152gat_37_, _210gat_49_, _259gat_55_, _36gat_6_, _55gat_9_, _75gat_15_, _159gat_40_, _237gat_52_, _138gat_33_, _8gat_1_, _219gat_50_, _26gat_4_, _74gat_14_, _153gat_38_, _59gat_10_, _207gat_48_, _261gat_57_, _88gat_20_, _183gat_44_, _149gat_36_, _260gat_56_, _13gat_2_, _73gat_13_, _116gat_28_, _130gat_31_, _246gat_53_, _89gat_21_, _111gat_27_, _189gat_45_, _68gat_11_, _72gat_12_, _268gat_59_, _90gat_22_, _143gat_34_, _201gat_47_, _267gat_58_, _101gat_25_, _171gat_42_, _29gat_5_, _228gat_51_, _91gat_23_, _146gat_35_, _51gat_8_, _80gat_16_, _87gat_19_, _165gat_41_, _255gat_54_, _156gat_39_, _177gat_43_, _42gat_7_, _86gat_18_, _17gat_3_, _96gat_24_, _106gat_26_, _121gat_29_, _195gat_46_, _126gat_30_;

output _768gat_334_, _388gat_133_, _420gat_158_, _423gat_155_, _419gat_164_, _850gat_404_, _389gat_132_, _767gat_349_, _874gat_433_, _418gat_168_, _421gat_162_, _422gat_161_, _878gat_442_, _450gat_173_, _447gat_182_, _879gat_441_, _449gat_176_, _863gat_424_, _446gat_183_, _866gat_426_, _880gat_440_, _391gat_124_, _448gat_179_, _865gat_422_, _390gat_131_, _864gat_423_;

wire n_n678, n_n661, n_n646, n_n641, n_n629, n_n623, n_n672, n_n669, n_n663, n_n638, n_n626, n_n645, n_n677, n_n628, n_n674, n_n664, n_n640, n_n668, n_n630, n_n621, n_n658, n_n634, n_n642, n_n622, n_n676, n_n665, n_n650, n_n647, n_n625, n_n657, n_n651, n_n633, n_n667, n_n666, n_n619, n_n656, n_n644, n_n631, n_n620, n_n653, n_n636, n_n673, n_n627, n_n655, n_n643, n_n670, n_n662, n_n659, n_n637, n_n624, n_n639, n_n635, n_n671, n_n660, n_n675, n_n654, n_n652, n_n649, n_n632, n_n648, n_n266, n_n598, n_n587, n_n576, n_n245, n_n236, n_n523, n_n511, n_n499, n_n488, n_n215, n_n466, n_n209, n_n440, n_n198, n_n187, n_n405, n_n388, n_n377, n_n180, n_n174, n_n325, n_n313, n_n298, n_n282, n_n279, n_n287, n_n144, n_n127, n_n118, n_n107, n_n353, n_n363, n_n91, n_n399, n_n60, n_n450, n_n53, n_n45, n_n480, n_n496, n_n260, n_n597, n_n254, n_n575, n_n246, n_n234, n_n232, n_n510, n_n500, n_n487, n_n216, n_n476, n_n208, n_n441, n_n197, n_n188, n_n403, n_n389, n_n376, n_n181, n_n335, n_n326, n_n165, n_n162, n_n160, n_n278, n_n288, n_n145, n_n319, n_n117, n_n108, n_n354, n_n362, n_n90, n_n84, n_n431, n_n449, n_n52, n_n46, n_n481, n_n35, n_n268, n_n261, n_n574, n_n243, n_n237, n_n233, n_n509, n_n497, n_n490, n_n217, n_n207, n_n438, n_n200, n_n189, n_n401, n_n386, n_n379, n_n182, n_n334, n_n170, n_n315, n_n303, n_n159, n_n281, n_n152, n_n146, n_n131, n_n332, n_n109, n_n97, n_n365, n_n93, n_n85, n_n70, n_n65, n_n460, n_n43, n_n479, n_n36, n_n267, n_n601, n_n573, n_n244, n_n552, n_n529, n_n508, n_n498, n_n489, n_n218, n_n206, n_n439, n_n199, n_n190, n_n400, n_n387, n_n378, n_n183, n_n333, n_n171, n_n314, n_n304, n_n158, n_n280, n_n286, n_n147, n_n130, n_n126, n_n119, n_n96, n_n364, n_n92, n_n396, n_n421, n_n426, n_n461, n_n44, n_n39, n_n495, n_n594, n_n252, n_n557, n_n532, n_n473, n_n213, n_n191, n_n398, n_n177, n_n343, n_n272, n_n156, n_n302, n_n137, n_n356, n_n367, n_n88, n_n404, n_n414, n_n462, n_n468, n_n482, n_n31, n_n604, n_n593, n_n584, n_n238, n_n535, n_n472, n_n463, n_n201, n_n385, n_n176, n_n344, n_n273, n_n157, n_n143, n_n312, n_n357, n_n366, n_n402, n_n406, n_n74, n_n51, n_n42, n_n492, n_n32, n_n259, n_n585, n_n578, n_n247, n_n475, n_n464, n_n442, n_n375, n_n178, n_n345, n_n289, n_n300, n_n311, n_n358, n_n390, n_n82, n_n50, n_n41, n_n38, n_n33, n_n258, n_n253, n_n251, n_n248, n_n474, n_n465, n_n210, n_n179, n_n355, n_n346, n_n290, n_n299, n_n301, n_n368, n_n89, n_n83, n_n49, n_n477, n_n37, n_n34, n_n617, n_n606, n_n255, n_n579, n_n225, n_n485, n_n469, n_n458, n_n445, n_n374, n_n350, n_n339, n_n328, n_n316, n_n140, n_n133, n_n129, n_n120, n_n110, n_n80, n_n73, n_n424, n_n429, n_n446, n_n56, n_n610, n_n616, n_n264, n_n589, n_n580, n_n224, n_n486, n_n214, n_n459, n_n202, n_n384, n_n349, n_n340, n_n172, n_n166, n_n139, n_n134, n_n128, n_n121, n_n100, n_n79, n_n418, n_n67, n_n62, n_n448, n_n57, n_n609, n_n265, n_n257, n_n581, n_n230, n_n506, n_n471, n_n211, n_n192, n_n397, n_n175, n_n341, n_n306, n_n292, n_n142, n_n135, n_n327, n_n112, n_n101, n_n408, n_n416, n_n66, n_n61, n_n443, n_n456, n_n608, n_n256, n_n582, n_n516, n_n507, n_n470, n_n212, n_n413, n_n412, n_n351, n_n342, n_n305, n_n293, n_n141, n_n136, n_n336, n_n111, n_n102, n_n81, n_n415, n_n425, n_n430, n_n444, n_n455, n_n607, n_n270, n_n602, n_n572, n_n241, n_n541, n_n231, n_n229, n_n504, n_n221, n_n219, n_n205, n_n436, n_n194, n_n184, n_n411, n_n394, n_n381, n_n370, n_n173, n_n320, n_n308, n_n294, n_n291, n_n275, n_n284, n_n148, n_n310, n_n321, n_n124, n_n114, n_n103, n_n359, n_n95, n_n86, n_n76, n_n71, n_n422, n_n427, n_n58, n_n454, n_n40, n_n494, n_n614, n_n269, n_n262, n_n250, n_n242, n_n538, n_n520, n_n514, n_n505, n_n491, n_n220, n_n204, n_n437, n_n193, n_n185, n_n410, n_n395, n_n380, n_n371, n_n331, n_n169, n_n307, n_n295, n_n161, n_n274, n_n153, n_n149, n_n318, n_n322, n_n125, n_n113, n_n104, n_n99, n_n94, n_n87, n_n75, n_n420, n_n69, n_n64, n_n433, n_n453, n_n478, n_n493, n_n613, n_n615, n_n263, n_n249, n_n239, n_n547, n_n521, n_n228, n_n226, n_n223, n_n483, n_n467, n_n203, n_n434, n_n196, n_n186, n_n409, n_n391, n_n383, n_n372, n_n348, n_n337, n_n330, n_n167, n_n164, n_n296, n_n285, n_n277, n_n155, n_n150, n_n138, n_n317, n_n323, n_n122, n_n116, n_n105, n_n98, n_n361, n_n393, n_n78, n_n419, n_n68, n_n63, n_n432, n_n452, n_n55, n_n47, n_n612, n_n271, n_n605, n_n569, n_n240, n_n543, n_n522, n_n512, n_n227, n_n222, n_n484, n_n457, n_n447, n_n435, n_n195, n_n417, n_n407, n_n392, n_n382, n_n373, n_n347, n_n338, n_n329, n_n168, n_n163, n_n297, n_n283, n_n276, n_n154, n_n151, n_n309, n_n132, n_n324, n_n123, n_n115, n_n106, n_n352, n_n360, n_n369, n_n77, n_n72, n_n423, n_n428, n_n59, n_n451, n_n54, n_n48, n_n611, n_n28, n_n517, n_n531, n_n17, n_n12, n_n29, n_n518, n_n530, n_n16, n_n553, n_n503, n_n519, n_n534, n_n545, n_n13, n_n502, n_n19, n_n533, n_n546, n_n551, n_n618, n_n501, n_n561, n_n10, n_n592, n_n0, n_n30, n_n562, n_n11, n_n595, n_n1, n_n563, n_n583, n_n7, n_n603, n_n564, n_n577, n_n6, n_n600, n_n536, n_n235, n_n556, n_n568, n_n590, n_n2, n_n537, n_n548, n_n558, n_n567, n_n591, n_n3, n_n23, n_n524, n_n559, n_n571, n_n9, n_n599, n_n22, n_n18, n_n560, n_n570, n_n8, n_n596, n_n24, n_n21, n_n526, n_n542, n_n550, n_n586, n_n4, n_n25, n_n20, n_n525, n_n544, n_n549, n_n588, n_n5, n_n26, n_n513, n_n528, n_n539, n_n14, n_n554, n_n566, n_n27, n_n515, n_n527, n_n540, n_n15, n_n555, n_n565;

assign n_n678 = ( _1gat_0_ ) ;
 assign n_n661 = ( _85gat_17_ ) ;
 assign _768gat_334_ = ( n_n410 ) ;
 assign n_n646 = ( _135gat_32_ ) ;
 assign n_n641 = ( _152gat_37_ ) ;
 assign n_n629 = ( _210gat_49_ ) ;
 assign n_n623 = ( _259gat_55_ ) ;
 assign _388gat_133_ = ( n_n579 ) ;
 assign n_n672 = ( _36gat_6_ ) ;
 assign n_n669 = ( _55gat_9_ ) ;
 assign n_n663 = ( _75gat_15_ ) ;
 assign _420gat_158_ = ( n_n555 ) ;
 assign _423gat_155_ = ( n_n557 ) ;
 assign n_n638 = ( _159gat_40_ ) ;
 assign n_n626 = ( _237gat_52_ ) ;
 assign _419gat_164_ = ( n_n548 ) ;
 assign _850gat_404_ = ( n_n312 ) ;
 assign n_n645 = ( _138gat_33_ ) ;
 assign _389gat_132_ = ( n_n580 ) ;
 assign n_n677 = ( _8gat_1_ ) ;
 assign n_n628 = ( _219gat_50_ ) ;
 assign n_n674 = ( _26gat_4_ ) ;
 assign n_n664 = ( _74gat_14_ ) ;
 assign n_n640 = ( _153gat_38_ ) ;
 assign _767gat_349_ = ( n_n388 ) ;
 assign n_n668 = ( _59gat_10_ ) ;
 assign n_n630 = ( _207gat_48_ ) ;
 assign n_n621 = ( _261gat_57_ ) ;
 assign n_n658 = ( _88gat_20_ ) ;
 assign n_n634 = ( _183gat_44_ ) ;
 assign n_n642 = ( _149gat_36_ ) ;
 assign n_n622 = ( _260gat_56_ ) ;
 assign _874gat_433_ = ( n_n281 ) ;
 assign n_n676 = ( _13gat_2_ ) ;
 assign n_n665 = ( _73gat_13_ ) ;
 assign n_n650 = ( _116gat_28_ ) ;
 assign n_n647 = ( _130gat_31_ ) ;
 assign n_n625 = ( _246gat_53_ ) ;
 assign _418gat_168_ = ( n_n544 ) ;
 assign n_n657 = ( _89gat_21_ ) ;
 assign n_n651 = ( _111gat_27_ ) ;
 assign n_n633 = ( _189gat_45_ ) ;
 assign n_n667 = ( _68gat_11_ ) ;
 assign n_n666 = ( _72gat_12_ ) ;
 assign _421gat_162_ = ( n_n550 ) ;
 assign _422gat_161_ = ( n_n551 ) ;
 assign _878gat_442_ = ( n_n272 ) ;
 assign n_n619 = ( _268gat_59_ ) ;
 assign n_n656 = ( _90gat_22_ ) ;
 assign n_n644 = ( _143gat_34_ ) ;
 assign n_n631 = ( _201gat_47_ ) ;
 assign n_n620 = ( _267gat_58_ ) ;
 assign _450gat_173_ = ( n_n530 ) ;
 assign n_n653 = ( _101gat_25_ ) ;
 assign n_n636 = ( _171gat_42_ ) ;
 assign n_n673 = ( _29gat_5_ ) ;
 assign n_n627 = ( _228gat_51_ ) ;
 assign _447gat_182_ = ( n_n525 ) ;
 assign n_n655 = ( _91gat_23_ ) ;
 assign n_n643 = ( _146gat_35_ ) ;
 assign _879gat_441_ = ( n_n273 ) ;
 assign n_n670 = ( _51gat_8_ ) ;
 assign n_n662 = ( _80gat_16_ ) ;
 assign n_n659 = ( _87gat_19_ ) ;
 assign n_n637 = ( _165gat_41_ ) ;
 assign _449gat_176_ = ( n_n528 ) ;
 assign _863gat_424_ = ( n_n288 ) ;
 assign _446gat_183_ = ( n_n524 ) ;
 assign _866gat_426_ = ( n_n286 ) ;
 assign _880gat_440_ = ( n_n274 ) ;
 assign n_n624 = ( _255gat_54_ ) ;
 assign n_n639 = ( _156gat_39_ ) ;
 assign n_n635 = ( _177gat_43_ ) ;
 assign _391gat_124_ = ( n_n589 ) ;
 assign n_n671 = ( _42gat_7_ ) ;
 assign n_n660 = ( _86gat_18_ ) ;
 assign _448gat_179_ = ( n_n526 ) ;
 assign _865gat_422_ = ( n_n290 ) ;
 assign n_n675 = ( _17gat_3_ ) ;
 assign n_n654 = ( _96gat_24_ ) ;
 assign n_n652 = ( _106gat_26_ ) ;
 assign n_n649 = ( _121gat_29_ ) ;
 assign n_n632 = ( _195gat_46_ ) ;
 assign _390gat_131_ = ( n_n576 ) ;
 assign _864gat_423_ = ( n_n289 ) ;
 assign n_n648 = ( _126gat_30_ ) ;
 assign n_n266 = ( n_n635  &  n_n636 ) ;
 assign n_n598 = ( n_n652  &  n_n629 ) ;
 assign n_n587 = ( n_n663  &  n_n662  &  n_n668 ) ;
 assign n_n576 = ( n_n672  &  n_n671  &  n_n673 ) ;
 assign n_n245 = ( n_n612  &  n_n611 ) ;
 assign n_n236 = ( n_n14  &  n_n15 ) ;
 assign n_n523 = ( n_n542  &  n_n540 ) ;
 assign n_n511 = ( n_n22  &  n_n23 ) ;
 assign n_n499 = ( n_n30  &  n_n32 ) ;
 assign n_n488 = ( n_n637  &  n_n503 ) ;
 assign n_n215 = ( n_n504  &  n_n647 ) ;
 assign n_n466 = ( n_n44  &  n_n45 ) ;
 assign n_n209 = ( n_n465  &  n_n513 ) ;
 assign n_n440 = ( n_n455  &  n_n625 ) ;
 assign n_n198 = ( n_n62  &  n_n63 ) ;
 assign n_n187 = ( n_n638  &  n_n452 ) ;
 assign n_n405 = ( n_n428  &  n_n429 ) ;
 assign n_n388 = ( n_n92  &  n_n93 ) ;
 assign n_n377 = ( n_n409  &  n_n627 ) ;
 assign n_n180 = ( n_n399  &  n_n423 ) ;
 assign n_n174 = ( n_n354  &  n_n427 ) ;
 assign n_n325 = ( n_n332  &  n_n400 ) ;
 assign n_n313 = ( n_n320  &  n_n628 ) ;
 assign n_n298 = ( n_n144  &  n_n145 ) ;
 assign n_n282 = ( n_n156  &  n_n157 ) ;
 assign n_n279 = ( (~ n_n159) ) ;
 assign n_n287 = ( (~ n_n161) ) ;
 assign n_n144 = ( (~ n_n307) ) ;
 assign n_n127 = ( (~ n_n605) ) ;
 assign n_n118 = ( (~ n_n354) ) ;
 assign n_n107 = ( (~ n_n373) ) ;
 assign n_n353 = ( (~ n_n176) ) ;
 assign n_n363 = ( (~ n_n402) ) ;
 assign n_n91 = ( (~ n_n435) ) ;
 assign n_n399 = ( (~ n_n424) ) ;
 assign n_n60 = ( (~ n_n632) ) ;
 assign n_n450 = ( (~ n_n204) ) ;
 assign n_n53 = ( (~ n_n585) ) ;
 assign n_n45 = ( (~ n_n485) ) ;
 assign n_n480 = ( (~ n_n218) ) ;
 assign n_n496 = ( (~ n_n225) ) ;
 assign n_n260 = ( n_n650  &  n_n651 ) ;
 assign n_n597 = ( n_n653  &  n_n629 ) ;
 assign n_n254 = ( n_n639  &  n_n668 ) ;
 assign n_n575 = ( n_n671  &  n_n675 ) ;
 assign n_n246 = ( n_n614  &  n_n613 ) ;
 assign n_n234 = ( n_n235  &  n_n19 ) ;
 assign n_n232 = ( n_n18  &  n_n19 ) ;
 assign n_n510 = ( n_n24  &  n_n25 ) ;
 assign n_n500 = ( n_n30  &  n_n31 ) ;
 assign n_n487 = ( n_n638  &  n_n503 ) ;
 assign n_n216 = ( n_n40  &  n_n41 ) ;
 assign n_n476 = ( n_n502  &  n_n648 ) ;
 assign n_n208 = ( n_n466  &  n_n513 ) ;
 assign n_n441 = ( n_n454  &  n_n625 ) ;
 assign n_n197 = ( n_n633  &  n_n455 ) ;
 assign n_n188 = ( n_n72  &  n_n73 ) ;
 assign n_n403 = ( n_n426  &  n_n427 ) ;
 assign n_n389 = ( n_n90  &  n_n91 ) ;
 assign n_n376 = ( n_n407  &  n_n627 ) ;
 assign n_n181 = ( n_n406  &  n_n429 ) ;
 assign n_n335 = ( n_n120  &  n_n121 ) ;
 assign n_n326 = ( n_n128  &  n_n129 ) ;
 assign n_n165 = ( n_n493  &  n_n350  &  n_n412  &  n_n316 ) ;
 assign n_n162 = ( n_n419  &  n_n317 ) ;
 assign n_n160 = ( n_n346  &  n_n395  &  n_n283 ) ;
 assign n_n278 = ( (~ n_n158) ) ;
 assign n_n288 = ( (~ n_n299) ) ;
 assign n_n145 = ( (~ n_n308) ) ;
 assign n_n319 = ( (~ n_n168) ) ;
 assign n_n117 = ( (~ n_n405) ) ;
 assign n_n108 = ( (~ n_n380) ) ;
 assign n_n354 = ( (~ n_n177) ) ;
 assign n_n362 = ( (~ n_n399) ) ;
 assign n_n90 = ( (~ n_n487) ) ;
 assign n_n84 = ( (~ n_n490) ) ;
 assign n_n431 = ( (~ n_n200) ) ;
 assign n_n449 = ( (~ n_n203) ) ;
 assign n_n52 = ( (~ n_n470) ) ;
 assign n_n46 = ( (~ n_n474) ) ;
 assign n_n481 = ( (~ n_n219) ) ;
 assign n_n35 = ( (~ n_n630) ) ;
 assign n_n268 = ( n_n633  &  n_n634 ) ;
 assign n_n261 = ( n_n2  &  n_n3 ) ;
 assign n_n574 = ( n_n10  &  n_n11 ) ;
 assign n_n243 = ( n_n608  &  n_n607 ) ;
 assign n_n237 = ( n_n12  &  n_n15 ) ;
 assign n_n233 = ( n_n553  &  n_n546 ) ;
 assign n_n509 = ( n_n516  &  n_n640 ) ;
 assign n_n497 = ( n_n30  &  n_n34 ) ;
 assign n_n490 = ( n_n635  &  n_n503 ) ;
 assign n_n217 = ( n_n510  &  n_n647 ) ;
 assign n_n207 = ( n_n467  &  n_n513 ) ;
 assign n_n438 = ( n_n449  &  n_n625 ) ;
 assign n_n200 = ( n_n60  &  n_n61 ) ;
 assign n_n189 = ( n_n637  &  n_n451 ) ;
 assign n_n401 = ( n_n82  &  n_n83 ) ;
 assign n_n386 = ( n_n94  &  n_n95 ) ;
 assign n_n379 = ( n_n393  &  n_n626 ) ;
 assign n_n182 = ( n_n431  &  n_n408  &  n_n429 ) ;
 assign n_n334 = ( n_n122  &  n_n123 ) ;
 assign n_n170 = ( n_n425  &  n_n332  &  n_n423 ) ;
 assign n_n315 = ( n_n134  &  n_n135 ) ;
 assign n_n303 = ( n_n317  &  n_n391 ) ;
 assign n_n159 = ( n_n345  &  n_n392  &  n_n282 ) ;
 assign n_n281 = ( (~ n_n284) ) ;
 assign n_n152 = ( (~ n_n291) ) ;
 assign n_n146 = ( (~ n_n305) ) ;
 assign n_n131 = ( (~ n_n326) ) ;
 assign n_n332 = ( (~ n_n173) ) ;
 assign n_n109 = ( (~ n_n372) ) ;
 assign n_n97 = ( (~ n_n386) ) ;
 assign n_n365 = ( (~ n_n181) ) ;
 assign n_n93 = ( (~ n_n445) ) ;
 assign n_n85 = ( (~ n_n438) ) ;
 assign n_n70 = ( (~ n_n637) ) ;
 assign n_n65 = ( (~ n_n456) ) ;
 assign n_n460 = ( (~ n_n211) ) ;
 assign n_n43 = ( (~ n_n486) ) ;
 assign n_n479 = ( (~ n_n217) ) ;
 assign n_n36 = ( (~ n_n511) ) ;
 assign n_n267 = ( n_n66  &  n_n68 ) ;
 assign n_n601 = ( n_n651  &  n_n629 ) ;
 assign n_n573 = ( n_n645  &  n_n675 ) ;
 assign n_n244 = ( n_n610  &  n_n609 ) ;
 assign n_n552 = ( n_n13  &  n_n15 ) ;
 assign n_n529 = ( n_n665  &  n_n552 ) ;
 assign n_n508 = ( n_n516  &  n_n642 ) ;
 assign n_n498 = ( n_n30  &  n_n33 ) ;
 assign n_n489 = ( n_n636  &  n_n503 ) ;
 assign n_n218 = ( n_n39  &  n_n41 ) ;
 assign n_n206 = ( n_n500  &  n_n457 ) ;
 assign n_n439 = ( n_n456  &  n_n625 ) ;
 assign n_n199 = ( n_n632  &  n_n454 ) ;
 assign n_n190 = ( n_n70  &  n_n71 ) ;
 assign n_n400 = ( n_n424  &  n_n425 ) ;
 assign n_n387 = ( n_n621  &  n_n409 ) ;
 assign n_n378 = ( n_n390  &  n_n626 ) ;
 assign n_n183 = ( n_n408  &  n_n431 ) ;
 assign n_n333 = ( n_n124  &  n_n125 ) ;
 assign n_n171 = ( n_n332  &  n_n425 ) ;
 assign n_n314 = ( n_n136  &  n_n137 ) ;
 assign n_n304 = ( n_n142  &  n_n143 ) ;
 assign n_n158 = ( n_n344  &  n_n389  &  n_n285 ) ;
 assign n_n280 = ( (~ n_n160) ) ;
 assign n_n286 = ( (~ n_n295) ) ;
 assign n_n147 = ( (~ n_n306) ) ;
 assign n_n130 = ( (~ n_n325) ) ;
 assign n_n126 = ( (~ n_n343) ) ;
 assign n_n119 = ( (~ n_n403) ) ;
 assign n_n96 = ( (~ n_n387) ) ;
 assign n_n364 = ( (~ n_n404) ) ;
 assign n_n92 = ( (~ n_n417) ) ;
 assign n_n396 = ( (~ n_n422) ) ;
 assign n_n421 = ( (~ n_n190) ) ;
 assign n_n426 = ( (~ n_n195) ) ;
 assign n_n461 = ( (~ n_n212) ) ;
 assign n_n44 = ( (~ n_n475) ) ;
 assign n_n39 = ( (~ n_n510) ) ;
 assign n_n495 = ( (~ n_n224) ) ;
 assign n_n594 = ( n_n654  &  n_n629 ) ;
 assign n_n252 = ( n_n666  &  n_n671  &  n_n667  &  n_n668 ) ;
 assign n_n557 = ( n_n590  &  n_n656 ) ;
 assign n_n532 = ( n_n559  &  n_n558 ) ;
 assign n_n473 = ( n_n502  &  n_n651 ) ;
 assign n_n213 = ( n_n482  &  n_n481 ) ;
 assign n_n191 = ( n_n636  &  n_n450 ) ;
 assign n_n398 = ( n_n84  &  n_n85 ) ;
 assign n_n177 = ( n_n416  &  n_n365  &  n_n367  &  n_n364 ) ;
 assign n_n343 = ( n_n355  &  n_n628 ) ;
 assign n_n272 = ( (~ n_n275) ) ;
 assign n_n156 = ( (~ n_n292) ) ;
 assign n_n302 = ( (~ n_n162) ) ;
 assign n_n137 = ( (~ n_n598) ) ;
 assign n_n356 = ( (~ n_n390) ) ;
 assign n_n367 = ( (~ n_n182) ) ;
 assign n_n88 = ( (~ n_n488) ) ;
 assign n_n404 = ( (~ n_n428) ) ;
 assign n_n414 = ( (~ n_n184) ) ;
 assign n_n462 = ( (~ n_n213) ) ;
 assign n_n468 = ( (~ n_n214) ) ;
 assign n_n482 = ( (~ n_n220) ) ;
 assign n_n31 = ( (~ n_n506) ) ;
 assign n_n604 = ( (~ n_n263) ) ;
 assign n_n593 = ( n_n655  &  n_n629 ) ;
 assign n_n584 = ( n_n663  &  n_n671  &  n_n668 ) ;
 assign n_n238 = ( n_n590  &  n_n657 ) ;
 assign n_n535 = ( n_n561  &  n_n560 ) ;
 assign n_n472 = ( n_n502  &  n_n652 ) ;
 assign n_n463 = ( n_n50  &  n_n51 ) ;
 assign n_n201 = ( n_n631  &  n_n453 ) ;
 assign n_n385 = ( n_n408  &  n_n626 ) ;
 assign n_n176 = ( n_n368  &  n_n415  &  n_n366 ) ;
 assign n_n344 = ( n_n112  &  n_n113 ) ;
 assign n_n273 = ( (~ n_n276) ) ;
 assign n_n157 = ( (~ n_n593) ) ;
 assign n_n143 = ( (~ n_n391) ) ;
 assign n_n312 = ( (~ n_n321) ) ;
 assign n_n357 = ( (~ n_n393) ) ;
 assign n_n366 = ( (~ n_n406) ) ;
 assign n_n402 = ( (~ n_n426) ) ;
 assign n_n406 = ( (~ n_n430) ) ;
 assign n_n74 = ( (~ n_n442) ) ;
 assign n_n51 = ( (~ n_n606) ) ;
 assign n_n42 = ( (~ n_n476) ) ;
 assign n_n492 = ( (~ n_n221) ) ;
 assign n_n32 = ( (~ n_n507) ) ;
 assign n_n259 = ( n_n4  &  n_n5 ) ;
 assign n_n585 = ( n_n645  &  n_n670 ) ;
 assign n_n578 = ( n_n663  &  n_n662  &  n_n673 ) ;
 assign n_n247 = ( n_n675  &  n_n677  &  n_n676  &  n_n678 ) ;
 assign n_n475 = ( n_n502  &  n_n649 ) ;
 assign n_n464 = ( n_n48  &  n_n49 ) ;
 assign n_n442 = ( n_n453  &  n_n625 ) ;
 assign n_n375 = ( n_n405  &  n_n627 ) ;
 assign n_n178 = ( n_n396  &  n_n421 ) ;
 assign n_n345 = ( n_n110  &  n_n111 ) ;
 assign n_n289 = ( (~ n_n300) ) ;
 assign n_n300 = ( (~ n_n310) ) ;
 assign n_n311 = ( (~ n_n165) ) ;
 assign n_n358 = ( (~ n_n178) ) ;
 assign n_n390 = ( (~ n_n418) ) ;
 assign n_n82 = ( (~ n_n491) ) ;
 assign n_n50 = ( (~ n_n472) ) ;
 assign n_n41 = ( (~ n_n647) ) ;
 assign n_n38 = ( (~ n_n505) ) ;
 assign n_n33 = ( (~ n_n508) ) ;
 assign n_n258 = ( n_n652  &  n_n653 ) ;
 assign n_n253 = ( n_n667  &  n_n664  &  n_n668 ) ;
 assign n_n251 = ( n_n667  &  n_n673 ) ;
 assign n_n248 = ( n_n675  &  n_n674  &  n_n676  &  n_n678 ) ;
 assign n_n474 = ( n_n502  &  n_n650 ) ;
 assign n_n465 = ( n_n46  &  n_n47 ) ;
 assign n_n210 = ( n_n464  &  n_n513 ) ;
 assign n_n179 = ( n_n423  &  n_n399  &  n_n421 ) ;
 assign n_n355 = ( n_n96  &  n_n97 ) ;
 assign n_n346 = ( n_n108  &  n_n109 ) ;
 assign n_n290 = ( (~ n_n301) ) ;
 assign n_n299 = ( (~ n_n309) ) ;
 assign n_n301 = ( (~ n_n311) ) ;
 assign n_n368 = ( (~ n_n183) ) ;
 assign n_n89 = ( (~ n_n436) ) ;
 assign n_n83 = ( (~ n_n439) ) ;
 assign n_n49 = ( (~ n_n483) ) ;
 assign n_n477 = ( (~ n_n215) ) ;
 assign n_n37 = ( (~ n_n646) ) ;
 assign n_n34 = ( (~ n_n509) ) ;
 assign n_n617 = ( n_n620  &  n_n624 ) ;
 assign n_n606 = ( n_n645  &  n_n641 ) ;
 assign n_n255 = ( n_n8  &  n_n9 ) ;
 assign n_n579 = ( n_n663  &  n_n671  &  n_n673 ) ;
 assign n_n225 = ( n_n35  &  n_n36 ) ;
 assign n_n485 = ( n_n501  &  n_n642 ) ;
 assign n_n469 = ( n_n502  &  n_n655 ) ;
 assign n_n458 = ( n_n54  &  n_n55 ) ;
 assign n_n445 = ( n_n462  &  n_n460 ) ;
 assign n_n374 = ( n_n403  &  n_n627 ) ;
 assign n_n350 = ( n_n100  &  n_n101 ) ;
 assign n_n339 = ( n_n353  &  n_n405 ) ;
 assign n_n328 = ( n_n333  &  n_n628 ) ;
 assign n_n316 = ( n_n132  &  n_n133 ) ;
 assign n_n140 = ( (~ n_n318) ) ;
 assign n_n133 = ( (~ n_n602) ) ;
 assign n_n129 = ( (~ n_n400) ) ;
 assign n_n120 = ( (~ n_n341) ) ;
 assign n_n110 = ( (~ n_n379) ) ;
 assign n_n80 = ( (~ n_n434) ) ;
 assign n_n73 = ( (~ n_n452) ) ;
 assign n_n424 = ( (~ n_n193) ) ;
 assign n_n429 = ( (~ n_n198) ) ;
 assign n_n446 = ( (~ n_n462) ) ;
 assign n_n56 = ( (~ n_n469) ) ;
 assign n_n610 = ( (~ n_n267) ) ;
 assign n_n616 = ( n_n622  &  n_n624 ) ;
 assign n_n264 = ( n_n637  &  n_n638 ) ;
 assign n_n589 = ( n_n660  &  n_n661 ) ;
 assign n_n580 = ( n_n672  &  n_n662  &  n_n673 ) ;
 assign n_n224 = ( n_n630  &  n_n511 ) ;
 assign n_n486 = ( n_n501  &  n_n640 ) ;
 assign n_n214 = ( n_n496  &  n_n495 ) ;
 assign n_n459 = ( n_n52  &  n_n53 ) ;
 assign n_n202 = ( n_n58  &  n_n59 ) ;
 assign n_n384 = ( n_n406  &  n_n626 ) ;
 assign n_n349 = ( n_n102  &  n_n103 ) ;
 assign n_n340 = ( n_n116  &  n_n117 ) ;
 assign n_n172 = ( n_n494  &  n_n351  &  n_n413  &  n_n331 ) ;
 assign n_n166 = ( n_n322  &  n_n358  &  n_n360  &  n_n357 ) ;
 assign n_n139 = ( (~ n_n397) ) ;
 assign n_n134 = ( (~ n_n329) ) ;
 assign n_n128 = ( (~ n_n332) ) ;
 assign n_n121 = ( (~ n_n342) ) ;
 assign n_n100 = ( (~ n_n384) ) ;
 assign n_n79 = ( (~ n_n615) ) ;
 assign n_n418 = ( (~ n_n187) ) ;
 assign n_n67 = ( (~ n_n449) ) ;
 assign n_n62 = ( (~ n_n633) ) ;
 assign n_n448 = ( (~ n_n468) ) ;
 assign n_n57 = ( (~ n_n572) ) ;
 assign n_n609 = ( (~ n_n266) ) ;
 assign n_n265 = ( n_n70  &  n_n72 ) ;
 assign n_n257 = ( n_n6  &  n_n7 ) ;
 assign n_n581 = ( n_n672  &  n_n662  &  n_n668 ) ;
 assign n_n230 = ( n_n578  &  n_n669  &  n_n525 ) ;
 assign n_n506 = ( n_n516  &  n_n644 ) ;
 assign n_n471 = ( n_n502  &  n_n653 ) ;
 assign n_n211 = ( n_n478  &  n_n477 ) ;
 assign n_n192 = ( n_n68  &  n_n69 ) ;
 assign n_n397 = ( n_n422  &  n_n423 ) ;
 assign n_n175 = ( n_n414  &  n_n369 ) ;
 assign n_n341 = ( n_n352  &  n_n407 ) ;
 assign n_n306 = ( n_n140  &  n_n141 ) ;
 assign n_n292 = ( n_n297  &  n_n628 ) ;
 assign n_n142 = ( (~ n_n317) ) ;
 assign n_n135 = ( (~ n_n601) ) ;
 assign n_n327 = ( (~ n_n172) ) ;
 assign n_n112 = ( (~ n_n378) ) ;
 assign n_n101 = ( (~ n_n376) ) ;
 assign n_n408 = ( (~ n_n432) ) ;
 assign n_n416 = ( (~ n_n186) ) ;
 assign n_n66 = ( (~ n_n635) ) ;
 assign n_n61 = ( (~ n_n454) ) ;
 assign n_n443 = ( (~ n_n460) ) ;
 assign n_n456 = ( (~ n_n210) ) ;
 assign n_n608 = ( (~ n_n265) ) ;
 assign n_n256 = ( n_n654  &  n_n655 ) ;
 assign n_n582 = ( n_n672  &  n_n671  &  n_n668 ) ;
 assign n_n516 = ( n_n525  &  n_n669  &  n_n588 ) ;
 assign n_n507 = ( n_n516  &  n_n643 ) ;
 assign n_n470 = ( n_n502  &  n_n654 ) ;
 assign n_n212 = ( n_n480  &  n_n479 ) ;
 assign n_n413 = ( n_n74  &  n_n75 ) ;
 assign n_n412 = ( n_n76  &  n_n77 ) ;
 assign n_n351 = ( n_n98  &  n_n99 ) ;
 assign n_n342 = ( n_n114  &  n_n115 ) ;
 assign n_n305 = ( n_n318  &  n_n394 ) ;
 assign n_n293 = ( n_n298  &  n_n628 ) ;
 assign n_n141 = ( (~ n_n394) ) ;
 assign n_n136 = ( (~ n_n328) ) ;
 assign n_n336 = ( (~ n_n174) ) ;
 assign n_n111 = ( (~ n_n371) ) ;
 assign n_n102 = ( (~ n_n383) ) ;
 assign n_n81 = ( (~ n_n447) ) ;
 assign n_n415 = ( (~ n_n185) ) ;
 assign n_n425 = ( (~ n_n194) ) ;
 assign n_n430 = ( (~ n_n199) ) ;
 assign n_n444 = ( (~ n_n461) ) ;
 assign n_n455 = ( (~ n_n209) ) ;
 assign n_n607 = ( (~ n_n264) ) ;
 assign n_n270 = ( n_n631  &  n_n632 ) ;
 assign n_n602 = ( n_n650  &  n_n629 ) ;
 assign n_n572 = ( n_n645  &  n_n677 ) ;
 assign n_n241 = ( n_n600  &  n_n599 ) ;
 assign n_n541 = ( n_n565  &  n_n564 ) ;
 assign n_n231 = ( n_n525  &  n_n668  &  n_n639  &  n_n547 ) ;
 assign n_n229 = ( n_n588  &  n_n675  &  n_n525 ) ;
 assign n_n504 = ( n_n28  &  n_n29 ) ;
 assign n_n221 = ( n_n633  &  n_n503 ) ;
 assign n_n219 = ( n_n646  &  n_n505 ) ;
 assign n_n205 = ( n_n499  &  n_n459 ) ;
 assign n_n436 = ( n_n451  &  n_n625 ) ;
 assign n_n194 = ( n_n66  &  n_n67 ) ;
 assign n_n184 = ( n_n621  &  n_n433 ) ;
 assign n_n411 = ( n_n78  &  n_n79 ) ;
 assign n_n394 = ( n_n420  &  n_n421 ) ;
 assign n_n381 = ( n_n399  &  n_n626 ) ;
 assign n_n370 = ( n_n391  &  n_n627 ) ;
 assign n_n173 = ( n_n363  &  n_n336 ) ;
 assign n_n320 = ( n_n130  &  n_n131 ) ;
 assign n_n308 = ( n_n138  &  n_n139 ) ;
 assign n_n294 = ( n_n150  &  n_n151 ) ;
 assign n_n291 = ( n_n296  &  n_n628 ) ;
 assign n_n275 = ( (~ n_n278) ) ;
 assign n_n284 = ( (~ n_n287) ) ;
 assign n_n148 = ( (~ n_n303) ) ;
 assign n_n310 = ( (~ n_n164) ) ;
 assign n_n321 = ( (~ n_n327) ) ;
 assign n_n124 = ( (~ n_n337) ) ;
 assign n_n114 = ( (~ n_n352) ) ;
 assign n_n103 = ( (~ n_n375) ) ;
 assign n_n359 = ( (~ n_n396) ) ;
 assign n_n95 = ( (~ n_n409) ) ;
 assign n_n86 = ( (~ n_n489) ) ;
 assign n_n76 = ( (~ n_n441) ) ;
 assign n_n71 = ( (~ n_n451) ) ;
 assign n_n422 = ( (~ n_n191) ) ;
 assign n_n427 = ( (~ n_n196) ) ;
 assign n_n58 = ( (~ n_n631) ) ;
 assign n_n454 = ( (~ n_n208) ) ;
 assign n_n40 = ( (~ n_n504) ) ;
 assign n_n494 = ( (~ n_n223) ) ;
 assign n_n614 = ( (~ n_n271) ) ;
 assign n_n269 = ( n_n62  &  n_n64 ) ;
 assign n_n262 = ( n_n648  &  n_n649 ) ;
 assign n_n250 = ( n_n669  &  n_n677  &  n_n676  &  n_n678 ) ;
 assign n_n242 = ( n_n604  &  n_n603 ) ;
 assign n_n538 = ( n_n563  &  n_n562 ) ;
 assign n_n520 = ( n_n533  &  n_n531 ) ;
 assign n_n514 = ( n_n675  &  n_n578  &  n_n525 ) ;
 assign n_n505 = ( n_n26  &  n_n27 ) ;
 assign n_n491 = ( n_n634  &  n_n503 ) ;
 assign n_n220 = ( n_n37  &  n_n38 ) ;
 assign n_n204 = ( n_n498  &  n_n458 ) ;
 assign n_n437 = ( n_n450  &  n_n625 ) ;
 assign n_n193 = ( n_n635  &  n_n449 ) ;
 assign n_n185 = ( n_n433  &  n_n621  &  n_n431 ) ;
 assign n_n410 = ( n_n80  &  n_n81 ) ;
 assign n_n395 = ( n_n86  &  n_n87 ) ;
 assign n_n380 = ( n_n396  &  n_n626 ) ;
 assign n_n371 = ( n_n394  &  n_n627 ) ;
 assign n_n331 = ( n_n126  &  n_n127 ) ;
 assign n_n169 = ( n_n332  &  n_n423  &  n_n425  &  n_n421 ) ;
 assign n_n307 = ( n_n319  &  n_n397 ) ;
 assign n_n295 = ( n_n302  &  n_n356 ) ;
 assign n_n161 = ( n_n347  &  n_n398  &  n_n294 ) ;
 assign n_n274 = ( (~ n_n277) ) ;
 assign n_n153 = ( (~ n_n543) ) ;
 assign n_n149 = ( (~ n_n304) ) ;
 assign n_n318 = ( (~ n_n167) ) ;
 assign n_n322 = ( (~ n_n169) ) ;
 assign n_n125 = ( (~ n_n338) ) ;
 assign n_n113 = ( (~ n_n370) ) ;
 assign n_n104 = ( (~ n_n382) ) ;
 assign n_n99 = ( (~ n_n377) ) ;
 assign n_n94 = ( (~ n_n621) ) ;
 assign n_n87 = ( (~ n_n437) ) ;
 assign n_n75 = ( (~ n_n617) ) ;
 assign n_n420 = ( (~ n_n189) ) ;
 assign n_n69 = ( (~ n_n450) ) ;
 assign n_n64 = ( (~ n_n634) ) ;
 assign n_n433 = ( (~ n_n202) ) ;
 assign n_n453 = ( (~ n_n207) ) ;
 assign n_n478 = ( (~ n_n216) ) ;
 assign n_n493 = ( (~ n_n222) ) ;
 assign n_n613 = ( (~ n_n270) ) ;
 assign n_n615 = ( n_n623  &  n_n624 ) ;
 assign n_n263 = ( n_n0  &  n_n1 ) ;
 assign n_n249 = ( n_n675  &  n_n677  &  n_n670  &  n_n678 ) ;
 assign n_n239 = ( n_n592  &  n_n591 ) ;
 assign n_n547 = ( n_n16  &  n_n17 ) ;
 assign n_n521 = ( n_n536  &  n_n534 ) ;
 assign n_n228 = ( n_n20  &  n_n21 ) ;
 assign n_n226 = ( n_n678  &  n_n515 ) ;
 assign n_n223 = ( n_n631  &  n_n503 ) ;
 assign n_n483 = ( n_n501  &  n_n644 ) ;
 assign n_n467 = ( n_n42  &  n_n43 ) ;
 assign n_n203 = ( n_n497  &  n_n463 ) ;
 assign n_n434 = ( n_n448  &  n_n444 ) ;
 assign n_n196 = ( n_n64  &  n_n65 ) ;
 assign n_n186 = ( n_n621  &  n_n431  &  n_n433  &  n_n429 ) ;
 assign n_n409 = ( n_n432  &  n_n433 ) ;
 assign n_n391 = ( n_n418  &  n_n419 ) ;
 assign n_n383 = ( n_n404  &  n_n626 ) ;
 assign n_n372 = ( n_n397  &  n_n627 ) ;
 assign n_n348 = ( n_n104  &  n_n105 ) ;
 assign n_n337 = ( n_n354  &  n_n403 ) ;
 assign n_n330 = ( n_n335  &  n_n628 ) ;
 assign n_n167 = ( n_n361  &  n_n323  &  n_n359 ) ;
 assign n_n164 = ( n_n492  &  n_n349  &  n_n411  &  n_n315 ) ;
 assign n_n296 = ( n_n148  &  n_n149 ) ;
 assign n_n285 = ( n_n152  &  n_n153 ) ;
 assign n_n277 = ( (~ n_n280) ) ;
 assign n_n155 = ( (~ n_n594) ) ;
 assign n_n150 = ( (~ n_n313) ) ;
 assign n_n138 = ( (~ n_n319) ) ;
 assign n_n317 = ( (~ n_n166) ) ;
 assign n_n323 = ( (~ n_n170) ) ;
 assign n_n122 = ( (~ n_n339) ) ;
 assign n_n116 = ( (~ n_n353) ) ;
 assign n_n105 = ( (~ n_n374) ) ;
 assign n_n98 = ( (~ n_n385) ) ;
 assign n_n361 = ( (~ n_n180) ) ;
 assign n_n393 = ( (~ n_n420) ) ;
 assign n_n78 = ( (~ n_n440) ) ;
 assign n_n419 = ( (~ n_n188) ) ;
 assign n_n68 = ( (~ n_n636) ) ;
 assign n_n63 = ( (~ n_n455) ) ;
 assign n_n432 = ( (~ n_n201) ) ;
 assign n_n452 = ( (~ n_n206) ) ;
 assign n_n55 = ( (~ n_n573) ) ;
 assign n_n47 = ( (~ n_n484) ) ;
 assign n_n612 = ( (~ n_n269) ) ;
 assign n_n271 = ( n_n58  &  n_n60 ) ;
 assign n_n605 = ( n_n649  &  n_n629 ) ;
 assign n_n569 = ( n_n674  &  n_n670  &  n_n678 ) ;
 assign n_n240 = ( n_n596  &  n_n595 ) ;
 assign n_n543 = ( n_n566  &  n_n629 ) ;
 assign n_n522 = ( n_n539  &  n_n537 ) ;
 assign n_n512 = ( n_n514  &  n_n618 ) ;
 assign n_n227 = ( n_n527  &  n_n518 ) ;
 assign n_n222 = ( n_n632  &  n_n503 ) ;
 assign n_n484 = ( n_n501  &  n_n643 ) ;
 assign n_n457 = ( n_n56  &  n_n57 ) ;
 assign n_n447 = ( n_n468  &  n_n461 ) ;
 assign n_n435 = ( n_n452  &  n_n625 ) ;
 assign n_n195 = ( n_n634  &  n_n456 ) ;
 assign n_n417 = ( n_n446  &  n_n443 ) ;
 assign n_n407 = ( n_n430  &  n_n431 ) ;
 assign n_n392 = ( n_n88  &  n_n89 ) ;
 assign n_n382 = ( n_n402  &  n_n626 ) ;
 assign n_n373 = ( n_n400  &  n_n627 ) ;
 assign n_n347 = ( n_n106  &  n_n107 ) ;
 assign n_n338 = ( n_n118  &  n_n119 ) ;
 assign n_n329 = ( n_n334  &  n_n628 ) ;
 assign n_n168 = ( n_n324  &  n_n362 ) ;
 assign n_n163 = ( n_n348  &  n_n401  &  n_n314 ) ;
 assign n_n297 = ( n_n146  &  n_n147 ) ;
 assign n_n283 = ( n_n154  &  n_n155 ) ;
 assign n_n276 = ( (~ n_n279) ) ;
 assign n_n154 = ( (~ n_n293) ) ;
 assign n_n151 = ( (~ n_n597) ) ;
 assign n_n309 = ( (~ n_n163) ) ;
 assign n_n132 = ( (~ n_n330) ) ;
 assign n_n324 = ( (~ n_n171) ) ;
 assign n_n123 = ( (~ n_n340) ) ;
 assign n_n115 = ( (~ n_n407) ) ;
 assign n_n106 = ( (~ n_n381) ) ;
 assign n_n352 = ( (~ n_n175) ) ;
 assign n_n360 = ( (~ n_n179) ) ;
 assign n_n369 = ( (~ n_n408) ) ;
 assign n_n77 = ( (~ n_n616) ) ;
 assign n_n72 = ( (~ n_n638) ) ;
 assign n_n423 = ( (~ n_n192) ) ;
 assign n_n428 = ( (~ n_n197) ) ;
 assign n_n59 = ( (~ n_n453) ) ;
 assign n_n451 = ( (~ n_n205) ) ;
 assign n_n54 = ( (~ n_n471) ) ;
 assign n_n48 = ( (~ n_n473) ) ;
 assign n_n611 = ( (~ n_n268) ) ;
 assign n_n28 = ( (~ n_n520) ) ;
 assign n_n517 = ( (~ n_n230) ) ;
 assign n_n531 = ( (~ n_n558) ) ;
 assign n_n17 = ( (~ n_n574) ) ;
 assign n_n12 = ( (~ n_n586) ) ;
 assign n_n29 = ( (~ n_n532) ) ;
 assign n_n518 = ( (~ n_n231) ) ;
 assign n_n530 = ( (~ n_n556) ) ;
 assign n_n16 = ( (~ n_n575) ) ;
 assign n_n553 = ( (~ n_n584) ) ;
 assign n_n503 = ( (~ n_n519) ) ;
 assign n_n519 = ( (~ n_n529) ) ;
 assign n_n534 = ( (~ n_n560) ) ;
 assign n_n545 = ( (~ n_n569) ) ;
 assign n_n13 = ( (~ n_n583) ) ;
 assign n_n502 = ( (~ n_n227) ) ;
 assign n_n19 = ( (~ n_n568) ) ;
 assign n_n533 = ( (~ n_n559) ) ;
 assign n_n546 = ( (~ n_n570) ) ;
 assign n_n551 = ( (~ n_n582) ) ;
 assign n_n618 = ( (~ n_n619) ) ;
 assign n_n501 = ( (~ n_n226) ) ;
 assign n_n561 = ( (~ n_n242) ) ;
 assign n_n10 = ( (~ n_n671) ) ;
 assign n_n592 = ( (~ n_n257) ) ;
 assign n_n0 = ( (~ n_n648) ) ;
 assign n_n30 = ( (~ n_n512) ) ;
 assign n_n562 = ( (~ n_n243) ) ;
 assign n_n11 = ( (~ n_n675) ) ;
 assign n_n595 = ( (~ n_n258) ) ;
 assign n_n1 = ( (~ n_n649) ) ;
 assign n_n563 = ( (~ n_n244) ) ;
 assign n_n583 = ( (~ n_n252) ) ;
 assign n_n7 = ( (~ n_n655) ) ;
 assign n_n603 = ( (~ n_n262) ) ;
 assign n_n564 = ( (~ n_n245) ) ;
 assign n_n577 = ( (~ n_n251) ) ;
 assign n_n6 = ( (~ n_n654) ) ;
 assign n_n600 = ( (~ n_n261) ) ;
 assign n_n536 = ( (~ n_n561) ) ;
 assign n_n235 = ( (~ n_n576) ) ;
 assign n_n556 = ( (~ n_n238) ) ;
 assign n_n568 = ( (~ n_n248) ) ;
 assign n_n590 = ( (~ n_n255) ) ;
 assign n_n2 = ( (~ n_n650) ) ;
 assign n_n537 = ( (~ n_n562) ) ;
 assign n_n548 = ( (~ n_n234) ) ;
 assign n_n558 = ( (~ n_n239) ) ;
 assign n_n567 = ( (~ n_n247) ) ;
 assign n_n591 = ( (~ n_n256) ) ;
 assign n_n3 = ( (~ n_n651) ) ;
 assign n_n23 = ( (~ n_n541) ) ;
 assign n_n524 = ( (~ n_n232) ) ;
 assign n_n559 = ( (~ n_n240) ) ;
 assign n_n571 = ( (~ n_n250) ) ;
 assign n_n9 = ( (~ n_n659) ) ;
 assign n_n599 = ( (~ n_n260) ) ;
 assign n_n22 = ( (~ n_n523) ) ;
 assign n_n18 = ( (~ n_n235) ) ;
 assign n_n560 = ( (~ n_n241) ) ;
 assign n_n570 = ( (~ n_n249) ) ;
 assign n_n8 = ( (~ n_n658) ) ;
 assign n_n596 = ( (~ n_n259) ) ;
 assign n_n24 = ( (~ n_n522) ) ;
 assign n_n21 = ( (~ n_n566) ) ;
 assign n_n526 = ( (~ n_n549) ) ;
 assign n_n542 = ( (~ n_n565) ) ;
 assign n_n550 = ( (~ n_n581) ) ;
 assign n_n586 = ( (~ n_n253) ) ;
 assign n_n4 = ( (~ n_n652) ) ;
 assign n_n25 = ( (~ n_n538) ) ;
 assign n_n20 = ( (~ n_n517) ) ;
 assign n_n525 = ( (~ n_n545) ) ;
 assign n_n544 = ( (~ n_n567) ) ;
 assign n_n549 = ( (~ n_n236) ) ;
 assign n_n588 = ( (~ n_n254) ) ;
 assign n_n5 = ( (~ n_n653) ) ;
 assign n_n26 = ( (~ n_n521) ) ;
 assign n_n513 = ( (~ n_n228) ) ;
 assign n_n528 = ( (~ n_n554) ) ;
 assign n_n539 = ( (~ n_n563) ) ;
 assign n_n14 = ( (~ n_n577) ) ;
 assign n_n554 = ( (~ n_n237) ) ;
 assign n_n566 = ( (~ n_n618) ) ;
 assign n_n27 = ( (~ n_n535) ) ;
 assign n_n515 = ( (~ n_n229) ) ;
 assign n_n527 = ( (~ n_n233) ) ;
 assign n_n540 = ( (~ n_n564) ) ;
 assign n_n15 = ( (~ n_n571) ) ;
 assign n_n555 = ( (~ n_n587) ) ;
 assign n_n565 = ( (~ n_n246) ) ;


endmodule

