module ex5p_mapped (
	i_7_, i_5_, i_6_, i_3_, i_4_, i_1_, i_2_, i_0_, 
	o_1_, o_19_, o_2_, o_0_, o_29_, o_60_, o_39_, o_38_, o_25_, o_12_, 
	o_37_, o_26_, o_11_, o_50_, o_36_, o_27_, o_14_, o_35_, o_28_, o_13_, 
	o_34_, o_21_, o_16_, o_40_, o_33_, o_22_, o_15_, o_32_, o_23_, o_18_, 
	o_31_, o_24_, o_17_, o_56_, o_43_, o_30_, o_55_, o_44_, o_58_, o_41_, 
	o_57_, o_42_, o_20_, o_52_, o_47_, o_51_, o_48_, o_54_, o_45_, o_10_, 
	o_53_, o_46_, o_61_, o_9_, o_62_, o_49_, o_7_, o_8_, o_5_, o_59_, 
	o_6_, o_3_, o_4_);

input i_7_, i_5_, i_6_, i_3_, i_4_, i_1_, i_2_, i_0_;

output o_1_, o_19_, o_2_, o_0_, o_29_, o_60_, o_39_, o_38_, o_25_, o_12_, o_37_, o_26_, o_11_, o_50_, o_36_, o_27_, o_14_, o_35_, o_28_, o_13_, o_34_, o_21_, o_16_, o_40_, o_33_, o_22_, o_15_, o_32_, o_23_, o_18_, o_31_, o_24_, o_17_, o_56_, o_43_, o_30_, o_55_, o_44_, o_58_, o_41_, o_57_, o_42_, o_20_, o_52_, o_47_, o_51_, o_48_, o_54_, o_45_, o_10_, o_53_, o_46_, o_61_, o_9_, o_62_, o_49_, o_7_, o_8_, o_5_, o_59_, o_6_, o_3_, o_4_;

wire wire3179, wire3180, wire3184, n_n744, wire248, n_n0, wire71, wire3188, wire3189, wire3190, wire3191, wire3204, wire3205, wire3209, n_n7, wire3266, wire3267, wire3268, wire3269, n_n136, wire3332, wire3333, wire3334, wire3377, wire3378, wire3381, n_n2, n_n5, n_n8, wire3417, wire3418, wire3424, wire3428, n_n17, n_n19, n_n6, wire3452, wire3453, wire3454, wire3455, wire3481, wire3482, n_n3, n_n4, n_n12, wire3502, wire3503, n_n11, wire3526, wire3527, wire3528, wire3566, wire3567, wire3568, wire3569, wire3598, wire3599, wire3600, wire3601, wire3614, wire3615, wire3618, n_n1017, wire3619, n_n13, n_n1, wire318, wire3605, wire180, wire3636, wire322, wire3639, wire3660, wire3663, n_n371, wire3705, wire3706, wire3710, wire3733, wire3743, wire3744, wire3745, wire3763, wire3764, wire321, wire3790, wire3795, wire3829, wire3830, wire3831, wire3832, wire314, wire3882, wire3908, wire3909, wire3910, wire3911, wire3921, wire3925, wire3966, wire3967, wire3968, wire3969, n_n476, wire263, wire264, wire4013, wire4014, wire4015, wire4016, wire3355, wire4031, wire4055, wire4056, wire4057, wire4058, wire4069, wire3344, wire3345, wire4093, wire4097, wire267, wire347, wire4108, wire4112, wire4117, wire4126, wire4127, wire4128, wire4129, wire4160, wire4161, wire4162, wire4163, wire4166, wire4167, wire4168, wire4169, n_n1154, n_n1245, n_n1215, n_n1274, n_n1305, n_n10, n_n9, n_n1121, n_n1180, n_n1211, n_n1271, n_n1302, wire246, wire354, n_n1168, n_n1321, n_n1169, wire73, wire92, wire93, wire94, wire146, wire147, wire186, wire208, wire249, n_n1120, n_n1083, wire236, wire3213, n_n1008, wire163, n_n1009, n_n18, n_n872, n_n958, n_n949, n_n1137, n_n14, wire108, wire85, n_n1021, n_n1020, wire115, n_n15, n_n1136, wire152, n_n864, wire69, wire187, n_n602, n_n1022, n_n1298, wire3218, wire192, wire222, n_n930, wire72, wire226, wire104, n_n1226, wire77, wire228, wire70, wire3221, wire3222, wire240, n_n1197, wire88, n_n955, wire3225, wire252, n_n950, n_n1208, wire551, wire280, wire254, wire269, wire301, wire194, n_n859, wire324, wire134, wire327, n_n387, wire3237, wire3238, wire330, wire300, wire127, wire331, n_n1133, wire3239, wire346, n_n1193, n_n1225, n_n936, n_n1194, wire285, wire3288, wire3290, wire3292, n_n1028, n_n1316, wire306, wire3296, n_n137, n_n1029, n_n1253, wire588, n_n935, wire184, wire209, n_n809, n_n1223, wire3299, wire218, wire197, wire270, n_n823, wire326, n_n1203, n_n1056, wire348, n_n1261, wire287, n_n1268, wire132, n_n573, n_n616, n_n617, n_n1024, n_n1025, wire568, wire76, wire114, wire128, wire162, wire243, wire298, n_n822, n_n826, wire138, wire3361, wire319, wire82, n_n1196, n_n1287, n_n1163, n_n1049, n_n1318, n_n1189, n_n1061, n_n756, n_n845, n_n215, n_n1135, wire66, n_n921, wire250, n_n468, wire140, wire297, wire98, n_n1166, wire309, wire229, wire3387, wire3388, wire333, n_n1076, n_n1077, wire337, wire237, wire139, wire3393, wire341, n_n895, wire173, wire343, n_n1181, n_n716, n_n427, n_n906, n_n1329, n_n459, n_n973, n_n1134, wire353, n_n904, n_n1037, wire3312, n_n996, n_n1033, wire483, wire87, wire216, wire3304, wire3305, wire3309, wire200, wire67, n_n909, wire261, n_n1256, n_n1229, n_n953, wire110, wire177, n_n858, wire3462, wire3464, wire182, wire279, n_n813, wire189, n_n821, wire421, wire310, wire102, wire84, n_n1283, n_n580, wire260, wire129, wire153, wire155, wire148, wire487, wire488, wire3311, wire201, wire221, n_n805, n_n1238, n_n1239, wire450, n_n803, wire3465, wire3467, wire159, n_n16, wire164, wire277, wire288, wire293, n_n1285, n_n923, n_n814, n_n1122, n_n1288, n_n963, n_n1006, n_n1204, wire86, n_n961, wire111, wire130, wire136, n_n1192, wire534, wire3535, wire154, wire253, wire274, wire434, wire276, wire291, wire305, n_n934, n_n797, wire345, n_n128, wire242, wire3573, n_n1002, wire592, wire156, wire193, n_n1074, n_n609, wire286, wire316, wire255, wire3577, wire284, n_n673, wire313, n_n1320, wire3216, wire332, n_n1010, n_n1272, n_n95, n_n1334, n_n1314, n_n1282, n_n925, n_n1013, n_n990, wire3621, wire179, wire174, wire3395, wire283, wire3359, wire238, n_n1300, wire3638, n_n490, n_n1231, wire135, wire545, wire546, n_n1258, n_n1275, n_n534, n_n926, wire266, n_n1018, n_n1301, wire64, wire83, wire183, wire109, wire112, wire247, wire257, n_n1254, n_n1330, wire268, n_n1040, n_n642, n_n574, wire3671, wire3672, wire3674, wire3676, wire259, n_n660, n_n1147, wire532, wire78, wire99, wire500, n_n1170, wire235, wire97, n_n817, wire315, n_n802, wire325, wire281, n_n1032, wire165, n_n1257, n_n745, wire181, n_n1227, wire3358, wire292, n_n1216, n_n1244, n_n554, n_n810, n_n1269, wire150, wire308, wire340, wire191, wire342, n_n1224, n_n937, wire3802, n_n711, n_n1284, wire95, wire3384, wire107, n_n1243, wire217, wire231, wire295, wire3485, wire3486, wire3804, n_n1034, wire504, wire505, n_n824, wire412, wire413, wire101, wire271, wire320, n_n1165, n_n989, n_n1322, wire106, wire3390, wire207, n_n1139, n_n553, n_n1138, wire113, wire158, wire161, n_n962, n_n799, wire3973, wire3978, wire265, n_n1155, wire466, n_n738, wire3273, wire473, wire471, wire160, wire323, wire561, n_n948, n_n1167, wire461, wire3341, wire3342, wire3348, n_n901, n_n582, n_n1148, n_n1104, n_n1119, n_n1303, n_n1023, n_n786, n_n1273, n_n1319, n_n825, wire549, wire273, n_n1153, n_n1230, wire507, wire3349, n_n1315, n_n931, n_n910, n_n792, wire515, wire3283, n_n1213, wire219, wire303, wire564, wire133, wire3363, wire493, wire414, wire426, wire456, wire462, wire468, wire512, wire3176, wire3177, wire3178, wire3195, wire3196, wire3203, wire3206, wire3236, wire3245, wire3248, wire3250, wire3251, wire3256, wire3257, wire3261, wire3262, wire3264, wire3277, wire3278, wire3279, wire3282, wire3285, wire3286, wire3287, wire3294, wire3313, wire3316, wire3317, wire3318, wire3319, wire3320, wire3321, wire3322, wire3327, wire3328, wire3329, wire3340, wire3350, wire3351, wire3353, wire3367, wire3368, wire3370, wire3373, wire3375, wire3383, wire3400, wire3404, wire3405, wire3406, wire3407, wire3408, wire3410, wire3411, wire3414, wire3420, wire3422, wire3432, wire3433, wire3434, wire3436, wire3437, wire3439, wire3440, wire3441, wire3442, wire3443, wire3447, wire3460, wire3470, wire3471, wire3472, wire3475, wire3477, wire3487, wire3488, wire3491, wire3493, wire3494, wire3495, wire3496, wire3497, wire3498, wire3505, wire3506, wire3507, wire3510, wire3511, wire3515, wire3516, wire3517, wire3518, wire3519, wire3520, wire3533, wire3541, wire3542, wire3545, wire3546, wire3548, wire3552, wire3554, wire3557, wire3558, wire3561, wire3579, wire3582, wire3585, wire3587, wire3588, wire3589, wire3590, wire3592, wire3607, wire3610, wire3612, wire3613, wire3616, wire3624, wire3628, wire3631, wire3641, wire3643, wire3644, wire3653, wire3654, wire3655, wire3667, wire3668, wire3669, wire3679, wire3682, wire3686, wire3687, wire3688, wire3689, wire3690, wire3692, wire3693, wire3695, wire3702, wire3703, wire3704, wire3712, wire3713, wire3714, wire3715, wire3716, wire3717, wire3719, wire3723, wire3724, wire3725, wire3736, wire3739, wire3754, wire3756, wire3758, wire3759, wire3760, wire3765, wire3770, wire3772, wire3774, wire3775, wire3777, wire3781, wire3782, wire3784, wire3786, wire3789, wire3792, wire3796, wire3797, wire3798, wire3800, wire3801, wire3806, wire3807, wire3808, wire3809, wire3810, wire3813, wire3816, wire3818, wire3820, wire3821, wire3822, wire3823, wire3827, wire3841, wire3842, wire3843, wire3844, wire3850, wire3853, wire3854, wire3855, wire3856, wire3857, wire3860, wire3864, wire3868, wire3870, wire3871, wire3872, wire3873, wire3874, wire3875, wire3877, wire3883, wire3890, wire3892, wire3897, wire3899, wire3900, wire3903, wire3905, wire3915, wire3916, wire3920, wire3926, wire3929, wire3937, wire3938, wire3939, wire3940, wire3941, wire3942, wire3944, wire3945, wire3950, wire3951, wire3952, wire3955, wire3957, wire3958, wire3962, wire3965, wire3975, wire3982, wire3983, wire3985, wire3993, wire3994, wire3995, wire3997, wire3998, wire4001, wire4005, wire4006, wire4007, wire4008, wire4009, wire4019, wire4020, wire4023, wire4024, wire4025, wire4027, wire4029, wire4037, wire4038, wire4039, wire4042, wire4044, wire4046, wire4047, wire4051, wire4053, wire4063, wire4065, wire4066, wire4071, wire4074, wire4076, wire4079, wire4081, wire4082, wire4083, wire4084, wire4086, wire4090, wire4091, wire4092, wire4094, wire4099, wire4100, wire4101, wire4105, wire4106, wire4109, wire4113, wire4115, wire4119, wire4122, wire4123, wire4125, wire4138, wire4139, wire4140, wire4141, wire4142, wire4144, wire4145, wire4149, wire4150, wire4151, wire4152, wire4153, wire4154, _88, _92, _94, _100, _111, _113, _115, _119, _121, _148, _173, _175, _177, _192, _225, _230, _233, _271, _302, _315, _327, _363, _420, _473, _475, _485, _540, _583, _605, _646, _713, _787, _6938, _6943, _6944, _6968, _7024, _7041, _7043, _7056, _7076, _7160, _7201, _7234, _7256, _7275, _7295, _7316, _7318, _7320, _7324, _7325, _7326, _7362, _7435, _7451, _7486, _7583, _7611, _7620, _7638, _7788, _7795, _7798, _7801, _7818, _7830, _7839, _7869, _7921, _7923, _7931, _7932, _7991, _7993, _7994, _8022, _8053, _8108, _8115, _8117, _8134, _8137, _8159, _8171, _8174, _8175, _8176, _8178, _8180, _8188, _8190, _8193, _8194, _8200, _8211, _8222, _8233, _8234, _8235, _8241, _8245, _8257, _8258, _8259, _8261, _8276, _8277, _8292, _8295, _8309, _8315, _8318, _8328, _8329, _8332, _8384, _8387, _8418, _8423, _8425, _8455, _8456, _8458, _8479, _8489, _8491, _8494, _8503, _8505, _8510, _8513, _8515, _8519, _8530, _8533, _8535, _8546, _8549, _8561, _8569, _8594, _8610, _8613, _8615, _8616, _8617, _8619, _8622, _8626, _8647, _8692, _8698, _8700, _8701, _8710, _8711, _8716, _8718, _8720, _8722, _8726, _8729, _8730, _8733, _8737, _8738, _8740, _8741, _8742, _8745, _8759, _8760, _8762, _8855, _8860, _8875, _8876, _8882, _8889, _8905, _8906, _8910, _8915, _8923, _8927, _8932, _8934, _8941, _8950, _8951, _8952, _8954, _8958, _8974, _8975, _8976, _9005, _9008, _9009, _9011, _9012, _9019, _9021, _9032, _9035, _9037, _9052, _9061, _9065, _9068, _9071, _9083, _9087, _9088, _9095, _9097, _9099, _9104, _9107, _9116, _9120, _9141, _9151, _9153, _9162, _9187, _9191;

assign o_1_ = ( wire3179 ) | ( wire3180 ) | ( wire3184 ) ;
 assign o_19_ = ( n_n744 ) | ( wire248 ) | ( n_n0  &  wire71 ) ;
 assign o_2_ = ( wire3188 ) | ( wire3189 ) | ( wire3190 ) | ( wire3191 ) ;
 assign o_0_ = ( wire3204 ) | ( wire3205 ) | ( wire3209 ) ;
 assign o_29_ = ( i_7_  &  (~ i_6_)  &  n_n0  &  n_n7 ) ;
 assign o_60_ = ( wire3266 ) | ( wire3267 ) | ( wire3268 ) | ( wire3269 ) ;
 assign o_39_ = ( n_n136 ) | ( wire3332 ) | ( wire3333 ) | ( wire3334 ) ;
 assign o_38_ = ( wire3377 ) | ( wire3378 ) | ( wire3381 ) ;
 assign o_25_ = ( (~ i_7_)  &  i_6_  &  n_n7  &  n_n2 ) ;
 assign o_12_ = ( i_7_  &  i_6_  &  n_n5  &  n_n8 ) ;
 assign o_37_ = ( wire3417 ) | ( wire3418 ) | ( wire3424 ) | ( wire3428 ) ;
 assign o_26_ = ( n_n7  &  n_n5  &  n_n17 ) | ( n_n7  &  n_n17  &  n_n19 ) ;
 assign o_11_ = ( i_7_  &  i_6_  &  n_n8  &  n_n6 ) ;
 assign o_50_ = ( wire3452 ) | ( wire3453 ) | ( wire3454 ) | ( wire3455 ) ;
 assign o_36_ = ( wire3481 ) | ( wire3477 ) | ( _8245 ) | ( _8295 ) ;
 assign o_27_ = ( (~ i_7_)  &  i_6_  &  n_n7  &  n_n3 ) ;
 assign o_14_ = ( i_7_  &  i_6_  &  n_n4  &  n_n12 ) ;
 assign o_35_ = ( wire3502 ) | ( wire3503 ) | ( wire3355 ) | ( _8235 ) ;
 assign o_28_ = ( i_7_  &  i_6_  &  n_n5  &  n_n11 ) ;
 assign o_13_ = ( i_7_  &  i_6_  &  n_n2  &  n_n12 ) ;
 assign o_34_ = ( n_n136 ) | ( wire3526 ) | ( wire3527 ) | ( wire3528 ) ;
 assign o_21_ = ( i_7_  &  (~ i_6_)  &  n_n4  &  n_n11 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n4  &  n_n11 ) ;
 assign o_16_ = ( i_7_  &  i_6_  &  n_n6  &  n_n12 ) ;
 assign o_40_ = ( wire3566 ) | ( wire3567 ) | ( wire3568 ) | ( wire3569 ) ;
 assign o_33_ = ( wire3598 ) | ( wire3599 ) | ( wire3600 ) | ( wire3601 ) ;
 assign o_22_ = ( n_n7  &  n_n17  &  n_n4 ) | ( n_n17  &  n_n4  &  n_n11 ) ;
 assign o_15_ = ( i_7_  &  i_6_  &  n_n3  &  n_n12 ) ;
 assign o_32_ = ( wire3614 ) | ( wire3615 ) | ( wire3618 ) ;
 assign o_23_ = ( n_n1017 ) | ( wire3619 ) ;
 assign o_18_ = ( i_7_  &  i_6_  &  n_n13  &  n_n1 ) | ( (~ i_7_)  &  i_6_  &  n_n13  &  n_n1 ) | ( i_7_  &  (~ i_6_)  &  n_n13  &  n_n1 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n13  &  n_n1 ) ;
 assign o_31_ = ( wire3355 ) | ( wire3631 ) | ( _8546 ) | ( _8549 ) ;
 assign o_24_ = ( (~ i_7_)  &  i_6_  &  n_n0  &  n_n7 ) ;
 assign o_17_ = ( wire180 ) | ( wire3636 ) ;
 assign o_56_ = ( wire3660 ) | ( wire3663 ) | ( _8619 ) ;
 assign o_43_ = ( n_n371 ) | ( wire3705 ) | ( wire3706 ) | ( wire3710 ) ;
 assign o_30_ = ( i_7_  &  i_6_  &  n_n7  &  n_n19 ) ;
 assign o_55_ = ( wire3733 ) | ( wire3717 ) | ( _8710 ) | ( _8718 ) ;
 assign o_44_ = ( wire3743 ) | ( wire3744 ) | ( _8733 ) ;
 assign o_58_ = ( wire3763 ) | ( wire3764 ) | ( wire3765 ) | ( _8760 ) ;
 assign o_41_ = ( wire322 ) | ( wire321 ) | ( wire3790 ) | ( wire3795 ) ;
 assign o_57_ = ( wire3829 ) | ( wire3830 ) | ( wire3831 ) | ( wire3832 ) ;
 assign o_42_ = ( wire3882 ) | ( wire3883 ) | ( _8905 ) | ( _8906 ) ;
 assign o_20_ = ( i_7_  &  (~ i_6_)  &  n_n7  &  n_n4 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n7  &  n_n4 ) ;
 assign o_52_ = ( wire3908 ) | ( wire3909 ) | ( wire3910 ) | ( wire3911 ) ;
 assign o_47_ = ( wire3925 ) | ( wire3926 ) | ( _8951 ) | ( _8952 ) ;
 assign o_51_ = ( wire3966 ) | ( wire3967 ) | ( wire3968 ) | ( wire3969 ) ;
 assign o_48_ = ( wire3355 ) | ( wire3978 ) | ( _9012 ) | ( _9021 ) ;
 assign o_54_ = ( wire4013 ) | ( wire4014 ) | ( wire4015 ) | ( wire4016 ) ;
 assign o_45_ = ( wire3355 ) | ( wire4031 ) | ( _9065 ) ;
 assign o_10_ = ( n_n8  &  n_n17  &  n_n3 ) | ( n_n17  &  n_n3  &  n_n12 ) ;
 assign o_53_ = ( wire4055 ) | ( wire4056 ) | ( wire4057 ) | ( wire4058 ) ;
 assign o_46_ = ( wire263 ) | ( wire4069 ) | ( wire4066 ) | ( _9097 ) ;
 assign o_61_ = ( wire3344 ) | ( wire3345 ) | ( wire4093 ) | ( wire4097 ) ;
 assign o_9_ = ( i_7_  &  i_6_  &  n_n7  &  n_n1 ) ;
 assign o_62_ = ( wire267 ) | ( wire347 ) | ( wire4108 ) | ( wire4112 ) ;
 assign o_49_ = ( wire3355 ) | ( wire3978 ) | ( _9012 ) | ( _9162 ) ;
 assign o_7_ = ( i_7_  &  i_6_  &  n_n2  &  n_n8 ) ;
 assign o_8_ = ( i_7_  &  i_6_  &  n_n8  &  n_n19 ) ;
 assign o_5_ = ( wire4126 ) | ( wire4127 ) | ( wire4128 ) | ( wire4129 ) ;
 assign o_59_ = ( wire4160 ) | ( wire4161 ) | ( wire4162 ) | ( wire4163 ) ;
 assign o_6_ = ( i_7_  &  (~ i_6_)  &  n_n11  &  n_n1 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n11  &  n_n1 ) ;
 assign o_3_ = ( (~ i_7_)  &  (~ i_6_)  &  n_n12 ) ;
 assign o_4_ = ( wire4166 ) | ( wire4167 ) | ( wire4168 ) | ( wire4169 ) ;
 assign wire3179 = ( n_n0  &  n_n7  &  n_n14 ) | ( n_n7  &  n_n4  &  n_n14 ) ;
 assign wire3180 = ( n_n7  &  n_n2  &  n_n14 ) | ( n_n7  &  n_n19  &  n_n14 ) ;
 assign wire3184 = ( n_n1305 ) | ( wire3176 ) | ( wire3177 ) | ( wire3178 ) ;
 assign n_n744 = ( i_7_  &  i_6_  &  n_n0  &  n_n10 ) | ( (~ i_7_)  &  i_6_  &  n_n0  &  n_n10 ) | ( i_7_  &  (~ i_6_)  &  n_n0  &  n_n10 ) ;
 assign wire248 = ( i_7_  &  (~ i_6_)  &  n_n0  &  n_n9 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n0  &  n_n9 ) ;
 assign n_n0 = ( (~ i_1_)  &  (~ i_2_)  &  (~ i_0_) ) ;
 assign wire71 = ( (~ i_7_)  &  (~ i_6_)  &  n_n10 ) | ( i_7_  &  i_6_  &  n_n9 ) | ( (~ i_7_)  &  i_6_  &  n_n9 ) ;
 assign wire3188 = ( n_n5  &  n_n8  &  n_n14 ) | ( n_n8  &  n_n19  &  n_n14 ) ;
 assign wire3189 = ( n_n2  &  n_n8  &  n_n14 ) | ( n_n8  &  n_n4  &  n_n14 ) ;
 assign wire3190 = ( n_n0  &  n_n8  &  n_n14 ) | ( n_n8  &  n_n1  &  n_n14 ) ;
 assign wire3191 = ( n_n8  &  n_n6  &  n_n14 ) | ( n_n8  &  n_n3  &  n_n14 ) ;
 assign wire3204 = ( o_20_ ) | ( n_n1320 ) | ( n_n1010 ) | ( wire135 ) ;
 assign wire3205 = ( n_n1169 ) | ( wire73 ) | ( wire92 ) | ( wire93 ) ;
 assign wire3209 = ( wire208 ) | ( wire249 ) | ( wire3203 ) | ( wire3206 ) ;
 assign n_n7 = ( (~ i_5_)  &  (~ i_3_)  &  (~ i_4_) ) ;
 assign wire3266 = ( wire240 ) | ( wire252 ) | ( wire324 ) | ( wire3250 ) ;
 assign wire3267 = ( wire3261 ) | ( wire3262 ) ;
 assign wire3268 = ( wire332 ) | ( wire3256 ) | ( _7234 ) ;
 assign wire3269 = ( wire115 ) | ( wire192 ) | ( wire3257 ) | ( wire3264 ) ;
 assign n_n136 = ( wire285 ) | ( wire3288 ) | ( wire3290 ) | ( wire3292 ) ;
 assign wire3332 = ( wire3327 ) | ( wire3328 ) | ( wire3329 ) ;
 assign wire3333 = ( n_n137 ) | ( wire200 ) | ( wire148 ) | ( wire150 ) ;
 assign wire3334 = ( wire330 ) | ( wire326 ) | ( wire221 ) | ( wire165 ) ;
 assign wire3377 = ( wire3216 ) | ( wire3370 ) | ( wire3373 ) | ( _7795 ) ;
 assign wire3378 = ( wire218 ) | ( wire189 ) | ( wire238 ) | ( wire3375 ) ;
 assign wire3381 = ( wire3355 ) | ( wire319 ) | ( _7993 ) | ( _7994 ) ;
 assign n_n2 = ( i_1_  &  (~ i_2_)  &  (~ i_0_) ) ;
 assign n_n5 = ( (~ i_1_)  &  i_2_  &  i_0_ ) ;
 assign n_n8 = ( i_5_  &  (~ i_3_)  &  (~ i_4_) ) ;
 assign wire3417 = ( wire128 ) | ( n_n845 ) | ( wire129 ) | ( wire107 ) ;
 assign wire3418 = ( wire337 ) | ( wire3216 ) | ( _8022 ) ;
 assign wire3424 = ( wire3406 ) | ( wire3407 ) | ( wire3414 ) | ( _8053 ) ;
 assign wire3428 = ( wire333 ) | ( wire3420 ) | ( wire3422 ) | ( _8159 ) ;
 assign n_n17 = ( i_7_  &  i_6_ ) ;
 assign n_n19 = ( i_1_  &  i_2_  &  i_0_ ) ;
 assign n_n6 = ( i_1_  &  (~ i_2_)  &  i_0_ ) ;
 assign wire3452 = ( n_n996 ) | ( wire87 ) | ( _8178 ) ;
 assign wire3453 = ( wire343 ) | ( wire107 ) | ( _8188 ) | ( _8190 ) ;
 assign wire3454 = ( wire3436 ) | ( wire3440 ) | ( _8211 ) ;
 assign wire3455 = ( wire330 ) | ( n_n427 ) | ( wire200 ) | ( wire3447 ) ;
 assign wire3481 = ( n_n996 ) | ( wire181 ) | ( _485 ) | ( _8259 ) ;
 assign wire3482 = ( wire182 ) | ( wire3475 ) | ( _8292 ) ;
 assign n_n3 = ( i_1_  &  i_2_  &  (~ i_0_) ) ;
 assign n_n4 = ( (~ i_1_)  &  (~ i_2_)  &  i_0_ ) ;
 assign n_n12 = ( i_5_  &  i_3_  &  (~ i_4_) ) ;
 assign wire3502 = ( wire181 ) | ( wire3460 ) | ( wire3494 ) | ( wire3495 ) ;
 assign wire3503 = ( wire318 ) | ( wire3496 ) | ( wire3497 ) | ( wire3498 ) ;
 assign n_n11 = ( (~ i_5_)  &  i_3_  &  (~ i_4_) ) ;
 assign wire3526 = ( wire216 ) | ( wire310 ) | ( _8329 ) | ( _8332 ) ;
 assign wire3527 = ( wire3516 ) | ( wire3517 ) | ( wire3518 ) | ( wire3519 ) ;
 assign wire3528 = ( wire301 ) | ( n_n137 ) | ( wire3520 ) ;
 assign wire3566 = ( wire87 ) | ( wire3533 ) | ( _8384 ) | ( _8387 ) ;
 assign wire3567 = ( wire154 ) | ( wire305 ) | ( wire3554 ) | ( wire3561 ) ;
 assign wire3568 = ( wire3436 ) | ( wire3557 ) | ( _8423 ) ;
 assign wire3569 = ( wire341 ) | ( n_n427 ) | ( n_n1006 ) | ( wire3558 ) ;
 assign wire3598 = ( wire229 ) | ( wire345 ) | ( n_n642 ) | ( wire3592 ) ;
 assign wire3599 = ( wire87 ) | ( wire3585 ) | ( _7788 ) | ( _8458 ) ;
 assign wire3600 = ( wire193 ) | ( wire255 ) | ( wire313 ) | ( wire3587 ) ;
 assign wire3601 = ( wire332 ) | ( wire3588 ) | ( wire3589 ) | ( wire3590 ) ;
 assign wire3614 = ( wire200 ) | ( wire148 ) | ( wire150 ) | ( wire3612 ) ;
 assign wire3615 = ( wire343 ) | ( wire3607 ) | ( _8513 ) ;
 assign wire3618 = ( wire3355 ) | ( wire3344 ) | ( wire3345 ) | ( wire3616 ) ;
 assign n_n1017 = ( (~ i_7_)  &  i_6_  &  n_n0  &  n_n12 ) | ( i_7_  &  (~ i_6_)  &  n_n0  &  n_n12 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n0  &  n_n12 ) ;
 assign wire3619 = ( n_n0  &  n_n18 ) | ( n_n0  &  n_n17  &  n_n12 ) ;
 assign n_n13 = ( (~ i_5_)  &  i_3_  &  i_4_ ) ;
 assign n_n1 = ( (~ i_1_)  &  i_2_  &  (~ i_0_) ) ;
 assign wire318 = ( wire270 ) | ( n_n826 ) | ( _7932 ) ;
 assign wire3605 = ( wire180 ) | ( n_n955 ) | ( wire273 ) | ( _8515 ) ;
 assign wire180 = ( i_7_  &  i_6_  &  n_n4  &  n_n13 ) | ( (~ i_7_)  &  i_6_  &  n_n4  &  n_n13 ) | ( i_7_  &  (~ i_6_)  &  n_n4  &  n_n13 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n4  &  n_n13 ) ;
 assign wire3636 = ( i_7_  &  i_6_  &  n_n4  &  n_n9 ) | ( (~ i_7_)  &  i_6_  &  n_n4  &  n_n9 ) | ( i_7_  &  (~ i_6_)  &  n_n4  &  n_n9 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n4  &  n_n9 ) ;
 assign wire322 = ( wire189 ) | ( n_n814 ) | ( wire97 ) | ( n_n817 ) ;
 assign wire3639 = ( wire3638 ) | ( n_n3  &  n_n13  &  wire64 ) ;
 assign wire3660 = ( wire177 ) | ( wire332 ) | ( wire3641 ) | ( wire3653 ) ;
 assign wire3663 = ( wire3355 ) | ( wire3655 ) | ( _8616 ) | ( _8617 ) ;
 assign n_n371 = ( wire3671 ) | ( wire3672 ) | ( wire3674 ) | ( wire3676 ) ;
 assign wire3705 = ( n_n387 ) | ( wire305 ) | ( n_n642 ) | ( wire3690 ) ;
 assign wire3706 = ( n_n574 ) | ( wire3692 ) | ( _8647 ) ;
 assign wire3710 = ( wire314 ) | ( wire3702 ) | ( wire3703 ) | ( wire3704 ) ;
 assign wire3733 = ( wire3723 ) | ( wire3724 ) | ( _8716 ) ;
 assign wire3743 = ( wire270 ) | ( wire333 ) | ( _8261 ) | ( _8720 ) ;
 assign wire3744 = ( wire267 ) | ( wire86 ) | ( wire193 ) | ( wire3736 ) ;
 assign wire3745 = ( wire314 ) | ( wire3739 ) | ( _8730 ) ;
 assign wire3763 = ( wire194 ) | ( wire3440 ) | ( wire3760 ) | ( _8200 ) ;
 assign wire3764 = ( n_n996 ) | ( wire345 ) | ( _8722 ) | ( _8742 ) ;
 assign wire321 = ( n_n845 ) | ( n_n858 ) | ( wire3462 ) | ( wire3464 ) ;
 assign wire3790 = ( wire342 ) | ( wire3341 ) | ( wire3342 ) | ( wire3786 ) ;
 assign wire3795 = ( wire200 ) | ( wire238 ) | ( wire3789 ) | ( wire3792 ) ;
 assign wire3829 = ( wire327 ) | ( n_n711 ) | ( wire231 ) | ( wire3823 ) ;
 assign wire3830 = ( n_n660 ) | ( wire295 ) | ( wire3813 ) | ( wire3818 ) ;
 assign wire3831 = ( wire347 ) | ( n_n427 ) | ( wire3820 ) ;
 assign wire3832 = ( wire3821 ) | ( wire3822 ) | ( wire3827 ) ;
 assign wire314 = ( wire85 ) | ( n_n1021 ) | ( n_n1020 ) | ( wire153 ) ;
 assign wire3882 = ( wire3870 ) | ( wire3871 ) | ( wire3877 ) ;
 assign wire3908 = ( n_n1008 ) | ( wire136 ) | ( _8910 ) | ( _8915 ) ;
 assign wire3909 = ( wire139 ) | ( wire154 ) | ( wire3903 ) | ( wire3905 ) ;
 assign wire3910 = ( wire218 ) | ( wire189 ) | ( wire238 ) | ( _8927 ) ;
 assign wire3911 = ( wire319 ) | ( wire3892 ) | ( _8934 ) ;
 assign wire3921 = ( n_n459 ) | ( wire129 ) | ( wire107 ) ;
 assign wire3925 = ( wire200 ) | ( wire201 ) | ( wire3439 ) | ( wire3440 ) ;
 assign wire3966 = ( wire252 ) | ( wire3296 ) | ( _8711 ) | ( _8954 ) ;
 assign wire3967 = ( wire342 ) | ( wire3950 ) | ( wire3951 ) | ( wire3952 ) ;
 assign wire3968 = ( wire3944 ) | ( wire3945 ) | ( wire3955 ) | ( wire3962 ) ;
 assign wire3969 = ( wire3957 ) | ( wire3958 ) | ( wire3965 ) ;
 assign n_n476 = ( wire138 ) | ( n_n574 ) | ( n_n799 ) | ( wire3973 ) ;
 assign wire263 = ( wire3355 ) | ( wire3978 ) | ( _9012 ) ;
 assign wire264 = ( n_n990 ) | ( n_n0  &  wire72 ) ;
 assign wire4013 = ( wire4008 ) | ( wire4009 ) ;
 assign wire4014 = ( n_n468 ) | ( wire3717 ) | ( _9032 ) | ( _9037 ) ;
 assign wire4015 = ( wire347 ) | ( wire3462 ) | ( wire3464 ) | ( _8762 ) ;
 assign wire4016 = ( n_n1006 ) | ( wire4005 ) | ( wire4006 ) | ( wire4007 ) ;
 assign wire3355 = ( n_n427 ) | ( n_n609 ) | ( wire3350 ) | ( wire3353 ) ;
 assign wire4031 = ( wire322 ) | ( wire267 ) | ( wire4027 ) | ( wire4029 ) ;
 assign wire4055 = ( wire140 ) | ( wire325 ) | ( _9068 ) | ( _9071 ) ;
 assign wire4056 = ( wire4046 ) | ( wire4047 ) | ( wire4051 ) ;
 assign wire4057 = ( wire154 ) | ( wire97 ) | ( _8701 ) | ( _9088 ) ;
 assign wire4058 = ( wire115 ) | ( wire192 ) | ( wire255 ) | ( wire4053 ) ;
 assign wire4069 = ( wire138 ) | ( wire4065 ) | ( _92 ) | ( _9104 ) ;
 assign wire3344 = ( wire461 ) | ( wire3341 ) | ( wire3342 ) ;
 assign wire3345 = ( _7931 ) | ( n_n10  &  wire93 ) | ( n_n10  &  wire466 ) ;
 assign wire4093 = ( wire343 ) | ( wire3607 ) | ( _9107 ) ;
 assign wire4097 = ( wire4091 ) | ( wire4092 ) | ( wire4094 ) ;
 assign wire267 = ( n_n996 ) | ( wire345 ) | ( n_n1040 ) | ( n_n1257 ) ;
 assign wire347 = ( n_n1002 ) | ( wire3485 ) | ( wire3486 ) | ( wire3804 ) ;
 assign wire4108 = ( n_n990 ) | ( wire3892 ) | ( _100 ) | ( _9141 ) ;
 assign wire4112 = ( wire4105 ) | ( wire4106 ) | ( wire4109 ) ;
 assign wire4117 = ( wire139 ) | ( wire129 ) | ( wire107 ) | ( wire4115 ) ;
 assign wire4126 = ( n_n1300 ) | ( n_n1315 ) | ( wire4119 ) ;
 assign wire4127 = ( n_n1269 ) | ( n_n1224 ) | ( n_n1284 ) | ( n_n1148 ) ;
 assign wire4128 = ( wire4122 ) | ( wire4123 ) ;
 assign wire4129 = ( n_n1133 ) | ( n_n1119 ) | ( wire4125 ) ;
 assign wire4160 = ( wire323 ) | ( n_n786 ) | ( wire4154 ) ;
 assign wire4161 = ( wire4149 ) | ( wire4150 ) | ( wire4151 ) | ( wire4152 ) ;
 assign wire4162 = ( wire218 ) | ( wire189 ) | ( wire238 ) | ( wire315 ) ;
 assign wire4163 = ( wire326 ) | ( wire193 ) | ( n_n989 ) | ( wire4153 ) ;
 assign wire4166 = ( n_n4  &  n_n11  &  n_n16 ) | ( n_n11  &  n_n1  &  n_n16 ) ;
 assign wire4167 = ( n_n2  &  n_n11  &  n_n16 ) | ( n_n5  &  n_n11  &  n_n16 ) ;
 assign wire4168 = ( n_n6  &  n_n11  &  n_n16 ) | ( n_n3  &  n_n11  &  n_n16 ) ;
 assign wire4169 = ( n_n0  &  n_n11  &  n_n16 ) | ( n_n19  &  n_n11  &  n_n16 ) ;
 assign n_n1154 = ( (~ i_7_)  &  (~ i_6_)  &  n_n7  &  n_n6 ) ;
 assign n_n1245 = ( (~ i_7_)  &  (~ i_6_)  &  n_n7  &  n_n3 ) ;
 assign n_n1215 = ( (~ i_7_)  &  (~ i_6_)  &  n_n7  &  n_n4 ) ;
 assign n_n1274 = ( (~ i_7_)  &  (~ i_6_)  &  n_n7  &  n_n2 ) ;
 assign n_n1305 = ( (~ i_7_)  &  (~ i_6_)  &  n_n7  &  n_n1 ) ;
 assign n_n10 = ( i_5_  &  (~ i_3_)  &  i_4_ ) ;
 assign n_n9 = ( (~ i_5_)  &  (~ i_3_)  &  i_4_ ) ;
 assign n_n1121 = ( (~ i_7_)  &  (~ i_6_)  &  n_n8  &  n_n19 ) ;
 assign n_n1180 = ( (~ i_7_)  &  (~ i_6_)  &  n_n5  &  n_n8 ) ;
 assign n_n1211 = ( (~ i_7_)  &  (~ i_6_)  &  n_n8  &  n_n4 ) ;
 assign n_n1271 = ( (~ i_7_)  &  (~ i_6_)  &  n_n2  &  n_n8 ) ;
 assign n_n1302 = ( (~ i_7_)  &  (~ i_6_)  &  n_n8  &  n_n1 ) ;
 assign wire246 = ( (~ i_7_)  &  (~ i_6_)  &  n_n8  &  n_n3 ) ;
 assign wire354 = ( (~ i_7_)  &  (~ i_6_)  &  n_n8  &  n_n6 ) ;
 assign n_n1168 = ( i_7_  &  (~ i_6_)  &  n_n5  &  n_n11 ) ;
 assign n_n1321 = ( (~ i_7_)  &  (~ i_6_)  &  n_n0  &  n_n11 ) ;
 assign n_n1169 = ( (~ i_7_)  &  (~ i_6_)  &  n_n5  &  n_n11 ) ;
 assign wire73 = ( i_7_  &  (~ i_6_)  &  n_n19  &  n_n11 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n19  &  n_n11 ) ;
 assign wire92 = ( i_7_  &  (~ i_6_)  &  n_n7  &  n_n6 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n7  &  n_n6 ) ;
 assign wire93 = ( i_7_  &  (~ i_6_)  &  n_n6  &  n_n11 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n6  &  n_n11 ) ;
 assign wire94 = ( i_7_  &  (~ i_6_)  &  n_n7  &  n_n19 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n7  &  n_n19 ) ;
 assign wire146 = ( i_7_  &  (~ i_6_)  &  n_n7  &  n_n3 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n7  &  n_n3 ) ;
 assign wire147 = ( i_7_  &  (~ i_6_)  &  n_n2  &  n_n11 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n2  &  n_n11 ) ;
 assign wire186 = ( i_7_  &  (~ i_6_)  &  n_n7  &  n_n5 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n7  &  n_n5 ) ;
 assign wire208 = ( i_7_  &  (~ i_6_)  &  n_n7  &  n_n2 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n7  &  n_n2 ) ;
 assign wire249 = ( i_7_  &  (~ i_6_)  &  n_n7  &  n_n1 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n7  &  n_n1 ) ;
 assign n_n1120 = ( i_7_  &  (~ i_6_)  &  n_n8  &  n_n19 ) ;
 assign n_n1083 = ( (~ i_7_)  &  i_6_  &  n_n19  &  n_n12 ) | ( i_7_  &  (~ i_6_)  &  n_n19  &  n_n12 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n19  &  n_n12 ) ;
 assign wire236 = ( i_7_  &  i_6_  &  n_n19  &  n_n11 ) | ( (~ i_7_)  &  i_6_  &  n_n19  &  n_n11 ) | ( i_7_  &  (~ i_6_)  &  n_n19  &  n_n11 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n19  &  n_n11 ) ;
 assign wire3213 = ( i_7_  &  i_6_  &  n_n8  &  n_n19 ) | ( (~ i_7_)  &  i_6_  &  n_n8  &  n_n19 ) ;
 assign n_n1008 = ( n_n1083 ) | ( wire236 ) | ( wire3213 ) ;
 assign wire163 = ( i_5_  &  i_3_  &  i_4_ ) | ( (~ i_5_)  &  i_3_  &  i_4_ ) ;
 assign n_n1009 = ( n_n19  &  wire163 ) | ( n_n17  &  n_n19  &  n_n12 ) ;
 assign n_n18 = ( i_5_  &  i_3_  &  i_4_ ) ;
 assign n_n872 = ( i_7_  &  i_6_  &  n_n6  &  n_n18 ) | ( (~ i_7_)  &  i_6_  &  n_n6  &  n_n18 ) | ( i_7_  &  (~ i_6_)  &  n_n6  &  n_n18 ) ;
 assign n_n958 = ( (~ i_7_)  &  i_6_  &  n_n4  &  n_n18 ) | ( i_7_  &  (~ i_6_)  &  n_n4  &  n_n18 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n4  &  n_n18 ) ;
 assign n_n949 = ( i_7_  &  i_6_  &  n_n7  &  n_n4 ) | ( (~ i_7_)  &  i_6_  &  n_n7  &  n_n4 ) | ( i_7_  &  (~ i_6_)  &  n_n7  &  n_n4 ) ;
 assign n_n1137 = ( (~ i_7_)  &  i_6_  &  n_n6  &  n_n11 ) ;
 assign n_n14 = ( (~ i_7_)  &  (~ i_6_) ) ;
 assign wire108 = ( _173 ) | ( n_n6  &  n_n11  &  _7316 ) ;
 assign wire85 = ( wire266 ) | ( n_n0  &  wire69 ) | ( n_n0  &  wire102 ) ;
 assign n_n1021 = ( (~ i_7_)  &  i_6_  &  n_n7  &  n_n1 ) | ( i_7_  &  (~ i_6_)  &  n_n7  &  n_n1 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n7  &  n_n1 ) ;
 assign n_n1020 = ( i_7_  &  i_6_  &  n_n0  &  n_n18 ) | ( (~ i_7_)  &  i_6_  &  n_n0  &  n_n18 ) | ( i_7_  &  (~ i_6_)  &  n_n0  &  n_n18 ) ;
 assign wire115 = ( wire85 ) | ( n_n1021 ) | ( n_n1020 ) ;
 assign n_n15 = ( i_7_  &  (~ i_6_) ) ;
 assign n_n1136 = ( i_7_  &  i_6_  &  n_n6  &  n_n11 ) ;
 assign wire152 = ( _192 ) | ( n_n6  &  n_n11  &  _7318 ) ;
 assign n_n864 = ( i_7_  &  i_6_  &  n_n5  &  n_n18 ) | ( (~ i_7_)  &  i_6_  &  n_n5  &  n_n18 ) | ( i_7_  &  (~ i_6_)  &  n_n5  &  n_n18 ) ;
 assign wire69 = ( i_7_  &  i_6_  &  n_n13 ) | ( (~ i_7_)  &  i_6_  &  n_n13 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n18 ) ;
 assign wire187 = ( n_n864 ) | ( n_n5  &  wire69 ) ;
 assign n_n602 = ( o_6_ ) | ( n_n1024 ) | ( n_n1025 ) | ( wire568 ) ;
 assign n_n1022 = ( o_9_ ) | ( n_n1302 ) | ( n_n1301 ) ;
 assign n_n1298 = ( (~ i_7_)  &  (~ i_6_)  &  n_n1  &  n_n9 ) ;
 assign wire3218 = ( i_7_  &  i_6_  &  n_n8  &  n_n1 ) | ( (~ i_7_)  &  i_6_  &  n_n8  &  n_n1 ) ;
 assign wire192 = ( n_n602 ) | ( n_n1022 ) | ( n_n1298 ) | ( wire3218 ) ;
 assign wire222 = ( i_7_  &  i_6_  &  n_n8  &  n_n6 ) | ( (~ i_7_)  &  i_6_  &  n_n8  &  n_n6 ) | ( i_7_  &  (~ i_6_)  &  n_n8  &  n_n6 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n8  &  n_n6 ) ;
 assign n_n930 = ( (~ i_7_)  &  i_6_  &  n_n2  &  n_n9 ) | ( i_7_  &  (~ i_6_)  &  n_n2  &  n_n9 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n2  &  n_n9 ) ;
 assign wire72 = ( i_7_  &  (~ i_6_)  &  n_n10 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n10 ) | ( i_7_  &  i_6_  &  n_n9 ) ;
 assign wire226 = ( n_n930 ) | ( n_n2  &  wire72 ) ;
 assign wire104 = ( (~ i_7_)  &  i_6_  &  n_n3  &  n_n12 ) | ( i_7_  &  (~ i_6_)  &  n_n3  &  n_n12 ) ;
 assign n_n1226 = ( (~ i_7_)  &  (~ i_6_)  &  n_n3  &  n_n12 ) ;
 assign wire77 = ( i_7_  &  i_6_  &  n_n3  &  n_n11 ) | ( (~ i_7_)  &  i_6_  &  n_n3  &  n_n11 ) ;
 assign wire228 = ( wire77 ) | ( _7056 ) ;
 assign wire70 = ( i_7_  &  i_6_  &  n_n13 ) | ( i_7_  &  (~ i_6_)  &  n_n18 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n18 ) ;
 assign wire3221 = ( (~ i_7_)  &  i_6_  &  n_n3  &  n_n13 ) | ( i_7_  &  (~ i_6_)  &  n_n3  &  n_n13 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n3  &  n_n13 ) ;
 assign wire3222 = ( o_15_ ) | ( n_n1215 ) | ( _6938 ) ;
 assign wire240 = ( _6943 ) | ( n_n3  &  wire70 ) ;
 assign n_n1197 = ( (~ i_7_)  &  i_6_  &  n_n4  &  n_n11 ) ;
 assign wire88 = ( i_7_  &  i_6_  &  n_n4  &  n_n12 ) | ( (~ i_7_)  &  i_6_  &  n_n4  &  n_n12 ) ;
 assign n_n955 = ( n_n1194 ) | ( n_n1196 ) | ( wire242 ) ;
 assign wire3225 = ( wire180 ) | ( n_n4  &  n_n11  &  wire66 ) ;
 assign wire252 = ( wire180 ) | ( n_n955 ) | ( _787 ) | ( _6968 ) ;
 assign n_n950 = ( (~ i_7_)  &  i_6_  &  n_n8  &  n_n4 ) | ( i_7_  &  (~ i_6_)  &  n_n8  &  n_n4 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n8  &  n_n4 ) ;
 assign n_n1208 = ( i_7_  &  i_6_  &  n_n8  &  n_n4 ) ;
 assign wire551 = ( i_7_  &  (~ i_6_)  &  n_n4  &  n_n9 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n4  &  n_n9 ) ;
 assign wire280 = ( n_n950 ) | ( n_n1208 ) | ( wire551 ) ;
 assign wire254 = ( i_7_  &  i_6_  &  n_n7  &  n_n2 ) | ( (~ i_7_)  &  i_6_  &  n_n7  &  n_n2 ) | ( i_7_  &  (~ i_6_)  &  n_n7  &  n_n2 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n7  &  n_n2 ) ;
 assign wire269 = ( i_7_  &  i_6_  &  n_n1  &  n_n18 ) | ( (~ i_7_)  &  i_6_  &  n_n1  &  n_n18 ) | ( i_7_  &  (~ i_6_)  &  n_n1  &  n_n18 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n1  &  n_n18 ) ;
 assign wire301 = ( o_18_ ) | ( n_n1271 ) | ( wire254 ) | ( wire269 ) ;
 assign wire194 = ( n_n1180 ) | ( n_n961 ) | ( wire271 ) | ( n_n962 ) ;
 assign n_n859 = ( n_n1169 ) | ( n_n1170 ) | ( wire549 ) ;
 assign wire324 = ( wire194 ) | ( n_n859 ) | ( n_n5  &  wire72 ) ;
 assign wire134 = ( i_7_  &  i_6_  &  n_n7  &  n_n19 ) | ( (~ i_7_)  &  i_6_  &  n_n7  &  n_n19 ) ;
 assign wire327 = ( n_n1121 ) | ( wire94 ) | ( wire134 ) ;
 assign n_n387 = ( n_n1231 ) | ( wire135 ) | ( wire545 ) | ( wire546 ) ;
 assign wire3237 = ( n_n1238 ) | ( n_n1239 ) | ( n_n937 ) ;
 assign wire3238 = ( wire246 ) | ( wire109 ) | ( n_n1243 ) | ( wire3236 ) ;
 assign wire330 = ( n_n387 ) | ( wire3237 ) | ( wire3238 ) ;
 assign wire300 = ( i_7_  &  i_6_  &  n_n2  &  n_n10 ) | ( (~ i_7_)  &  i_6_  &  n_n2  &  n_n10 ) ;
 assign wire127 = ( i_7_  &  i_6_  &  n_n2  &  n_n11 ) | ( (~ i_7_)  &  i_6_  &  n_n2  &  n_n11 ) ;
 assign wire331 = ( wire147 ) | ( wire300 ) | ( wire127 ) ;
 assign n_n1133 = ( (~ i_7_)  &  i_6_  &  n_n6  &  n_n12 ) ;
 assign wire3239 = ( n_n6  &  n_n13 ) | ( n_n17  &  n_n6  &  n_n12 ) ;
 assign wire346 = ( n_n1133 ) | ( wire3239 ) | ( n_n6  &  wire69 ) ;
 assign n_n1193 = ( (~ i_7_)  &  i_6_  &  n_n4  &  n_n12 ) ;
 assign n_n1225 = ( i_7_  &  (~ i_6_)  &  n_n3  &  n_n12 ) ;
 assign n_n936 = ( i_1_  &  (~ i_2_)  &  (~ i_0_)  &  wire69 ) ;
 assign n_n1194 = ( i_7_  &  (~ i_6_)  &  n_n4  &  n_n12 ) ;
 assign wire285 = ( n_n468 ) | ( wire140 ) | ( _7435 ) ;
 assign wire3288 = ( wire297 ) | ( wire3279 ) | ( wire3286 ) ;
 assign wire3290 = ( n_n1009 ) | ( n_n786 ) | ( wire515 ) | ( wire3283 ) ;
 assign wire3292 = ( wire337 ) | ( wire323 ) | ( wire3277 ) | ( wire3287 ) ;
 assign n_n1028 = ( i_7_  &  i_6_  &  n_n12  &  n_n1 ) | ( (~ i_7_)  &  i_6_  &  n_n12  &  n_n1 ) | ( i_7_  &  (~ i_6_)  &  n_n12  &  n_n1 ) ;
 assign n_n1316 = ( i_7_  &  (~ i_6_)  &  n_n0  &  n_n12 ) ;
 assign wire306 = ( wire76 ) | ( n_n1322 ) | ( _7611 ) ;
 assign wire3296 = ( n_n906 ) | ( n_n1329 ) | ( n_n909 ) | ( n_n910 ) ;
 assign n_n137 = ( wire306 ) | ( wire3296 ) | ( _7638 ) ;
 assign n_n1029 = ( (~ i_7_)  &  i_6_  &  n_n13  &  n_n1 ) | ( i_7_  &  (~ i_6_)  &  n_n13  &  n_n1 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n13  &  n_n1 ) ;
 assign n_n1253 = ( (~ i_7_)  &  (~ i_6_)  &  n_n2  &  n_n13 ) ;
 assign wire588 = ( i_7_  &  (~ i_6_)  &  n_n2  &  n_n13 ) ;
 assign n_n935 = ( o_13_ ) | ( n_n1253 ) | ( wire588 ) ;
 assign wire184 = ( (~ i_7_)  &  i_6_  &  n_n2  &  n_n12 ) | ( i_7_  &  (~ i_6_)  &  n_n2  &  n_n12 ) ;
 assign wire209 = ( i_7_  &  i_6_  &  n_n3  &  n_n12 ) | ( (~ i_7_)  &  i_6_  &  n_n3  &  n_n12 ) ;
 assign n_n809 = ( i_7_  &  i_6_  &  n_n3  &  n_n13 ) | ( (~ i_7_)  &  i_6_  &  n_n3  &  n_n13 ) | ( i_7_  &  (~ i_6_)  &  n_n3  &  n_n13 ) ;
 assign n_n1223 = ( (~ i_7_)  &  (~ i_6_)  &  n_n3  &  n_n13 ) ;
 assign wire3299 = ( i_7_  &  i_6_  &  n_n3  &  n_n18 ) | ( (~ i_7_)  &  i_6_  &  n_n3  &  n_n18 ) | ( i_7_  &  (~ i_6_)  &  n_n3  &  n_n18 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n3  &  n_n18 ) ;
 assign wire218 = ( wire209 ) | ( n_n809 ) | ( n_n1223 ) | ( wire3299 ) ;
 assign wire197 = ( n_n822 ) | ( n_n821 ) | ( wire291 ) | ( wire500 ) ;
 assign wire270 = ( o_12_ ) | ( wire504 ) | ( wire505 ) | ( n_n825 ) ;
 assign n_n823 = ( n_n1180 ) | ( n_n1181 ) | ( wire507 ) ;
 assign wire326 = ( wire197 ) | ( wire270 ) | ( n_n823 ) ;
 assign n_n1203 = ( (~ i_7_)  &  (~ i_6_)  &  n_n4  &  n_n10 ) ;
 assign n_n1056 = ( i_7_  &  i_6_  &  n_n4  &  n_n9 ) | ( (~ i_7_)  &  i_6_  &  n_n4  &  n_n9 ) | ( i_7_  &  (~ i_6_)  &  n_n4  &  n_n9 ) ;
 assign wire348 = ( n_n1056 ) | ( _7583 ) ;
 assign n_n1261 = ( i_7_  &  i_6_  &  n_n2  &  n_n10 ) ;
 assign wire287 = ( i_7_  &  i_6_  &  n_n7  &  n_n2 ) | ( (~ i_7_)  &  i_6_  &  n_n7  &  n_n2 ) | ( i_7_  &  (~ i_6_)  &  n_n7  &  n_n2 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n7  &  n_n2 ) ;
 assign n_n1268 = ( (~ i_7_)  &  (~ i_6_)  &  n_n2  &  n_n9 ) ;
 assign wire132 = ( i_7_  &  i_6_  &  n_n2  &  n_n8 ) | ( (~ i_7_)  &  i_6_  &  n_n2  &  n_n8 ) | ( i_7_  &  (~ i_6_)  &  n_n2  &  n_n8 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n2  &  n_n8 ) ;
 assign n_n573 = ( wire287 ) | ( n_n1268 ) | ( wire132 ) ;
 assign n_n616 = ( i_7_  &  i_6_  &  n_n2  &  n_n9 ) | ( (~ i_7_)  &  i_6_  &  n_n2  &  n_n9 ) | ( i_7_  &  (~ i_6_)  &  n_n2  &  n_n9 ) ;
 assign n_n617 = ( (~ i_7_)  &  i_6_  &  n_n2  &  n_n10 ) | ( i_7_  &  (~ i_6_)  &  n_n2  &  n_n10 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n2  &  n_n10 ) ;
 assign n_n1024 = ( i_7_  &  i_6_  &  n_n1  &  n_n9 ) | ( (~ i_7_)  &  i_6_  &  n_n1  &  n_n9 ) | ( i_7_  &  (~ i_6_)  &  n_n1  &  n_n9 ) ;
 assign n_n1025 = ( (~ i_7_)  &  i_6_  &  n_n1  &  n_n10 ) | ( i_7_  &  (~ i_6_)  &  n_n1  &  n_n10 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n1  &  n_n10 ) ;
 assign wire568 = ( i_7_  &  i_6_  &  n_n1  &  n_n10 ) ;
 assign wire76 = ( i_7_  &  i_6_  &  n_n0  &  n_n11 ) | ( (~ i_7_)  &  i_6_  &  n_n0  &  n_n11 ) ;
 assign wire114 = ( n_n1017 ) | ( wire76 ) ;
 assign wire128 = ( i_7_  &  i_6_  &  n_n0  &  n_n8 ) | ( (~ i_7_)  &  i_6_  &  n_n0  &  n_n8 ) | ( i_7_  &  (~ i_6_)  &  n_n0  &  n_n8 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n0  &  n_n8 ) ;
 assign wire162 = ( i_7_  &  i_6_  &  n_n11  &  n_n1 ) | ( (~ i_7_)  &  i_6_  &  n_n11  &  n_n1 ) ;
 assign wire243 = ( (~ i_7_)  &  (~ i_6_)  &  n_n12  &  n_n1 ) ;
 assign wire298 = ( n_n1028 ) | ( wire162 ) | ( wire243 ) ;
 assign n_n822 = ( (~ i_7_)  &  i_6_  &  n_n7  &  n_n5 ) | ( i_7_  &  (~ i_6_)  &  n_n7  &  n_n5 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n7  &  n_n5 ) ;
 assign n_n826 = ( (~ i_7_)  &  i_6_  &  n_n5  &  n_n10 ) | ( i_7_  &  (~ i_6_)  &  n_n5  &  n_n10 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n5  &  n_n10 ) ;
 assign wire138 = ( wire127 ) | ( n_n1256 ) | ( n_n797 ) | ( wire3363 ) ;
 assign wire3361 = ( n_n1244 ) | ( n_n2  &  wire70 ) ;
 assign wire319 = ( wire138 ) | ( wire3361 ) | ( _7991 ) ;
 assign wire82 = ( i_7_  &  i_6_  &  n_n8 ) ;
 assign n_n1196 = ( i_7_  &  i_6_  &  n_n4  &  n_n11 ) ;
 assign n_n1287 = ( i_7_  &  i_6_  &  n_n11  &  n_n1 ) ;
 assign n_n1163 = ( i_7_  &  i_6_  &  n_n5  &  n_n12 ) ;
 assign n_n1049 = ( (~ i_7_)  &  i_6_  &  n_n3  &  n_n12 ) | ( i_7_  &  (~ i_6_)  &  n_n3  &  n_n12 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n3  &  n_n12 ) ;
 assign n_n1318 = ( i_7_  &  i_6_  &  n_n0  &  n_n11 ) ;
 assign n_n1189 = ( i_7_  &  i_6_  &  n_n4  &  n_n13 ) ;
 assign n_n1061 = ( (~ i_7_)  &  i_6_  &  n_n4  &  n_n13 ) | ( i_7_  &  (~ i_6_)  &  n_n4  &  n_n13 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n4  &  n_n13 ) ;
 assign n_n756 = ( i_7_  &  i_6_  &  n_n19  &  n_n10 ) | ( (~ i_7_)  &  i_6_  &  n_n19  &  n_n10 ) | ( i_7_  &  (~ i_6_)  &  n_n19  &  n_n10 ) ;
 assign n_n845 = ( i_7_  &  i_6_  &  n_n0  &  n_n7 ) | ( (~ i_7_)  &  i_6_  &  n_n0  &  n_n7 ) | ( i_7_  &  (~ i_6_)  &  n_n0  &  n_n7 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n0  &  n_n7 ) ;
 assign n_n215 = ( wire128 ) | ( n_n845 ) ;
 assign n_n1135 = ( (~ i_7_)  &  (~ i_6_)  &  n_n6  &  n_n12 ) ;
 assign wire66 = ( i_7_  &  (~ i_6_) ) | ( (~ i_7_)  &  (~ i_6_) ) ;
 assign n_n921 = ( i_7_  &  i_6_  &  n_n1  &  n_n10 ) | ( (~ i_7_)  &  i_6_  &  n_n1  &  n_n10 ) | ( i_7_  &  (~ i_6_)  &  n_n1  &  n_n10 ) ;
 assign wire250 = ( n_n921 ) | ( n_n11  &  n_n1  &  wire66 ) ;
 assign n_n468 = ( wire3273 ) | ( n_n6  &  n_n18 ) | ( n_n6  &  wire70 ) ;
 assign wire140 = ( wire113 ) | ( wire71  &  n_n19 ) ;
 assign wire297 = ( n_n5  &  n_n13 ) | ( n_n5  &  wire70 ) ;
 assign wire98 = ( (~ i_7_)  &  i_6_  &  n_n5  &  n_n12 ) | ( i_7_  &  (~ i_6_)  &  n_n5  &  n_n12 ) ;
 assign n_n1166 = ( (~ i_7_)  &  (~ i_6_)  &  n_n5  &  n_n12 ) ;
 assign wire309 = ( o_28_ ) | ( wire98 ) | ( n_n1166 ) ;
 assign wire229 = ( wire112 ) | ( _8108 ) ;
 assign wire3387 = ( wire146 ) | ( n_n3  &  wire72 ) ;
 assign wire3388 = ( n_n1238 ) | ( n_n1239 ) | ( wire434 ) | ( wire268 ) ;
 assign wire333 = ( wire3387 ) | ( wire3388 ) | ( _8134 ) ;
 assign n_n1076 = ( i_7_  &  i_6_  &  n_n6  &  n_n12 ) | ( (~ i_7_)  &  i_6_  &  n_n6  &  n_n12 ) | ( i_7_  &  (~ i_6_)  &  n_n6  &  n_n12 ) ;
 assign n_n1077 = ( (~ i_7_)  &  i_6_  &  n_n6  &  n_n13 ) | ( i_7_  &  (~ i_6_)  &  n_n6  &  n_n13 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n6  &  n_n13 ) ;
 assign wire337 = ( n_n1136 ) | ( n_n1076 ) | ( n_n1077 ) ;
 assign wire237 = ( wire174 ) | ( wire3395 ) | ( n_n0  &  wire70 ) ;
 assign wire139 = ( n_n1301 ) | ( wire106 ) | ( wire3390 ) ;
 assign wire3393 = ( wire249 ) | ( wire183 ) | ( wire207 ) | ( wire426 ) ;
 assign wire341 = ( wire237 ) | ( wire139 ) | ( wire3393 ) ;
 assign n_n895 = ( n_n949 ) | ( n_n950 ) | ( n_n1208 ) | ( wire551 ) ;
 assign wire173 = ( wire3221 ) | ( n_n3  &  wire70 ) ;
 assign wire343 = ( wire3222 ) | ( n_n895 ) | ( wire173 ) ;
 assign n_n1181 = ( i_7_  &  i_6_  &  n_n7  &  n_n5 ) ;
 assign n_n716 = ( n_n1083 ) | ( wire236 ) | ( wire473 ) ;
 assign n_n427 = ( wire140 ) | ( n_n716 ) | ( _7869 ) ;
 assign n_n906 = ( (~ i_7_)  &  i_6_  &  n_n0  &  n_n7 ) | ( i_7_  &  (~ i_6_)  &  n_n0  &  n_n7 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n0  &  n_n7 ) ;
 assign n_n1329 = ( (~ i_7_)  &  (~ i_6_)  &  n_n0  &  n_n9 ) ;
 assign n_n459 = ( wire128 ) | ( n_n906 ) | ( n_n1329 ) ;
 assign n_n973 = ( i_7_  &  i_6_  &  n_n6  &  n_n13 ) | ( (~ i_7_)  &  i_6_  &  n_n6  &  n_n13 ) | ( i_7_  &  (~ i_6_)  &  n_n6  &  n_n13 ) ;
 assign n_n1134 = ( i_7_  &  (~ i_6_)  &  n_n6  &  n_n12 ) ;
 assign wire353 = ( i_5_  &  i_3_  &  i_4_  &  _7921 ) ;
 assign n_n904 = ( n_n1121 ) | ( _7923 ) | ( n_n18  &  _7921 ) ;
 assign n_n1037 = ( (~ i_7_)  &  i_6_  &  n_n2  &  n_n11 ) | ( i_7_  &  (~ i_6_)  &  n_n2  &  n_n11 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n2  &  n_n11 ) ;
 assign wire3312 = ( i_7_  &  i_6_  &  n_n2  &  n_n10 ) | ( (~ i_7_)  &  i_6_  &  n_n2  &  n_n10 ) | ( i_7_  &  (~ i_6_)  &  n_n2  &  n_n10 ) ;
 assign n_n996 = ( n_n1037 ) | ( wire3312 ) | ( wire71  &  n_n2 ) ;
 assign n_n1033 = ( (~ i_7_)  &  i_6_  &  n_n2  &  n_n8 ) | ( i_7_  &  (~ i_6_)  &  n_n2  &  n_n8 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n2  &  n_n8 ) ;
 assign wire483 = ( i_7_  &  (~ i_6_)  &  n_n2  &  n_n9 ) ;
 assign wire87 = ( o_7_ ) | ( n_n1268 ) | ( n_n1033 ) | ( wire483 ) ;
 assign wire216 = ( wire249 ) | ( n_n792 ) | ( wire493 ) ;
 assign wire3304 = ( i_7_  &  i_6_  &  n_n0  &  n_n12 ) | ( (~ i_7_)  &  i_6_  &  n_n0  &  n_n12 ) ;
 assign wire3305 = ( i_7_  &  i_6_  &  n_n0  &  n_n13 ) | ( (~ i_7_)  &  i_6_  &  n_n0  &  n_n13 ) | ( i_7_  &  (~ i_6_)  &  n_n0  &  n_n13 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n0  &  n_n13 ) ;
 assign wire3309 = ( n_n1302 ) | ( wire106 ) | ( n_n553 ) ;
 assign wire200 = ( wire216 ) | ( wire3304 ) | ( wire3305 ) | ( wire3309 ) ;
 assign wire67 = ( (~ i_7_)  &  i_6_ ) | ( i_7_  &  (~ i_6_) ) | ( (~ i_7_)  &  (~ i_6_) ) ;
 assign n_n909 = ( i_7_  &  i_6_  &  n_n0  &  n_n9 ) | ( (~ i_7_)  &  i_6_  &  n_n0  &  n_n9 ) | ( i_7_  &  (~ i_6_)  &  n_n0  &  n_n9 ) ;
 assign wire261 = ( n_n909 ) | ( n_n0  &  n_n10  &  wire67 ) ;
 assign n_n1256 = ( (~ i_7_)  &  (~ i_6_)  &  n_n2  &  n_n12 ) ;
 assign n_n1229 = ( i_7_  &  (~ i_6_)  &  n_n3  &  n_n11 ) ;
 assign n_n953 = ( i_7_  &  i_6_  &  n_n4  &  n_n10 ) | ( (~ i_7_)  &  i_6_  &  n_n4  &  n_n10 ) | ( i_7_  &  (~ i_6_)  &  n_n4  &  n_n10 ) ;
 assign wire110 = ( n_n1029 ) | ( n_n1  &  wire70 ) ;
 assign wire177 = ( wire270 ) | ( _8261 ) ;
 assign n_n858 = ( (~ i_7_)  &  i_6_  &  n_n0  &  n_n8 ) | ( i_7_  &  (~ i_6_)  &  n_n0  &  n_n8 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n0  &  n_n8 ) ;
 assign wire3462 = ( wire248 ) | ( n_n0  &  wire71 ) | ( n_n0  &  wire82 ) ;
 assign wire3464 = ( n_n744 ) | ( wire153 ) | ( wire155 ) ;
 assign wire182 = ( n_n858 ) | ( wire3462 ) | ( wire3464 ) ;
 assign wire279 = ( i_7_  &  i_6_  &  n_n7  &  n_n4 ) | ( (~ i_7_)  &  i_6_  &  n_n7  &  n_n4 ) ;
 assign n_n813 = ( i_7_  &  i_6_  &  n_n8  &  n_n4 ) | ( (~ i_7_)  &  i_6_  &  n_n8  &  n_n4 ) | ( i_7_  &  (~ i_6_)  &  n_n8  &  n_n4 ) ;
 assign wire189 = ( o_20_ ) | ( n_n1211 ) | ( wire279 ) | ( n_n813 ) ;
 assign n_n821 = ( i_7_  &  i_6_  &  n_n4  &  n_n18 ) | ( (~ i_7_)  &  i_6_  &  n_n4  &  n_n18 ) | ( i_7_  &  (~ i_6_)  &  n_n4  &  n_n18 ) ;
 assign wire421 = ( (~ i_7_)  &  (~ i_6_)  &  n_n4  &  n_n18 ) ;
 assign wire310 = ( n_n822 ) | ( n_n821 ) | ( wire421 ) ;
 assign wire102 = ( i_7_  &  i_6_  &  n_n12 ) ;
 assign wire84 = ( wire3304 ) | ( wire3305 ) ;
 assign n_n1283 = ( i_7_  &  i_6_  &  n_n12  &  n_n1 ) ;
 assign n_n580 = ( (~ i_7_)  &  i_6_  &  n_n12  &  n_n1 ) | ( i_7_  &  (~ i_6_)  &  n_n12  &  n_n1 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n12  &  n_n1 ) ;
 assign wire260 = ( i_7_  &  (~ i_6_)  &  n_n13  &  n_n1 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n13  &  n_n1 ) ;
 assign wire129 = ( n_n1283 ) | ( n_n580 ) | ( wire260 ) ;
 assign wire153 = ( i_7_  &  i_6_  &  n_n0  &  n_n11 ) | ( (~ i_7_)  &  i_6_  &  n_n0  &  n_n11 ) | ( i_7_  &  (~ i_6_)  &  n_n0  &  n_n11 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n0  &  n_n11 ) ;
 assign wire155 = ( i_7_  &  (~ i_6_)  &  n_n0  &  n_n12 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n0  &  n_n12 ) ;
 assign wire148 = ( n_n554 ) | ( n_n1  &  wire72 ) ;
 assign wire487 = ( i_7_  &  i_6_  &  n_n1  &  n_n10 ) | ( (~ i_7_)  &  i_6_  &  n_n1  &  n_n10 ) ;
 assign wire488 = ( (~ i_7_)  &  (~ i_6_)  &  n_n11  &  n_n1 ) ;
 assign wire3311 = ( i_7_  &  i_6_  &  n_n11  &  n_n1 ) | ( (~ i_7_)  &  i_6_  &  n_n11  &  n_n1 ) | ( i_7_  &  (~ i_6_)  &  n_n11  &  n_n1 ) ;
 assign wire201 = ( n_n554 ) | ( _8180 ) | ( n_n1  &  wire72 ) ;
 assign wire221 = ( n_n996 ) | ( n_n2  &  n_n17  &  n_n11 ) ;
 assign n_n805 = ( i_7_  &  i_6_  &  n_n3  &  n_n10 ) | ( (~ i_7_)  &  i_6_  &  n_n3  &  n_n10 ) | ( i_7_  &  (~ i_6_)  &  n_n3  &  n_n10 ) ;
 assign n_n1238 = ( (~ i_7_)  &  (~ i_6_)  &  n_n3  &  n_n9 ) ;
 assign n_n1239 = ( i_7_  &  i_6_  &  n_n8  &  n_n3 ) ;
 assign wire450 = ( i_7_  &  (~ i_6_)  &  n_n3  &  n_n9 ) ;
 assign n_n803 = ( n_n1238 ) | ( n_n1239 ) | ( wire450 ) ;
 assign wire3465 = ( i_7_  &  i_6_  &  n_n3  &  n_n18 ) | ( (~ i_7_)  &  i_6_  &  n_n3  &  n_n18 ) | ( i_7_  &  (~ i_6_)  &  n_n3  &  n_n18 ) ;
 assign wire3467 = ( o_15_ ) | ( n_n1223 ) | ( wire414 ) ;
 assign wire159 = ( (~ i_7_)  &  i_6_  &  n_n2  &  n_n8 ) | ( i_7_  &  (~ i_6_)  &  n_n2  &  n_n8 ) ;
 assign n_n16 = ( (~ i_7_)  &  i_6_ ) ;
 assign wire164 = ( wire88 ) | ( n_n4  &  n_n11  &  n_n16 ) ;
 assign wire277 = ( i_7_  &  i_6_  &  n_n2  &  n_n18 ) | ( (~ i_7_)  &  i_6_  &  n_n2  &  n_n18 ) ;
 assign wire288 = ( i_7_  &  (~ i_6_)  &  n_n4  &  n_n10 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n4  &  n_n10 ) ;
 assign wire293 = ( n_n4  &  n_n12  &  n_n15 ) | ( n_n4  &  n_n11  &  n_n15 ) ;
 assign n_n1285 = ( i_7_  &  (~ i_6_)  &  n_n12  &  n_n1 ) ;
 assign n_n923 = ( wire243 ) | ( n_n1287 ) | ( n_n1285 ) ;
 assign n_n814 = ( (~ i_7_)  &  i_6_  &  n_n4  &  n_n9 ) | ( i_7_  &  (~ i_6_)  &  n_n4  &  n_n9 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n4  &  n_n9 ) ;
 assign n_n1122 = ( (~ i_7_)  &  i_6_  &  n_n7  &  n_n19 ) ;
 assign n_n1288 = ( (~ i_7_)  &  i_6_  &  n_n11  &  n_n1 ) ;
 assign n_n963 = ( (~ i_1_)  &  i_2_  &  i_0_  &  wire72 ) ;
 assign n_n1006 = ( n_n1137 ) | ( n_n1135 ) | ( wire337 ) ;
 assign n_n1204 = ( i_7_  &  i_6_  &  n_n4  &  n_n9 ) ;
 assign wire86 = ( n_n1211 ) | ( wire279 ) | ( n_n813 ) ;
 assign n_n961 = ( i_7_  &  i_6_  &  n_n5  &  n_n8 ) | ( (~ i_7_)  &  i_6_  &  n_n5  &  n_n8 ) | ( i_7_  &  (~ i_6_)  &  n_n5  &  n_n8 ) ;
 assign wire111 = ( n_n961 ) | ( n_n5  &  n_n9  &  wire67 ) ;
 assign wire130 = ( i_7_  &  i_6_  &  n_n12  &  n_n1 ) | ( (~ i_7_)  &  i_6_  &  n_n12  &  n_n1 ) ;
 assign wire136 = ( n_n6  &  n_n18 ) | ( n_n6  &  wire70 ) ;
 assign n_n1192 = ( (~ i_7_)  &  (~ i_6_)  &  n_n4  &  n_n13 ) ;
 assign wire534 = ( i_7_  &  (~ i_6_)  &  n_n4  &  n_n13 ) ;
 assign wire3535 = ( (~ i_7_)  &  i_6_  &  n_n4  &  n_n12 ) | ( i_7_  &  (~ i_6_)  &  n_n4  &  n_n12 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n4  &  n_n12 ) ;
 assign wire154 = ( o_14_ ) | ( n_n1192 ) | ( wire534 ) | ( wire3535 ) ;
 assign wire253 = ( wire3312 ) | ( wire71  &  n_n2 ) ;
 assign wire274 = ( i_7_  &  i_6_  &  n_n4  &  n_n11 ) | ( (~ i_7_)  &  i_6_  &  n_n4  &  n_n11 ) ;
 assign wire434 = ( (~ i_7_)  &  i_6_  &  n_n3  &  n_n9 ) | ( i_7_  &  (~ i_6_)  &  n_n3  &  n_n9 ) ;
 assign wire276 = ( n_n1238 ) | ( n_n1239 ) | ( wire434 ) ;
 assign wire291 = ( i_7_  &  i_6_  &  n_n4  &  n_n13 ) | ( (~ i_7_)  &  i_6_  &  n_n4  &  n_n13 ) ;
 assign wire305 = ( i_7_  &  i_6_  &  n_n2  &  n_n11 ) | ( (~ i_7_)  &  i_6_  &  n_n2  &  n_n11 ) | ( i_7_  &  (~ i_6_)  &  n_n2  &  n_n11 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n2  &  n_n11 ) ;
 assign n_n934 = ( (~ i_7_)  &  i_6_  &  n_n2  &  n_n12 ) | ( i_7_  &  (~ i_6_)  &  n_n2  &  n_n12 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n2  &  n_n12 ) ;
 assign n_n797 = ( i_7_  &  i_6_  &  n_n2  &  n_n12 ) | ( (~ i_7_)  &  i_6_  &  n_n2  &  n_n12 ) | ( i_7_  &  (~ i_6_)  &  n_n2  &  n_n12 ) ;
 assign wire345 = ( n_n1253 ) | ( n_n934 ) | ( n_n797 ) ;
 assign n_n128 = ( wire94 ) | ( n_n973 ) | ( n_n6  &  n_n18 ) ;
 assign wire242 = ( (~ i_7_)  &  (~ i_6_)  &  n_n4  &  n_n12 ) ;
 assign wire3573 = ( i_7_  &  i_6_  &  n_n4  &  n_n12 ) | ( (~ i_7_)  &  i_6_  &  n_n4  &  n_n12 ) | ( i_7_  &  (~ i_6_)  &  n_n4  &  n_n12 ) ;
 assign n_n1002 = ( n_n1061 ) | ( wire274 ) | ( wire242 ) | ( wire3573 ) ;
 assign wire592 = ( i_7_  &  i_6_  &  n_n4  &  n_n18 ) ;
 assign wire156 = ( wire186 ) | ( n_n958 ) | ( wire592 ) ;
 assign wire193 = ( o_6_ ) | ( wire568 ) | ( wire298 ) | ( wire110 ) ;
 assign n_n1074 = ( (~ i_7_)  &  i_6_  &  n_n8  &  n_n6 ) | ( i_7_  &  (~ i_6_)  &  n_n8  &  n_n6 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n8  &  n_n6 ) ;
 assign n_n609 = ( wire3349 ) | ( n_n5  &  n_n13 ) | ( n_n5  &  wire70 ) ;
 assign wire286 = ( i_7_  &  i_6_  &  n_n5  &  n_n18 ) | ( (~ i_7_)  &  i_6_  &  n_n5  &  n_n18 ) ;
 assign wire316 = ( i_7_  &  i_6_  &  n_n7  &  n_n6 ) | ( (~ i_7_)  &  i_6_  &  n_n7  &  n_n6 ) | ( i_7_  &  (~ i_6_)  &  n_n7  &  n_n6 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n7  &  n_n6 ) ;
 assign wire255 = ( n_n1074 ) | ( n_n609 ) | ( wire286 ) | ( wire316 ) ;
 assign wire3577 = ( n_n19  &  wire163 ) | ( n_n19  &  n_n10  &  wire64 ) ;
 assign wire284 = ( n_n1083 ) | ( wire236 ) | ( wire3577 ) ;
 assign n_n673 = ( o_11_ ) | ( n_n1147 ) | ( wire532 ) ;
 assign wire313 = ( n_n1136 ) | ( n_n1134 ) | ( n_n673 ) ;
 assign n_n1320 = ( i_7_  &  (~ i_6_)  &  n_n0  &  n_n11 ) ;
 assign wire3216 = ( n_n1013 ) | ( n_n0  &  wire72 ) ;
 assign wire332 = ( n_n1017 ) | ( wire76 ) | ( wire3216 ) | ( _7160 ) ;
 assign n_n1010 = ( i_7_  &  (~ i_6_)  &  n_n0  &  n_n7 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n0  &  n_n7 ) ;
 assign n_n1272 = ( i_7_  &  i_6_  &  n_n7  &  n_n2 ) ;
 assign n_n95 = ( n_n930 ) | ( wire132 ) | ( _8519 ) ;
 assign n_n1334 = ( i_7_  &  i_6_  &  n_n0  &  n_n7 ) ;
 assign n_n1314 = ( i_7_  &  i_6_  &  n_n0  &  n_n12 ) ;
 assign n_n1282 = ( (~ i_7_)  &  (~ i_6_)  &  n_n13  &  n_n1 ) ;
 assign n_n925 = ( i_7_  &  i_6_  &  n_n13  &  n_n1 ) | ( (~ i_7_)  &  i_6_  &  n_n13  &  n_n1 ) | ( i_7_  &  (~ i_6_)  &  n_n13  &  n_n1 ) ;
 assign n_n1013 = ( (~ i_7_)  &  i_6_  &  n_n0  &  n_n9 ) | ( i_7_  &  (~ i_6_)  &  n_n0  &  n_n9 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n0  &  n_n9 ) ;
 assign n_n990 = ( wire128 ) | ( n_n1013 ) | ( _8530 ) ;
 assign wire3621 = ( wire71  &  n_n1 ) | ( n_n11  &  n_n1  &  n_n16 ) ;
 assign wire179 = ( o_6_ ) | ( n_n921 ) | ( n_n923 ) | ( wire3621 ) ;
 assign wire174 = ( i_7_  &  i_6_  &  n_n0  &  n_n12 ) | ( (~ i_7_)  &  i_6_  &  n_n0  &  n_n12 ) | ( i_7_  &  (~ i_6_)  &  n_n0  &  n_n12 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n0  &  n_n12 ) ;
 assign wire3395 = ( (~ i_7_)  &  i_6_  &  n_n0  &  n_n13 ) | ( i_7_  &  (~ i_6_)  &  n_n0  &  n_n13 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n0  &  n_n13 ) ;
 assign wire283 = ( wire3358 ) | ( _7830 ) ;
 assign wire3359 = ( n_n805 ) | ( wire135 ) ;
 assign wire238 = ( n_n803 ) | ( _7839 ) | ( wire71  &  _7818 ) ;
 assign n_n1300 = ( (~ i_7_)  &  i_6_  &  n_n8  &  n_n1 ) ;
 assign wire3638 = ( i_7_  &  i_6_  &  n_n3  &  n_n18 ) | ( (~ i_7_)  &  i_6_  &  n_n3  &  n_n18 ) | ( i_7_  &  (~ i_6_)  &  n_n3  &  n_n18 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n3  &  n_n18 ) ;
 assign n_n490 = ( wire189 ) | ( wire97 ) | ( _8569 ) | ( _9005 ) ;
 assign n_n1231 = ( i_7_  &  i_6_  &  n_n3  &  n_n10 ) ;
 assign wire135 = ( i_7_  &  (~ i_6_)  &  n_n3  &  n_n11 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n3  &  n_n11 ) ;
 assign wire545 = ( (~ i_7_)  &  i_6_  &  n_n3  &  n_n10 ) | ( i_7_  &  (~ i_6_)  &  n_n3  &  n_n10 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n3  &  n_n10 ) ;
 assign wire546 = ( i_7_  &  i_6_  &  n_n3  &  n_n9 ) | ( (~ i_7_)  &  i_6_  &  n_n3  &  n_n9 ) | ( i_7_  &  (~ i_6_)  &  n_n3  &  n_n9 ) ;
 assign n_n1258 = ( (~ i_7_)  &  i_6_  &  n_n2  &  n_n11 ) ;
 assign n_n1275 = ( i_7_  &  i_6_  &  n_n1  &  n_n18 ) ;
 assign n_n534 = ( wire254 ) | ( wire132 ) | ( n_n1275 ) ;
 assign n_n926 = ( (~ i_7_)  &  i_6_  &  n_n1  &  n_n18 ) | ( i_7_  &  (~ i_6_)  &  n_n1  &  n_n18 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n1  &  n_n18 ) ;
 assign wire266 = ( i_7_  &  (~ i_6_)  &  n_n0  &  n_n13 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n0  &  n_n13 ) ;
 assign n_n1018 = ( wire266 ) | ( n_n0  &  n_n17  &  n_n12 ) ;
 assign n_n1301 = ( i_7_  &  (~ i_6_)  &  n_n8  &  n_n1 ) ;
 assign wire64 = ( i_7_  &  i_6_ ) | ( (~ i_7_)  &  i_6_ ) | ( i_7_  &  (~ i_6_) ) ;
 assign wire83 = ( n_n1021 ) | ( n_n0  &  n_n18  &  wire64 ) ;
 assign wire183 = ( i_7_  &  (~ i_6_)  &  n_n1  &  n_n9 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n1  &  n_n9 ) ;
 assign wire109 = ( (~ i_7_)  &  i_6_  &  n_n8  &  n_n3 ) | ( i_7_  &  (~ i_6_)  &  n_n8  &  n_n3 ) ;
 assign wire112 = ( i_7_  &  i_6_  &  n_n7  &  n_n3 ) | ( (~ i_7_)  &  i_6_  &  n_n7  &  n_n3 ) ;
 assign wire247 = ( n_n3  &  n_n13  &  n_n14 ) | ( n_n3  &  n_n9  &  n_n14 ) ;
 assign wire257 = ( i_7_  &  i_6_  &  n_n2  &  n_n12 ) | ( (~ i_7_)  &  i_6_  &  n_n2  &  n_n12 ) | ( i_7_  &  (~ i_6_)  &  n_n2  &  n_n12 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n2  &  n_n12 ) ;
 assign n_n1254 = ( (~ i_7_)  &  i_6_  &  n_n2  &  n_n12 ) ;
 assign n_n1330 = ( i_7_  &  i_6_  &  n_n0  &  n_n8 ) ;
 assign wire268 = ( i_7_  &  i_6_  &  n_n2  &  n_n18 ) | ( (~ i_7_)  &  i_6_  &  n_n2  &  n_n18 ) | ( i_7_  &  (~ i_6_)  &  n_n2  &  n_n18 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n2  &  n_n18 ) ;
 assign n_n1040 = ( i_7_  &  i_6_  &  n_n2  &  n_n13 ) | ( (~ i_7_)  &  i_6_  &  n_n2  &  n_n13 ) | ( i_7_  &  (~ i_6_)  &  n_n2  &  n_n13 ) ;
 assign n_n642 = ( wire146 ) | ( wire268 ) | ( n_n1040 ) ;
 assign n_n574 = ( wire147 ) | ( n_n1261 ) | ( n_n616 ) | ( n_n617 ) ;
 assign wire3671 = ( n_n859 ) | ( wire297 ) | ( n_n963 ) | ( wire3279 ) ;
 assign wire3672 = ( wire113 ) | ( _8626 ) | ( wire71  &  n_n19 ) ;
 assign wire3674 = ( n_n128 ) | ( wire3283 ) | ( wire3282 ) | ( wire3667 ) ;
 assign wire3676 = ( wire152 ) | ( n_n673 ) | ( wire3668 ) | ( wire3669 ) ;
 assign wire259 = ( (~ i_7_)  &  i_6_  &  n_n0  &  n_n8 ) | ( i_7_  &  (~ i_6_)  &  n_n0  &  n_n8 ) ;
 assign n_n660 = ( wire306 ) | ( wire237 ) | ( wire139 ) | ( wire3393 ) ;
 assign n_n1147 = ( (~ i_7_)  &  (~ i_6_)  &  n_n6  &  n_n9 ) ;
 assign wire532 = ( n_n6  &  n_n10 ) | ( n_n6  &  n_n9  &  wire64 ) ;
 assign wire78 = ( (~ i_7_)  &  i_6_  &  n_n5  &  n_n11 ) | ( i_7_  &  (~ i_6_)  &  n_n5  &  n_n11 ) ;
 assign wire99 = ( o_28_ ) | ( n_n1166 ) | ( wire78 ) ;
 assign wire500 = ( (~ i_7_)  &  (~ i_6_)  &  n_n4  &  n_n18 ) ;
 assign n_n1170 = ( i_7_  &  i_6_  &  n_n5  &  n_n10 ) ;
 assign wire235 = ( n_n1169 ) | ( n_n826 ) | ( n_n1170 ) ;
 assign wire97 = ( n_n1204 ) | ( wire413 ) | ( _8561 ) ;
 assign n_n817 = ( i_7_  &  i_6_  &  n_n4  &  n_n11 ) | ( (~ i_7_)  &  i_6_  &  n_n4  &  n_n11 ) | ( i_7_  &  (~ i_6_)  &  n_n4  &  n_n11 ) ;
 assign wire315 = ( n_n814 ) | ( wire154 ) | ( wire97 ) | ( n_n817 ) ;
 assign n_n802 = ( (~ i_7_)  &  i_6_  &  n_n8  &  n_n3 ) | ( i_7_  &  (~ i_6_)  &  n_n8  &  n_n3 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n8  &  n_n3 ) ;
 assign wire325 = ( o_10_ ) | ( wire112 ) | ( n_n802 ) ;
 assign wire281 = ( i_7_  &  i_6_  &  n_n1  &  n_n18 ) | ( (~ i_7_)  &  i_6_  &  n_n1  &  n_n18 ) ;
 assign n_n1032 = ( i_7_  &  i_6_  &  n_n7  &  n_n2 ) | ( (~ i_7_)  &  i_6_  &  n_n7  &  n_n2 ) | ( i_7_  &  (~ i_6_)  &  n_n7  &  n_n2 ) ;
 assign wire165 = ( n_n1274 ) | ( wire87 ) | ( wire281 ) | ( n_n1032 ) ;
 assign n_n1257 = ( i_7_  &  i_6_  &  n_n2  &  n_n11 ) ;
 assign n_n745 = ( (~ i_7_)  &  i_6_  &  n_n0  &  n_n11 ) | ( i_7_  &  (~ i_6_)  &  n_n0  &  n_n11 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n0  &  n_n11 ) ;
 assign wire181 = ( wire3387 ) | ( wire3388 ) | ( wire112 ) | ( _8108 ) ;
 assign n_n1227 = ( i_7_  &  i_6_  &  n_n3  &  n_n11 ) ;
 assign wire3358 = ( i_7_  &  (~ i_6_)  &  n_n3  &  n_n12 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n3  &  n_n12 ) ;
 assign wire292 = ( i_7_  &  i_6_  &  n_n3  &  n_n10 ) | ( (~ i_7_)  &  i_6_  &  n_n3  &  n_n10 ) ;
 assign n_n1216 = ( i_7_  &  i_6_  &  n_n3  &  n_n18 ) ;
 assign n_n1244 = ( i_7_  &  (~ i_6_)  &  n_n7  &  n_n3 ) ;
 assign n_n554 = ( (~ i_7_)  &  i_6_  &  n_n1  &  n_n9 ) | ( i_7_  &  (~ i_6_)  &  n_n1  &  n_n9 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n1  &  n_n9 ) ;
 assign n_n810 = ( (~ i_7_)  &  i_6_  &  n_n3  &  n_n18 ) | ( i_7_  &  (~ i_6_)  &  n_n3  &  n_n18 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n3  &  n_n18 ) ;
 assign n_n1269 = ( (~ i_7_)  &  i_6_  &  n_n2  &  n_n8 ) ;
 assign wire150 = ( wire487 ) | ( wire488 ) | ( wire3311 ) ;
 assign wire308 = ( (~ i_7_)  &  i_6_  &  n_n6  &  n_n11 ) | ( i_7_  &  (~ i_6_)  &  n_n6  &  n_n11 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n6  &  n_n11 ) ;
 assign wire340 = ( wire138 ) | ( n_n574 ) | ( n_n2  &  wire70 ) ;
 assign wire191 = ( wire564 ) | ( _7076 ) ;
 assign wire342 = ( wire187 ) | ( wire99 ) | ( wire564 ) | ( _7076 ) ;
 assign n_n1224 = ( (~ i_7_)  &  i_6_  &  n_n3  &  n_n12 ) ;
 assign n_n937 = ( i_7_  &  i_6_  &  n_n2  &  n_n18 ) | ( (~ i_7_)  &  i_6_  &  n_n2  &  n_n18 ) | ( i_7_  &  (~ i_6_)  &  n_n2  &  n_n18 ) ;
 assign wire3802 = ( (~ i_7_)  &  i_6_  &  n_n7  &  n_n3 ) | ( i_7_  &  (~ i_6_)  &  n_n7  &  n_n3 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n7  &  n_n3 ) ;
 assign n_n711 = ( n_n937 ) | ( wire3802 ) | ( n_n2  &  wire69 ) ;
 assign n_n1284 = ( (~ i_7_)  &  i_6_  &  n_n12  &  n_n1 ) ;
 assign wire95 = ( wire3465 ) | ( n_n3  &  wire69 ) ;
 assign wire3384 = ( i_7_  &  i_6_  &  n_n1  &  n_n18 ) | ( (~ i_7_)  &  i_6_  &  n_n1  &  n_n18 ) | ( i_7_  &  (~ i_6_)  &  n_n1  &  n_n18 ) ;
 assign wire107 = ( wire3384 ) | ( n_n1  &  wire69 ) ;
 assign n_n1243 = ( i_7_  &  i_6_  &  n_n7  &  n_n3 ) ;
 assign wire217 = ( wire246 ) | ( wire109 ) | ( n_n1243 ) ;
 assign wire231 = ( wire132 ) | ( n_n7  &  n_n2  &  n_n16 ) ;
 assign wire295 = ( o_13_ ) | ( n_n1253 ) | ( wire588 ) | ( n_n934 ) ;
 assign wire3485 = ( o_20_ ) | ( n_n8  &  n_n4  &  n_n15 ) ;
 assign wire3486 = ( n_n1211 ) | ( wire279 ) | ( wire512 ) | ( wire3294 ) ;
 assign wire3804 = ( o_21_ ) | ( n_n1203 ) | ( n_n1056 ) | ( n_n953 ) ;
 assign n_n1034 = ( o_7_ ) | ( n_n1268 ) | ( wire483 ) ;
 assign wire504 = ( (~ i_7_)  &  (~ i_6_)  &  n_n5  &  n_n9 ) ;
 assign wire505 = ( (~ i_7_)  &  i_6_  &  n_n5  &  n_n8 ) ;
 assign n_n824 = ( o_12_ ) | ( wire504 ) | ( wire505 ) ;
 assign wire412 = ( i_7_  &  i_6_  &  n_n4  &  n_n10 ) | ( (~ i_7_)  &  i_6_  &  n_n4  &  n_n10 ) ;
 assign wire413 = ( (~ i_7_)  &  (~ i_6_)  &  n_n4  &  n_n11 ) ;
 assign wire101 = ( i_7_  &  (~ i_6_)  &  n_n8 ) ;
 assign wire271 = ( i_7_  &  i_6_  &  n_n7  &  n_n5 ) | ( (~ i_7_)  &  i_6_  &  n_n7  &  n_n5 ) ;
 assign wire320 = ( wire180 ) | ( wire186 ) | ( n_n958 ) | ( wire592 ) ;
 assign n_n1165 = ( i_7_  &  (~ i_6_)  &  n_n5  &  n_n12 ) ;
 assign n_n989 = ( n_n1008 ) | ( wire136 ) | ( _8910 ) ;
 assign n_n1322 = ( i_7_  &  i_6_  &  n_n0  &  n_n10 ) ;
 assign wire106 = ( i_7_  &  i_6_  &  n_n7  &  n_n1 ) | ( (~ i_7_)  &  i_6_  &  n_n7  &  n_n1 ) ;
 assign wire3390 = ( (~ i_7_)  &  i_6_  &  n_n8  &  n_n1 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n8  &  n_n1 ) ;
 assign wire207 = ( i_7_  &  i_6_  &  n_n8  &  n_n1 ) ;
 assign n_n1139 = ( (~ i_7_)  &  (~ i_6_)  &  n_n6  &  n_n11 ) ;
 assign n_n553 = ( i_7_  &  i_6_  &  n_n8  &  n_n1 ) | ( (~ i_7_)  &  i_6_  &  n_n8  &  n_n1 ) | ( i_7_  &  (~ i_6_)  &  n_n8  &  n_n1 ) ;
 assign n_n1138 = ( i_7_  &  (~ i_6_)  &  n_n6  &  n_n11 ) ;
 assign wire113 = ( (~ i_7_)  &  i_6_  &  n_n8  &  n_n19 ) | ( i_7_  &  (~ i_6_)  &  n_n8  &  n_n19 ) ;
 assign wire158 = ( (~ i_7_)  &  i_6_  &  n_n8  &  n_n6 ) | ( i_7_  &  (~ i_6_)  &  n_n8  &  n_n6 ) ;
 assign wire161 = ( i_7_  &  i_6_  &  n_n19  &  n_n11 ) | ( (~ i_7_)  &  i_6_  &  n_n19  &  n_n11 ) ;
 assign n_n962 = ( (~ i_7_)  &  i_6_  &  n_n5  &  n_n9 ) | ( i_7_  &  (~ i_6_)  &  n_n5  &  n_n9 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n5  &  n_n9 ) ;
 assign n_n799 = ( i_1_  &  (~ i_2_)  &  (~ i_0_)  &  wire70 ) ;
 assign wire3973 = ( n_n1268 ) | ( wire132 ) | ( n_n1272 ) ;
 assign wire3978 = ( wire270 ) | ( wire238 ) | ( _8261 ) | ( _9011 ) ;
 assign wire265 = ( i_7_  &  i_6_  &  n_n0  &  n_n10 ) | ( (~ i_7_)  &  i_6_  &  n_n0  &  n_n10 ) ;
 assign n_n1155 = ( i_7_  &  i_6_  &  n_n5  &  n_n18 ) ;
 assign wire466 = ( n_n6  &  n_n10 ) | ( n_n6  &  n_n9  &  wire64 ) ;
 assign n_n738 = ( wire93 ) | ( wire466 ) ;
 assign wire3273 = ( i_7_  &  i_6_  &  n_n7  &  n_n19 ) | ( (~ i_7_)  &  i_6_  &  n_n7  &  n_n19 ) | ( i_7_  &  (~ i_6_)  &  n_n7  &  n_n19 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n7  &  n_n19 ) ;
 assign wire473 = ( i_7_  &  i_6_  &  n_n19  &  n_n10 ) | ( (~ i_7_)  &  i_6_  &  n_n19  &  n_n10 ) ;
 assign wire471 = ( i_7_  &  (~ i_6_)  &  n_n19  &  n_n10 ) ;
 assign wire160 = ( i_7_  &  i_6_  &  n_n7  &  n_n6 ) | ( (~ i_7_)  &  i_6_  &  n_n7  &  n_n6 ) ;
 assign wire323 = ( wire354 ) | ( wire92 ) | ( wire158 ) | ( wire160 ) ;
 assign wire561 = ( (~ i_7_)  &  i_6_  &  n_n3  &  n_n18 ) ;
 assign n_n948 = ( n_n1215 ) | ( n_n1216 ) | ( wire561 ) ;
 assign n_n1167 = ( (~ i_7_)  &  i_6_  &  n_n5  &  n_n11 ) ;
 assign wire461 = ( i_7_  &  i_6_  &  wire93 ) | ( (~ i_7_)  &  i_6_  &  wire93 ) | ( i_7_  &  i_6_  &  wire466 ) | ( (~ i_7_)  &  i_6_  &  wire466 ) ;
 assign wire3341 = ( n_n1136 ) | ( n_n1135 ) | ( n_n1134 ) ;
 assign wire3342 = ( n_n973 ) | ( wire468 ) | ( wire3340 ) ;
 assign wire3348 = ( n_n1147 ) | ( wire160 ) | ( n_n1153 ) | ( wire456 ) ;
 assign n_n901 = ( wire222 ) | ( wire3348 ) ;
 assign n_n582 = ( (~ i_7_)  &  i_6_  &  n_n7  &  n_n2 ) | ( i_7_  &  (~ i_6_)  &  n_n7  &  n_n2 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n7  &  n_n2 ) ;
 assign n_n1148 = ( (~ i_7_)  &  i_6_  &  n_n8  &  n_n6 ) ;
 assign n_n1104 = ( (~ i_7_)  &  i_6_  &  n_n19  &  n_n12 ) ;
 assign n_n1119 = ( (~ i_7_)  &  i_6_  &  n_n8  &  n_n19 ) ;
 assign n_n1303 = ( (~ i_7_)  &  i_6_  &  n_n7  &  n_n1 ) ;
 assign n_n1023 = ( wire3218 ) | ( n_n1  &  n_n9  &  n_n14 ) ;
 assign n_n786 = ( n_n1147 ) | ( wire532 ) | ( n_n1139 ) ;
 assign n_n1273 = ( i_7_  &  (~ i_6_)  &  n_n7  &  n_n2 ) ;
 assign n_n1319 = ( (~ i_7_)  &  i_6_  &  n_n0  &  n_n11 ) ;
 assign n_n825 = ( i_7_  &  i_6_  &  n_n5  &  n_n9 ) | ( (~ i_7_)  &  i_6_  &  n_n5  &  n_n9 ) | ( i_7_  &  (~ i_6_)  &  n_n5  &  n_n9 ) ;
 assign wire549 = ( (~ i_7_)  &  i_6_  &  n_n5  &  n_n10 ) ;
 assign wire273 = ( i_7_  &  i_6_  &  n_n4  &  n_n9 ) | ( (~ i_7_)  &  i_6_  &  n_n4  &  n_n9 ) ;
 assign n_n1153 = ( i_7_  &  (~ i_6_)  &  n_n7  &  n_n6 ) ;
 assign n_n1230 = ( (~ i_7_)  &  (~ i_6_)  &  n_n3  &  n_n11 ) ;
 assign wire507 = ( i_7_  &  (~ i_6_)  &  n_n5  &  n_n8 ) ;
 assign wire3349 = ( i_7_  &  i_6_  &  n_n5  &  n_n12 ) | ( (~ i_7_)  &  i_6_  &  n_n5  &  n_n12 ) | ( i_7_  &  (~ i_6_)  &  n_n5  &  n_n12 ) ;
 assign n_n1315 = ( (~ i_7_)  &  i_6_  &  n_n0  &  n_n12 ) ;
 assign n_n931 = ( i_1_  &  (~ i_2_)  &  (~ i_0_)  &  wire72 ) ;
 assign n_n910 = ( (~ i_7_)  &  i_6_  &  n_n0  &  n_n10 ) | ( i_7_  &  (~ i_6_)  &  n_n0  &  n_n10 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n0  &  n_n10 ) ;
 assign n_n792 = ( (~ i_7_)  &  i_6_  &  n_n0  &  n_n18 ) | ( i_7_  &  (~ i_6_)  &  n_n0  &  n_n18 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n0  &  n_n18 ) ;
 assign wire515 = ( i_7_  &  (~ i_6_)  &  n_n19  &  n_n12 ) ;
 assign wire3283 = ( wire236 ) | ( n_n756 ) | ( n_n1104 ) ;
 assign n_n1213 = ( (~ i_7_)  &  i_6_  &  n_n7  &  n_n4 ) ;
 assign wire219 = ( (~ i_7_)  &  i_6_  &  n_n12  &  n_n1 ) | ( i_7_  &  (~ i_6_)  &  n_n12  &  n_n1 ) ;
 assign wire303 = ( _175 ) | ( n_n1  &  n_n10  &  _7275 ) ;
 assign wire564 = ( i_7_  &  (~ i_6_)  &  n_n5  &  n_n13 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n5  &  n_n13 ) ;
 assign wire133 = ( i_7_  &  (~ i_6_)  &  n_n19  &  n_n9 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n19  &  n_n9 ) ;
 assign wire3363 = ( (~ i_7_)  &  i_6_  &  n_n2  &  n_n13 ) | ( i_7_  &  (~ i_6_)  &  n_n2  &  n_n13 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n2  &  n_n13 ) ;
 assign wire493 = ( i_7_  &  i_6_  &  n_n0  &  n_n18 ) ;
 assign wire414 = ( i_7_  &  (~ i_6_)  &  n_n3  &  n_n13 ) ;
 assign wire426 = ( i_7_  &  i_6_  &  n_n0  &  n_n18 ) | ( (~ i_7_)  &  i_6_  &  n_n0  &  n_n18 ) ;
 assign wire456 = ( i_7_  &  (~ i_6_)  &  n_n6  &  n_n9 ) ;
 assign wire462 = ( n_n10  &  wire93 ) | ( n_n10  &  wire466 ) ;
 assign wire468 = ( (~ i_7_)  &  (~ i_6_)  &  n_n6  &  n_n13 ) ;
 assign wire512 = ( (~ i_7_)  &  (~ i_6_)  &  n_n4  &  n_n9 ) ;
 assign wire3176 = ( (~ i_5_)  &  i_3_  &  i_4_  &  n_n14 ) | ( (~ i_5_)  &  (~ i_3_)  &  i_4_  &  n_n14 ) ;
 assign wire3177 = ( n_n11  &  n_n14 ) | ( n_n7  &  n_n5  &  n_n14 ) ;
 assign wire3178 = ( n_n7  &  n_n6  &  n_n14 ) | ( n_n7  &  n_n3  &  n_n14 ) ;
 assign wire3195 = ( i_7_  &  (~ i_6_)  &  n_n11 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n11 ) ;
 assign wire3196 = ( n_n4  &  n_n11  &  wire66 ) | ( n_n11  &  n_n1  &  wire66 ) ;
 assign wire3203 = ( n_n1168 ) | ( n_n1321 ) | ( wire3196 ) ;
 assign wire3206 = ( wire94 ) | ( wire146 ) | ( wire147 ) | ( wire186 ) ;
 assign wire3236 = ( (~ i_7_)  &  i_6_  &  n_n7  &  n_n3 ) | ( i_7_  &  (~ i_6_)  &  n_n7  &  n_n3 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n7  &  n_n3 ) ;
 assign wire3245 = ( o_7_ ) | ( wire186 ) | ( n_n1120 ) | ( wire592 ) ;
 assign wire3248 = ( wire93 ) | ( n_n872 ) | ( wire159 ) | ( wire219 ) ;
 assign wire3250 = ( n_n1083 ) | ( wire236 ) | ( wire3213 ) | ( _7043 ) ;
 assign wire3251 = ( wire354 ) | ( wire92 ) | ( wire222 ) | ( wire160 ) ;
 assign wire3256 = ( wire187 ) | ( wire226 ) | ( wire3248 ) ;
 assign wire3257 = ( wire295 ) | ( _7324 ) | ( _7325 ) | ( _7326 ) ;
 assign wire3261 = ( wire228 ) | ( wire99 ) | ( wire191 ) | ( wire3251 ) ;
 assign wire3262 = ( wire280 ) | ( wire327 ) | ( wire331 ) | ( wire346 ) ;
 assign wire3264 = ( wire301 ) | ( n_n387 ) | ( wire3237 ) | ( wire3238 ) ;
 assign wire3277 = ( _583 ) | ( n_n8  &  n_n6  &  _7486 ) ;
 assign wire3278 = ( n_n5  &  n_n12  &  n_n16 ) | ( n_n5  &  n_n18  &  n_n16 ) ;
 assign wire3279 = ( n_n1163 ) | ( wire564 ) | ( wire3278 ) ;
 assign wire3282 = ( n_n1009 ) | ( n_n19  &  n_n12  &  n_n15 ) ;
 assign wire3285 = ( (~ i_7_)  &  i_6_  &  n_n6  &  n_n11 ) | ( i_7_  &  (~ i_6_)  &  n_n6  &  n_n11 ) ;
 assign wire3286 = ( o_28_ ) | ( wire78 ) | ( n_n1165 ) ;
 assign wire3287 = ( n_n1169 ) | ( n_n826 ) | ( n_n1170 ) | ( wire3285 ) ;
 assign wire3294 = ( i_7_  &  i_6_  &  n_n8  &  n_n4 ) | ( (~ i_7_)  &  i_6_  &  n_n8  &  n_n4 ) ;
 assign wire3313 = ( n_n4  &  n_n10 ) | ( n_n4  &  n_n11  &  wire66 ) ;
 assign wire3316 = ( n_n8  &  n_n4  &  n_n15 ) | ( n_n4  &  n_n12  &  n_n15 ) ;
 assign wire3317 = ( o_20_ ) | ( n_n2  &  wire69 ) ;
 assign wire3318 = ( n_n1029 ) | ( n_n1  &  wire70 ) ;
 assign wire3319 = ( wire184 ) | ( wire3313 ) ;
 assign wire3320 = ( n_n1211 ) | ( n_n1197 ) | ( n_n1193 ) | ( n_n1225 ) ;
 assign wire3321 = ( o_14_ ) | ( n_n1192 ) | ( wire534 ) | ( wire3316 ) ;
 assign wire3322 = ( n_n1028 ) | ( wire512 ) | ( wire3294 ) ;
 assign wire3327 = ( wire77 ) | ( n_n935 ) | ( n_n1213 ) | ( wire3322 ) ;
 assign wire3328 = ( wire3317 ) | ( wire3318 ) | ( wire3319 ) | ( wire3320 ) ;
 assign wire3329 = ( wire218 ) | ( n_n1056 ) | ( wire3321 ) | ( _7583 ) ;
 assign wire3340 = ( i_7_  &  i_6_  &  n_n6  &  n_n12 ) | ( (~ i_7_)  &  i_6_  &  n_n6  &  n_n12 ) ;
 assign wire3350 = ( n_n1154 ) | ( n_n1169 ) | ( n_n1170 ) ;
 assign wire3351 = ( o_28_ ) | ( n_n1166 ) | ( wire286 ) | ( wire78 ) ;
 assign wire3353 = ( wire222 ) | ( wire3348 ) | ( wire3351 ) ;
 assign wire3367 = ( n_n1194 ) | ( n_n1261 ) | ( n_n1320 ) | ( n_n1010 ) ;
 assign wire3368 = ( wire147 ) | ( n_n616 ) | ( wire274 ) | ( wire242 ) ;
 assign wire3370 = ( n_n602 ) | ( n_n1022 ) | ( n_n1298 ) | ( wire3218 ) ;
 assign wire3373 = ( wire85 ) | ( n_n1021 ) | ( _473 ) | ( _7801 ) ;
 assign wire3375 = ( wire114 ) | ( wire298 ) | ( wire3367 ) | ( wire3368 ) ;
 assign wire3383 = ( _363 ) | ( n_n2  &  n_n11  &  _8137 ) ;
 assign wire3400 = ( i_7_  &  i_6_  &  n_n19  &  n_n11 ) | ( i_7_  &  (~ i_6_)  &  n_n19  &  n_n11 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n19  &  n_n11 ) ;
 assign wire3404 = ( n_n921 ) | ( wire71  &  n_n1 ) | ( n_n1  &  wire3195 ) ;
 assign wire3405 = ( o_21_ ) | ( n_n1168 ) | ( n_n1196 ) | ( n_n953 ) ;
 assign wire3406 = ( n_n1287 ) | ( n_n1163 ) | ( n_n1318 ) | ( n_n1189 ) ;
 assign wire3407 = ( n_n1203 ) | ( n_n756 ) | ( n_n1135 ) | ( wire273 ) ;
 assign wire3408 = ( n_n1049 ) | ( n_n1227 ) | ( wire3358 ) ;
 assign wire3410 = ( wire93 ) | ( wire186 ) | ( wire3400 ) ;
 assign wire3411 = ( n_n1083 ) | ( n_n1009 ) | ( n_n864 ) | ( n_n1061 ) ;
 assign wire3414 = ( wire297 ) | ( wire309 ) | ( wire3408 ) ;
 assign wire3420 = ( wire345 ) | ( wire3383 ) | ( wire3410 ) | ( wire3411 ) ;
 assign wire3422 = ( wire324 ) | ( wire343 ) | ( wire3404 ) | ( wire3405 ) ;
 assign wire3432 = ( wire77 ) | ( n_n1231 ) | ( wire135 ) | ( _7056 ) ;
 assign wire3433 = ( n_n1169 ) | ( n_n1147 ) | ( _8193 ) ;
 assign wire3434 = ( wire354 ) | ( wire92 ) | ( wire222 ) | ( wire160 ) ;
 assign wire3436 = ( wire187 ) | ( wire99 ) | ( wire191 ) | ( wire3434 ) ;
 assign wire3437 = ( wire88 ) | ( n_n5  &  wire72 ) ;
 assign wire3439 = ( wire194 ) | ( _8200 ) ;
 assign wire3440 = ( n_n955 ) | ( wire320 ) | ( wire3437 ) ;
 assign wire3441 = ( wire155 ) | ( n_n0  &  n_n11  &  n_n16 ) ;
 assign wire3442 = ( n_n1137 ) | ( n_n1135 ) | ( n_n1134 ) ;
 assign wire3443 = ( n_n973 ) | ( wire468 ) | ( wire3340 ) ;
 assign wire3447 = ( n_n936 ) | ( wire261 ) | ( wire295 ) | ( wire3442 ) ;
 assign wire3460 = ( wire292 ) | ( n_n1230 ) | ( _8258 ) ;
 assign wire3470 = ( i_7_  &  i_6_  &  n_n4  &  n_n10 ) | ( (~ i_7_)  &  i_6_  &  n_n4  &  n_n10 ) | ( i_7_  &  (~ i_6_)  &  n_n4  &  n_n10 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n4  &  n_n10 ) ;
 assign wire3471 = ( o_21_ ) | ( n_n1229 ) | ( _8241 ) ;
 assign wire3472 = ( n_n1029 ) | ( wire3470 ) | ( n_n1  &  wire70 ) ;
 assign wire3475 = ( n_n602 ) | ( n_n1022 ) | ( n_n1023 ) | ( wire3472 ) ;
 assign wire3477 = ( wire298 ) | ( wire216 ) | ( wire84 ) | ( wire3471 ) ;
 assign wire3487 = ( n_n13 ) | ( n_n7  &  n_n2  &  n_n14 ) ;
 assign wire3488 = ( i_7_  &  (~ i_6_)  &  n_n2  &  n_n12 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n2  &  n_n12 ) ;
 assign wire3491 = ( n_n1056 ) | ( n_n1229 ) | ( wire3488 ) ;
 assign wire3493 = ( n_n1283 ) | ( n_n580 ) | ( wire260 ) | ( wire153 ) ;
 assign wire3494 = ( n_n955 ) | ( wire3225 ) | ( wire164 ) | ( wire3491 ) ;
 assign wire3495 = ( o_20_ ) | ( wire3486 ) | ( _302 ) | ( _8309 ) ;
 assign wire3496 = ( wire87 ) | ( wire216 ) | ( wire3309 ) | ( n_n1032 ) ;
 assign wire3497 = ( n_n996 ) | ( wire150 ) | ( _8315 ) ;
 assign wire3498 = ( wire3305 ) | ( wire3487 ) | ( wire3493 ) | ( _8318 ) ;
 assign wire3505 = ( n_n2  &  n_n8  &  n_n17 ) | ( n_n8  &  n_n17  &  n_n4 ) ;
 assign wire3506 = ( n_n805 ) | ( wire71  &  n_n3 ) ;
 assign wire3507 = ( wire104 ) | ( wire412 ) | ( wire413 ) ;
 assign wire3510 = ( o_20_ ) | ( wire135 ) | ( wire3505 ) ;
 assign wire3511 = ( n_n930 ) | ( n_n1028 ) | ( n_n2  &  wire72 ) ;
 assign wire3515 = ( wire162 ) | ( wire159 ) | ( wire288 ) | ( wire293 ) ;
 assign wire3516 = ( wire331 ) | ( n_n797 ) | ( wire3363 ) ;
 assign wire3517 = ( wire3467 ) | ( wire95 ) | ( wire3510 ) ;
 assign wire3518 = ( wire77 ) | ( n_n950 ) | ( n_n1213 ) | ( wire3511 ) ;
 assign wire3519 = ( n_n803 ) | ( wire164 ) | ( wire3506 ) | ( wire3507 ) ;
 assign wire3520 = ( n_n602 ) | ( n_n1022 ) | ( n_n1023 ) | ( wire3515 ) ;
 assign wire3533 = ( wire77 ) | ( n_n3  &  wire72 ) ;
 assign wire3541 = ( wire94 ) | ( wire71  &  n_n1 ) ;
 assign wire3542 = ( o_6_ ) | ( n_n921 ) | ( n_n5  &  wire72 ) ;
 assign wire3545 = ( n_n1274 ) | ( n_n1121 ) | ( n_n1180 ) | ( n_n1321 ) ;
 assign wire3546 = ( n_n814 ) | ( n_n1122 ) | ( n_n1288 ) | ( n_n1204 ) ;
 assign wire3548 = ( wire243 ) | ( n_n822 ) | ( n_n1287 ) | ( n_n1285 ) ;
 assign wire3552 = ( wire76 ) | ( wire130 ) | ( wire274 ) | ( wire291 ) ;
 assign wire3554 = ( wire3467 ) | ( wire86 ) | ( wire95 ) ;
 assign wire3557 = ( wire111 ) | ( wire136 ) | ( wire253 ) | ( wire276 ) ;
 assign wire3558 = ( wire3541 ) | ( wire3542 ) | ( wire3552 ) ;
 assign wire3561 = ( wire345 ) | ( wire112 ) | ( n_n642 ) | ( _8108 ) ;
 assign wire3579 = ( wire133 ) | ( n_n8  &  n_n19  &  n_n14 ) ;
 assign wire3582 = ( n_n961 ) | ( n_n962 ) | ( wire468 ) | ( wire3340 ) ;
 assign wire3585 = ( n_n859 ) | ( n_n128 ) | ( n_n5  &  wire72 ) ;
 assign wire3587 = ( n_n1121 ) | ( wire140 ) | ( wire133 ) | ( wire3582 ) ;
 assign wire3588 = ( wire85 ) | ( wire276 ) | ( _8491 ) ;
 assign wire3589 = ( n_n602 ) | ( n_n1022 ) | ( n_n215 ) | ( n_n1023 ) ;
 assign wire3590 = ( wire3486 ) | ( wire3533 ) | ( _8494 ) ;
 assign wire3592 = ( wire348 ) | ( wire3467 ) | ( n_n1002 ) | ( wire95 ) ;
 assign wire3607 = ( wire546 ) | ( wire295 ) | ( _230 ) | ( _233 ) ;
 assign wire3610 = ( n_n1283 ) | ( n_n580 ) | ( n_n1334 ) ;
 assign wire3612 = ( wire331 ) | ( wire3610 ) | ( _8505 ) ;
 assign wire3613 = ( n_n858 ) | ( wire3462 ) | ( wire3464 ) | ( n_n95 ) ;
 assign wire3616 = ( wire318 ) | ( wire3605 ) | ( wire3613 ) ;
 assign wire3624 = ( n_n950 ) | ( n_n1208 ) | ( wire551 ) | ( wire153 ) ;
 assign wire3628 = ( o_18_ ) | ( wire237 ) | ( wire130 ) | ( wire3624 ) ;
 assign wire3631 = ( wire139 ) | ( wire3393 ) | ( wire179 ) | ( wire3628 ) ;
 assign wire3641 = ( wire197 ) | ( wire154 ) ;
 assign wire3643 = ( wire146 ) | ( n_n1  &  n_n18  &  wire67 ) ;
 assign wire3644 = ( wire183 ) | ( n_n0  &  wire69 ) ;
 assign wire3653 = ( n_n1022 ) | ( n_n1018 ) | ( wire3643 ) | ( wire3644 ) ;
 assign wire3654 = ( n_n215 ) | ( wire250 ) | ( n_n923 ) | ( wire3621 ) ;
 assign wire3655 = ( o_18_ ) | ( n_n387 ) | ( wire130 ) | ( _8613 ) ;
 assign wire3667 = ( n_n1122 ) | ( wire78 ) | ( n_n1165 ) ;
 assign wire3668 = ( n_n1137 ) | ( n_n962 ) | ( wire468 ) | ( wire3340 ) ;
 assign wire3669 = ( n_n864 ) | ( wire316 ) | ( wire158 ) ;
 assign wire3679 = ( n_n2  &  n_n12  &  n_n15 ) | ( n_n4  &  n_n12  &  n_n15 ) ;
 assign wire3682 = ( wire71  &  n_n1 ) | ( n_n1  &  n_n10  &  wire64 ) ;
 assign wire3686 = ( n_n1238 ) | ( n_n1239 ) | ( n_n1300 ) | ( n_n1315 ) ;
 assign wire3687 = ( o_9_ ) | ( n_n1301 ) | ( wire259 ) ;
 assign wire3688 = ( o_13_ ) | ( o_7_ ) | ( n_n1253 ) | ( n_n1268 ) ;
 assign wire3689 = ( o_6_ ) | ( n_n1225 ) | ( wire3679 ) ;
 assign wire3690 = ( n_n1316 ) | ( n_n1334 ) | ( n_n1254 ) | ( n_n1330 ) ;
 assign wire3692 = ( n_n1197 ) | ( wire88 ) | ( n_n822 ) ;
 assign wire3693 = ( n_n813 ) | ( wire183 ) | ( wire207 ) ;
 assign wire3695 = ( n_n961 ) | ( n_n1010 ) | ( wire109 ) | ( wire112 ) ;
 assign wire3702 = ( wire162 ) | ( wire159 ) | ( wire3682 ) | ( wire3693 ) ;
 assign wire3703 = ( wire3686 ) | ( wire3687 ) | ( wire3695 ) ;
 assign wire3704 = ( wire218 ) | ( wire3688 ) | ( wire3689 ) ;
 assign wire3712 = ( (~ i_7_)  &  i_6_  &  n_n7  &  n_n19 ) | ( i_7_  &  (~ i_6_)  &  n_n7  &  n_n19 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n7  &  n_n19 ) ;
 assign wire3713 = ( n_n1137 ) | ( n_n1135 ) | ( wire3712 ) ;
 assign wire3714 = ( i_7_  &  i_6_  &  n_n7  &  n_n2 ) | ( (~ i_7_)  &  i_6_  &  n_n7  &  n_n2 ) ;
 assign wire3715 = ( wire269 ) | ( wire3714 ) ;
 assign wire3716 = ( o_18_ ) | ( n_n1033 ) | ( wire130 ) ;
 assign wire3717 = ( wire250 ) | ( n_n923 ) | ( wire3621 ) | ( wire3715 ) ;
 assign wire3719 = ( o_30_ ) | ( o_7_ ) | ( wire127 ) ;
 assign wire3723 = ( wire77 ) | ( n_n1049 ) | ( wire99 ) | ( wire235 ) ;
 assign wire3724 = ( wire270 ) | ( n_n823 ) | ( wire189 ) ;
 assign wire3725 = ( n_n1136 ) | ( n_n1076 ) | ( n_n673 ) | ( wire3713 ) ;
 assign wire3736 = ( n_n1017 ) | ( n_n906 ) ;
 assign wire3739 = ( n_n1022 ) | ( wire3218 ) | ( _315 ) | ( _8729 ) ;
 assign wire3754 = ( n_n1017 ) | ( n_n1029 ) | ( n_n1  &  wire70 ) ;
 assign wire3756 = ( wire209 ) | ( n_n845 ) | ( wire292 ) ;
 assign wire3758 = ( n_n744 ) | ( n_n1215 ) | ( n_n745 ) | ( wire3754 ) ;
 assign wire3759 = ( n_n895 ) | ( n_n858 ) | ( wire3462 ) ;
 assign wire3760 = ( wire85 ) | ( wire3358 ) | ( wire3756 ) | ( _7830 ) ;
 assign wire3765 = ( wire165 ) | ( wire181 ) | ( wire3758 ) | ( wire3759 ) ;
 assign wire3770 = ( (~ i_7_)  &  i_6_  &  n_n2  &  n_n8 ) | ( i_7_  &  (~ i_6_)  &  n_n2  &  n_n8 ) ;
 assign wire3772 = ( o_7_ ) | ( n_n1268 ) | ( n_n554 ) ;
 assign wire3774 = ( n_n1271 ) | ( n_n1189 ) | ( n_n1  &  wire72 ) ;
 assign wire3775 = ( n_n1216 ) | ( n_n1244 ) | ( wire3770 ) ;
 assign wire3777 = ( wire186 ) | ( wire209 ) | ( n_n1223 ) | ( n_n1061 ) ;
 assign wire3781 = ( n_n1245 ) | ( wire287 ) | ( wire277 ) | ( wire308 ) ;
 assign wire3782 = ( n_n809 ) | ( n_n810 ) | ( wire3772 ) | ( wire3777 ) ;
 assign wire3784 = ( n_n904 ) | ( wire129 ) | ( wire107 ) ;
 assign wire3786 = ( wire112 ) | ( n_n802 ) | ( wire150 ) | ( wire3781 ) ;
 assign wire3789 = ( wire324 ) | ( wire3774 ) | ( wire3775 ) | ( wire3784 ) ;
 assign wire3792 = ( n_n427 ) | ( wire340 ) | ( wire3782 ) ;
 assign wire3796 = ( i_7_  &  i_6_  &  n_n5  &  n_n8 ) | ( (~ i_7_)  &  i_6_  &  n_n5  &  n_n8 ) | ( i_7_  &  (~ i_6_)  &  n_n5  &  n_n8 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n5  &  n_n8 ) ;
 assign wire3797 = ( wire3796 ) | ( n_n5  &  n_n14  &  wire72 ) ;
 assign wire3798 = ( wire271 ) | ( n_n17  &  n_n4  &  n_n13 ) ;
 assign wire3800 = ( n_n5  &  n_n12  &  n_n15 ) | ( n_n5  &  n_n10  &  n_n15 ) ;
 assign wire3801 = ( o_28_ ) | ( n_n1166 ) | ( wire78 ) | ( wire3800 ) ;
 assign wire3806 = ( n_n3  &  n_n12  &  n_n16 ) | ( n_n12  &  n_n1  &  n_n16 ) ;
 assign wire3807 = ( i_7_  &  (~ i_6_)  &  n_n2  &  n_n11 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n2  &  n_n11 ) ;
 assign wire3808 = ( n_n3  &  n_n13  &  n_n15 ) | ( n_n3  &  n_n9  &  n_n15 ) ;
 assign wire3809 = ( n_n1137 ) | ( n_n1135 ) | ( wire71  &  n_n3 ) ;
 assign wire3810 = ( wire127 ) | ( wire247 ) ;
 assign wire3813 = ( n_n1076 ) | ( wire3465 ) | ( n_n3  &  wire69 ) ;
 assign wire3816 = ( wire260 ) | ( wire3806 ) | ( wire3807 ) | ( wire3808 ) ;
 assign wire3818 = ( wire297 ) | ( n_n1147 ) | ( wire532 ) | ( wire3279 ) ;
 assign wire3820 = ( wire107 ) | ( wire217 ) | ( wire3809 ) | ( wire3810 ) ;
 assign wire3821 = ( wire250 ) | ( n_n923 ) | ( wire3621 ) | ( wire3816 ) ;
 assign wire3822 = ( wire270 ) | ( wire156 ) | ( wire3797 ) | ( wire3798 ) ;
 assign wire3823 = ( n_n859 ) | ( wire283 ) | ( wire3359 ) | ( wire3801 ) ;
 assign wire3827 = ( wire3296 ) | ( wire323 ) | ( _8855 ) ;
 assign wire3841 = ( wire134 ) | ( wire78 ) | ( wire158 ) | ( n_n825 ) ;
 assign wire3842 = ( o_8_ ) | ( wire346 ) | ( wire140 ) | ( wire133 ) ;
 assign wire3843 = ( wire187 ) | ( wire316 ) | ( wire235 ) | ( wire308 ) ;
 assign wire3844 = ( wire3841 ) | ( _8875 ) ;
 assign wire3850 = ( n_n1243 ) | ( n_n0  &  wire71 ) ;
 assign wire3853 = ( wire293 ) | ( wire109 ) ;
 assign wire3854 = ( o_9_ ) | ( n_n1300 ) | ( n_n1301 ) | ( n_n1315 ) ;
 assign wire3855 = ( wire259 ) | ( wire271 ) ;
 assign wire3856 = ( n_n1316 ) | ( n_n1287 ) | ( n_n814 ) | ( wire101 ) ;
 assign wire3857 = ( o_20_ ) | ( wire159 ) | ( wire135 ) | ( wire219 ) ;
 assign wire3860 = ( n_n813 ) | ( wire183 ) | ( wire207 ) ;
 assign wire3864 = ( n_n744 ) | ( wire104 ) | ( wire184 ) | ( n_n805 ) ;
 assign wire3868 = ( wire287 ) | ( wire305 ) ;
 assign wire3870 = ( n_n803 ) | ( wire97 ) | ( wire71  &  n_n3 ) ;
 assign wire3871 = ( wire77 ) | ( n_n935 ) | ( n_n1213 ) | ( wire3857 ) ;
 assign wire3872 = ( n_n1197 ) | ( wire88 ) | ( wire253 ) | ( wire3860 ) ;
 assign wire3873 = ( wire107 ) | ( n_n1034 ) | ( _8889 ) ;
 assign wire3874 = ( n_n824 ) | ( wire3850 ) | ( wire3864 ) ;
 assign wire3875 = ( wire3853 ) | ( wire3854 ) | ( wire3855 ) | ( wire3856 ) ;
 assign wire3877 = ( wire250 ) | ( wire3621 ) | ( n_n711 ) | ( wire3868 ) ;
 assign wire3883 = ( wire3872 ) | ( wire3873 ) | ( wire3874 ) | ( wire3875 ) ;
 assign wire3890 = ( wire93 ) | ( n_n1155 ) | ( wire160 ) ;
 assign wire3892 = ( wire3279 ) | ( wire3890 ) | ( _8932 ) ;
 assign wire3897 = ( n_n1169 ) | ( n_n821 ) | ( n_n1314 ) | ( n_n1165 ) ;
 assign wire3899 = ( n_n1180 ) | ( n_n817 ) | ( wire271 ) ;
 assign wire3900 = ( wire162 ) | ( n_n961 ) | ( wire291 ) | ( wire500 ) ;
 assign wire3903 = ( wire99 ) | ( n_n1322 ) | ( wire207 ) | ( wire3899 ) ;
 assign wire3905 = ( wire97 ) | ( wire3897 ) | ( _8923 ) ;
 assign wire3915 = ( o_10_ ) | ( n_n3  &  n_n12  &  n_n16 ) ;
 assign wire3916 = ( o_27_ ) | ( n_n1215 ) | ( wire277 ) ;
 assign wire3920 = ( wire261 ) | ( wire217 ) | ( wire3915 ) | ( wire3916 ) ;
 assign wire3926 = ( n_n573 ) | ( wire340 ) | ( wire3920 ) ;
 assign wire3929 = ( n_n17  &  n_n12 ) | ( n_n1  &  n_n10 ) ;
 assign wire3937 = ( n_n1238 ) | ( n_n1239 ) | ( n_n926 ) ;
 assign wire3938 = ( n_n930 ) | ( wire113 ) ;
 assign wire3939 = ( wire158 ) | ( wire161 ) ;
 assign wire3940 = ( o_9_ ) | ( o_8_ ) | ( n_n1302 ) | ( n_n872 ) ;
 assign wire3941 = ( n_n953 ) | ( n_n1288 ) | ( n_n1322 ) | ( n_n1139 ) ;
 assign wire3942 = ( n_n1203 ) | ( n_n1138 ) | ( wire273 ) | ( wire3929 ) ;
 assign wire3944 = ( wire354 ) | ( n_n1226 ) | ( wire77 ) | ( wire160 ) ;
 assign wire3945 = ( n_n1021 ) | ( n_n553 ) ;
 assign wire3950 = ( wire346 ) | ( wire3941 ) ;
 assign wire3951 = ( n_n859 ) | ( _8958 ) | ( wire72  &  _8622 ) ;
 assign wire3952 = ( o_18_ ) | ( wire130 ) | ( wire156 ) ;
 assign wire3955 = ( n_n923 ) | ( wire217 ) | ( wire3942 ) ;
 assign wire3957 = ( n_n1083 ) | ( wire104 ) | ( wire148 ) | ( _8976 ) ;
 assign wire3958 = ( wire3937 ) | ( wire3938 ) | ( wire3939 ) | ( wire3940 ) ;
 assign wire3962 = ( wire194 ) | ( n_n387 ) | ( n_n711 ) | ( wire295 ) ;
 assign wire3965 = ( wire3222 ) | ( n_n895 ) | ( wire173 ) | ( n_n534 ) ;
 assign wire3975 = ( wire209 ) | ( n_n1223 ) | ( wire112 ) | ( n_n802 ) ;
 assign wire3982 = ( o_9_ ) | ( n_n1302 ) | ( n_n553 ) ;
 assign wire3983 = ( n_n1021 ) | ( n_n1010 ) | ( wire265 ) ;
 assign wire3985 = ( n_n1017 ) | ( wire76 ) | ( wire3982 ) | ( wire3983 ) ;
 assign wire3993 = ( wire183 ) | ( n_n0  &  wire69 ) ;
 assign wire3994 = ( n_n1300 ) | ( wire266 ) | ( n_n1315 ) ;
 assign wire3995 = ( o_7_ ) | ( n_n1238 ) | ( n_n1147 ) | ( n_n1155 ) ;
 assign wire3997 = ( n_n1009 ) | ( wire127 ) | ( n_n1256 ) | ( wire471 ) ;
 assign wire3998 = ( wire147 ) | ( wire184 ) | ( wire545 ) | ( wire546 ) ;
 assign wire4001 = ( n_n1021 ) | ( n_n1020 ) | ( wire77 ) | ( n_n1049 ) ;
 assign wire4005 = ( wire3993 ) | ( wire3994 ) | ( wire3998 ) ;
 assign wire4006 = ( wire270 ) | ( wire229 ) | ( n_n642 ) | ( wire3797 ) ;
 assign wire4007 = ( n_n859 ) | ( wire156 ) | ( wire3798 ) | ( wire3801 ) ;
 assign wire4008 = ( wire140 ) | ( wire323 ) | ( wire3579 ) | ( wire3995 ) ;
 assign wire4009 = ( wire297 ) | ( n_n738 ) | ( wire3279 ) | ( wire4001 ) ;
 assign wire4019 = ( n_n1017 ) | ( n_n1024 ) | ( n_n1025 ) ;
 assign wire4020 = ( n_n1022 ) | ( n_n1298 ) | ( wire3218 ) | ( wire4019 ) ;
 assign wire4023 = ( n_n744 ) | ( n_n906 ) | ( wire268 ) | ( n_n745 ) ;
 assign wire4024 = ( n_n858 ) | ( wire3462 ) | ( wire325 ) ;
 assign wire4025 = ( wire298 ) | ( wire110 ) | ( wire303 ) | ( wire4023 ) ;
 assign wire4027 = ( wire270 ) | ( wire4024 ) | ( _8261 ) | ( _9052 ) ;
 assign wire4029 = ( wire4020 ) | ( wire4025 ) | ( _9061 ) ;
 assign wire4037 = ( o_30_ ) | ( n_n1261 ) | ( n_n1268 ) | ( n_n756 ) ;
 assign wire4038 = ( n_n949 ) | ( wire162 ) | ( wire243 ) ;
 assign wire4039 = ( n_n950 ) | ( wire159 ) | ( wire219 ) ;
 assign wire4042 = ( n_n1083 ) | ( wire127 ) | ( n_n616 ) | ( n_n617 ) ;
 assign wire4044 = ( wire77 ) | ( wire257 ) | ( _9083 ) ;
 assign wire4046 = ( wire173 ) | ( wire99 ) | ( wire235 ) | ( n_n948 ) ;
 assign wire4047 = ( wire135 ) | ( wire161 ) | ( wire4037 ) | ( wire4042 ) ;
 assign wire4051 = ( wire4038 ) | ( wire4039 ) | ( wire4044 ) ;
 assign wire4053 = ( wire301 ) | ( wire197 ) | ( wire270 ) | ( n_n823 ) ;
 assign wire4063 = ( n_n1321 ) | ( wire147 ) | ( wire281 ) | ( wire265 ) ;
 assign wire4065 = ( wire110 ) | ( n_n1320 ) | ( n_n1010 ) | ( wire4063 ) ;
 assign wire4066 = ( wire85 ) | ( wire132 ) | ( _148 ) | ( _9095 ) ;
 assign wire4071 = ( n_n10 ) | ( n_n7  &  n_n6  &  n_n14 ) ;
 assign wire4074 = ( wire88 ) | ( n_n5  &  wire72 ) ;
 assign wire4076 = ( n_n1163 ) | ( n_n1282 ) | ( wire4071 ) ;
 assign wire4079 = ( wire208 ) | ( wire269 ) | ( n_n1167 ) ;
 assign wire4081 = ( n_n953 ) | ( wire4076 ) | ( _7041 ) | ( _9116 ) ;
 assign wire4082 = ( wire76 ) | ( wire237 ) | ( n_n1322 ) | ( _7611 ) ;
 assign wire4083 = ( n_n955 ) | ( wire309 ) | ( _9120 ) ;
 assign wire4084 = ( wire130 ) | ( n_n925 ) | ( wire4074 ) | ( wire4079 ) ;
 assign wire4086 = ( wire139 ) | ( wire3393 ) | ( wire320 ) ;
 assign wire4090 = ( wire3296 ) | ( wire128 ) | ( n_n95 ) | ( n_n1334 ) ;
 assign wire4091 = ( wire331 ) | ( wire179 ) | ( n_n931 ) | ( wire4086 ) ;
 assign wire4092 = ( n_n901 ) | ( wire4081 ) | ( wire4082 ) | ( wire4083 ) ;
 assign wire4094 = ( n_n427 ) | ( wire4084 ) | ( wire4090 ) ;
 assign wire4099 = ( n_n1321 ) | ( wire3467 ) | ( wire95 ) | ( wire265 ) ;
 assign wire4100 = ( wire77 ) | ( n_n1049 ) | ( n_n1010 ) | ( _9151 ) ;
 assign wire4101 = ( wire270 ) | ( wire156 ) | ( wire3797 ) | ( wire3798 ) ;
 assign wire4105 = ( wire85 ) | ( wire83 ) | ( wire4020 ) | ( wire4101 ) ;
 assign wire4106 = ( n_n859 ) | ( wire333 ) | ( wire3801 ) | ( wire4099 ) ;
 assign wire4109 = ( wire193 ) | ( n_n989 ) | ( _9153 ) ;
 assign wire4113 = ( n_n0 ) | ( n_n8  &  n_n17  &  n_n1 ) ;
 assign wire4115 = ( wire162 ) | ( n_n582 ) | ( wire4113 ) ;
 assign wire4119 = ( n_n2  &  n_n12  &  n_n16 ) | ( n_n4  &  n_n12  &  n_n16 ) ;
 assign wire4122 = ( n_n0  &  n_n8  &  n_n16 ) | ( n_n8  &  n_n3  &  n_n16 ) ;
 assign wire4123 = ( n_n5  &  n_n12  &  n_n16 ) | ( n_n19  &  n_n12  &  n_n16 ) ;
 assign wire4125 = ( n_n5  &  n_n8  &  n_n16 ) | ( n_n8  &  n_n4  &  n_n16 ) ;
 assign wire4138 = ( n_n1137 ) | ( n_n826 ) | ( n_n1135 ) ;
 assign wire4139 = ( n_n1024 ) | ( n_n1  &  n_n10  &  wire67 ) ;
 assign wire4140 = ( o_11_ ) | ( n_n1302 ) | ( n_n1163 ) | ( n_n1256 ) ;
 assign wire4141 = ( n_n1258 ) | ( n_n1138 ) | ( n_n1167 ) | ( n_n1303 ) ;
 assign wire4142 = ( n_n1077 ) | ( n_n1301 ) | ( n_n1170 ) | ( n_n1273 ) ;
 assign wire4144 = ( n_n1076 ) | ( n_n909 ) | ( n_n910 ) ;
 assign wire4145 = ( n_n1274 ) | ( n_n1298 ) | ( wire3218 ) | ( wire281 ) ;
 assign wire4149 = ( n_n797 ) | ( n_n1322 ) | ( _8171 ) | ( _9191 ) ;
 assign wire4150 = ( wire226 ) | ( wire309 ) | ( wire4144 ) ;
 assign wire4151 = ( wire147 ) | ( wire300 ) | ( wire4138 ) | ( wire4145 ) ;
 assign wire4152 = ( wire4139 ) | ( wire4140 ) | ( wire4141 ) | ( wire4142 ) ;
 assign wire4153 = ( n_n459 ) | ( wire216 ) | ( wire3304 ) | ( wire3305 ) ;
 assign wire4154 = ( wire132 ) | ( wire3361 ) | ( _148 ) | ( _9187 ) ;
 assign _88 = ( (~ i_7_)  &  (~ i_6_)  &  n_n5  &  n_n8 ) ;
 assign _92 = ( i_1_  &  (~ i_2_)  &  (~ i_0_)  &  wire70 ) ;
 assign _94 = ( i_7_  &  i_6_  &  n_n6  &  n_n11 ) ;
 assign _100 = ( (~ i_1_)  &  (~ i_2_)  &  (~ i_0_)  &  wire72 ) ;
 assign _111 = ( (~ i_7_)  &  i_6_  &  n_n0  &  n_n11 ) ;
 assign _113 = ( i_7_  &  (~ i_6_)  &  n_n8  &  n_n19 ) ;
 assign _115 = ( (~ i_7_)  &  (~ i_6_)  &  n_n8  &  n_n19 ) ;
 assign _119 = ( i_7_  &  i_6_  &  n_n0  &  n_n8 ) ;
 assign _121 = ( i_7_  &  i_6_  &  n_n12  &  n_n1 ) ;
 assign _148 = ( (~ i_7_)  &  i_6_  &  n_n7  &  n_n2 ) ;
 assign _173 = ( (~ i_7_)  &  (~ i_6_)  &  n_n6  &  n_n12 ) ;
 assign _175 = ( i_7_  &  (~ i_6_)  &  n_n11  &  n_n1 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n11  &  n_n1 ) ;
 assign _177 = ( i_7_  &  i_6_  &  n_n1  &  n_n9 ) | ( (~ i_7_)  &  i_6_  &  n_n1  &  n_n9 ) | ( i_7_  &  (~ i_6_)  &  n_n1  &  n_n9 ) ;
 assign _192 = ( i_7_  &  (~ i_6_)  &  n_n6  &  n_n12 ) ;
 assign _225 = ( i_7_  &  i_6_  &  n_n9 ) ;
 assign _230 = ( i_1_  &  (~ i_2_)  &  (~ i_0_)  &  wire69 ) ;
 assign _233 = ( (~ i_7_)  &  i_6_  &  n_n3  &  n_n10 ) | ( i_7_  &  (~ i_6_)  &  n_n3  &  n_n10 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n3  &  n_n10 ) ;
 assign _271 = ( (~ i_7_)  &  i_6_  &  n_n5  &  n_n9 ) | ( i_7_  &  (~ i_6_)  &  n_n5  &  n_n9 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n5  &  n_n9 ) ;
 assign _302 = ( i_7_  &  (~ i_6_)  &  n_n8  &  n_n4 ) ;
 assign _315 = ( (~ i_7_)  &  (~ i_6_)  &  n_n1  &  n_n9 ) ;
 assign _327 = ( i_1_  &  i_2_  &  (~ i_0_)  &  wire69 ) ;
 assign _363 = ( i_7_  &  i_6_  &  n_n2  &  n_n13 ) | ( (~ i_7_)  &  i_6_  &  n_n2  &  n_n13 ) | ( i_7_  &  (~ i_6_)  &  n_n2  &  n_n13 ) ;
 assign _420 = ( (~ i_7_)  &  (~ i_6_)  &  n_n7  &  n_n3 ) ;
 assign _473 = ( i_7_  &  i_6_  &  n_n0  &  n_n18 ) | ( (~ i_7_)  &  i_6_  &  n_n0  &  n_n18 ) | ( i_7_  &  (~ i_6_)  &  n_n0  &  n_n18 ) ;
 assign _475 = ( (~ i_7_)  &  i_6_  &  n_n2  &  n_n10 ) | ( i_7_  &  (~ i_6_)  &  n_n2  &  n_n10 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n2  &  n_n10 ) ;
 assign _485 = ( i_7_  &  i_6_  &  n_n2  &  n_n11 ) ;
 assign _540 = ( i_7_  &  i_6_  &  n_n0  &  n_n7 ) ;
 assign _583 = ( i_7_  &  i_6_  &  n_n5  &  n_n18 ) ;
 assign _605 = ( i_7_  &  i_6_  &  n_n8  &  n_n19 ) ;
 assign _646 = ( (~ i_7_)  &  i_6_  &  n_n4  &  n_n18 ) | ( i_7_  &  (~ i_6_)  &  n_n4  &  n_n18 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n4  &  n_n18 ) ;
 assign _713 = ( (~ i_7_)  &  (~ i_6_)  &  n_n0  &  n_n11 ) ;
 assign _787 = ( i_7_  &  (~ i_6_)  &  n_n4  &  n_n11 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n4  &  n_n11 ) ;
 assign _6938 = ( i_7_  &  i_6_  &  n_n3  &  n_n18 ) | ( (~ i_7_)  &  i_6_  &  n_n3  &  n_n18 ) ;
 assign _6943 = ( o_15_ ) | ( n_n1215 ) | ( wire3221 ) | ( _6938 ) ;
 assign _6944 = ( i_6_  &  (~ i_7_) ) ;
 assign _6968 = ( wire88 ) | ( n_n4  &  n_n11  &  _6944 ) ;
 assign _7024 = ( (~ i_6_)  &  (~ i_7_) ) ;
 assign _7041 = ( (~ i_7_)  &  i_6_  &  n_n4  &  n_n11 ) | ( i_7_  &  (~ i_6_)  &  n_n4  &  n_n11 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n4  &  n_n11 ) ;
 assign _7043 = ( n_n1203 ) | ( n_n953 ) | ( wire273 ) | ( _7041 ) ;
 assign _7056 = ( (~ i_7_)  &  i_6_  &  n_n3  &  n_n12 ) | ( i_7_  &  (~ i_6_)  &  n_n3  &  n_n12 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n3  &  n_n12 ) ;
 assign _7076 = ( i_7_  &  i_6_  &  n_n5  &  n_n12 ) | ( (~ i_7_)  &  i_6_  &  n_n5  &  n_n12 ) | ( i_7_  &  (~ i_6_)  &  n_n5  &  n_n12 ) ;
 assign _7160 = ( n_n1320 ) | ( wire265 ) | ( _713 ) ;
 assign _7201 = ( n_n949 ) | ( wire162 ) | ( wire243 ) ;
 assign _7234 = ( n_n845 ) | ( n_n858 ) | ( wire3245 ) | ( _7201 ) ;
 assign _7256 = ( n_n1020 ) | ( n_n1021 ) ;
 assign _7275 = ( i_6_  &  i_7_ ) ;
 assign _7295 = ( i_1_  &  (~ i_2_)  &  (~ i_0_) ) ;
 assign _7316 = ( i_6_  &  (~ i_7_) ) ;
 assign _7318 = ( i_6_  &  i_7_ ) ;
 assign _7320 = ( (~ i_6_)  &  (~ i_7_) ) ;
 assign _7324 = ( i_7_  &  i_6_  &  n_n6  &  n_n11 ) | ( (~ i_7_)  &  i_6_  &  n_n6  &  n_n11 ) ;
 assign _7325 = ( i_7_  &  (~ i_6_)  &  n_n6  &  n_n12 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n6  &  n_n12 ) ;
 assign _7326 = ( n_n1009 ) | ( _646 ) | ( wire69  &  _7295 ) ;
 assign _7362 = ( i_6_  &  i_7_ ) ;
 assign _7435 = ( n_n1121 ) | ( wire133 ) | ( _605 ) ;
 assign _7451 = ( (~ i_6_)  &  i_7_ ) ;
 assign _7486 = ( i_6_  &  i_7_ ) ;
 assign _7583 = ( (~ i_7_)  &  i_6_  &  n_n4  &  n_n10 ) | ( i_7_  &  (~ i_6_)  &  n_n4  &  n_n10 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n4  &  n_n10 ) ;
 assign _7611 = ( i_7_  &  (~ i_6_)  &  n_n0  &  n_n11 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n0  &  n_n11 ) ;
 assign _7620 = ( (~ i_6_)  &  (~ i_7_) ) ;
 assign _7638 = ( n_n1316 ) | ( wire128 ) | ( _540 ) ;
 assign _7788 = ( n_n1274 ) | ( wire281 ) | ( n_n1032 ) ;
 assign _7795 = ( n_n1321 ) | ( wire88 ) | ( wire265 ) | ( _475 ) ;
 assign _7798 = ( i_6_  &  i_7_ ) ;
 assign _7801 = ( wire128 ) | ( n_n0  &  n_n7  &  _7798 ) ;
 assign _7818 = ( i_1_  &  i_2_  &  (~ i_0_) ) ;
 assign _7830 = ( i_7_  &  i_6_  &  n_n3  &  n_n11 ) | ( (~ i_7_)  &  i_6_  &  n_n3  &  n_n11 ) ;
 assign _7839 = ( n_n805 ) | ( wire135 ) | ( wire3358 ) | ( _7830 ) ;
 assign _7869 = ( n_n1009 ) | ( wire471 ) | ( wire133 ) | ( _605 ) ;
 assign _7921 = ( i_1_  &  (~ i_2_)  &  i_0_ ) ;
 assign _7923 = ( i_7_  &  i_6_  &  n_n7  &  n_n19 ) | ( (~ i_7_)  &  i_6_  &  n_n7  &  n_n19 ) | ( i_7_  &  (~ i_6_)  &  n_n7  &  n_n19 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n7  &  n_n19 ) ;
 assign _7931 = ( n_n1121 ) | ( wire353 ) | ( wire308 ) | ( _7923 ) ;
 assign _7932 = ( n_n1180 ) | ( n_n822 ) | ( n_n1181 ) | ( wire507 ) ;
 assign _7991 = ( wire277 ) | ( wire112 ) | ( n_n802 ) | ( _420 ) ;
 assign _7993 = ( wire270 ) | ( n_n573 ) | ( n_n826 ) | ( _7932 ) ;
 assign _7994 = ( wire3344 ) | ( wire462 ) | ( _7931 ) ;
 assign _8022 = ( n_n1320 ) | ( wire265 ) | ( _713 ) ;
 assign _8053 = ( wire287 ) | ( n_n1268 ) | ( wire132 ) | ( n_n574 ) ;
 assign _8108 = ( (~ i_7_)  &  i_6_  &  n_n8  &  n_n3 ) | ( i_7_  &  (~ i_6_)  &  n_n8  &  n_n3 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n8  &  n_n3 ) ;
 assign _8115 = ( (~ i_6_)  &  (~ i_7_) ) ;
 assign _8117 = ( i_7_  &  (~ i_6_)  &  n_n3  &  n_n11 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n3  &  n_n11 ) ;
 assign _8134 = ( wire112 ) | ( wire292 ) | ( _8108 ) | ( _8117 ) ;
 assign _8137 = ( i_6_  &  i_7_ ) ;
 assign _8159 = ( wire285 ) | ( wire237 ) | ( wire139 ) | ( wire3393 ) ;
 assign _8171 = ( i_7_  &  (~ i_6_)  &  n_n0  &  n_n11 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n0  &  n_n11 ) ;
 assign _8174 = ( wire155 ) | ( n_n1322 ) | ( n_n1319 ) | ( _8171 ) ;
 assign _8175 = ( wire128 ) | ( n_n0  &  n_n9  &  _7620 ) ;
 assign _8176 = ( n_n1121 ) | ( n_n906 ) | ( wire353 ) | ( _7923 ) ;
 assign _8178 = ( wire3443 ) | ( _8174 ) | ( _8175 ) | ( _8176 ) ;
 assign _8180 = ( wire487 ) | ( wire488 ) | ( wire3311 ) ;
 assign _8188 = ( n_n1283 ) | ( n_n580 ) | ( wire260 ) | ( n_n582 ) ;
 assign _8190 = ( wire148 ) | ( wire3432 ) | ( _8180 ) ;
 assign _8193 = ( i_7_  &  i_6_  &  n_n5  &  n_n10 ) | ( (~ i_7_)  &  i_6_  &  n_n5  &  n_n10 ) ;
 assign _8194 = ( wire466 ) | ( wire93 ) ;
 assign _8200 = ( n_n1203 ) | ( n_n953 ) | ( wire273 ) | ( _7041 ) ;
 assign _8211 = ( wire194 ) | ( wire3433 ) | ( _8194 ) | ( _8200 ) ;
 assign _8222 = ( wire461 ) | ( wire3341 ) | ( wire3342 ) ;
 assign _8233 = ( o_15_ ) | ( n_n1223 ) | ( wire3465 ) | ( wire414 ) ;
 assign _8234 = ( wire77 ) | ( n_n1049 ) | ( _327 ) | ( _8233 ) ;
 assign _8235 = ( wire462 ) | ( _7931 ) | ( _8222 ) | ( _8234 ) ;
 assign _8241 = ( i_7_  &  (~ i_6_)  &  n_n2  &  n_n12 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n2  &  n_n12 ) ;
 assign _8245 = ( n_n822 ) | ( wire189 ) | ( n_n821 ) | ( wire421 ) ;
 assign _8257 = ( wire292 ) | ( n_n3  &  n_n11  &  _8115 ) ;
 assign _8258 = ( o_13_ ) | ( n_n1253 ) | ( n_n1254 ) | ( n_n1040 ) ;
 assign _8259 = ( wire87 ) | ( _7788 ) | ( _8257 ) | ( _8258 ) ;
 assign _8261 = ( n_n1180 ) | ( n_n826 ) | ( n_n1181 ) | ( wire507 ) ;
 assign _8276 = ( wire88 ) | ( n_n4  &  n_n11  &  _6944 ) ;
 assign _8277 = ( n_n1194 ) | ( n_n1196 ) | ( n_n845 ) | ( wire242 ) ;
 assign _8292 = ( wire270 ) | ( _8261 ) | ( _8276 ) | ( _8277 ) ;
 assign _8295 = ( wire3482 ) | ( wire3355 ) | ( _8235 ) ;
 assign _8309 = ( n_n845 ) | ( wire128 ) ;
 assign _8315 = ( n_n1257 ) | ( n_n554 ) | ( n_n1  &  wire72 ) ;
 assign _8318 = ( i_7_  &  i_6_  &  n_n0  &  n_n12 ) | ( (~ i_7_)  &  i_6_  &  n_n0  &  n_n12 ) | ( i_7_  &  (~ i_6_)  &  n_n0  &  n_n12 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n0  &  n_n12 ) ;
 assign _8328 = ( n_n1245 ) | ( wire277 ) | ( wire112 ) | ( n_n802 ) ;
 assign _8329 = ( wire3305 ) | ( wire3304 ) ;
 assign _8332 = ( wire270 ) | ( n_n823 ) | ( wire3361 ) | ( _8328 ) ;
 assign _8384 = ( n_n1032 ) | ( wire292 ) | ( _8117 ) ;
 assign _8387 = ( wire128 ) | ( wire3545 ) | ( wire3546 ) | ( _540 ) ;
 assign _8418 = ( n_n1049 ) | ( n_n1320 ) | ( n_n1010 ) ;
 assign _8423 = ( wire3433 ) | ( wire3548 ) | ( _8194 ) | ( _8418 ) ;
 assign _8425 = ( n_n1137 ) | ( n_n6  &  n_n12  &  _7320 ) ;
 assign _8455 = ( n_n1083 ) | ( wire3577 ) ;
 assign _8456 = ( wire186 ) | ( wire236 ) | ( n_n958 ) | ( wire592 ) ;
 assign _8458 = ( n_n996 ) | ( _485 ) | ( _8455 ) | ( _8456 ) ;
 assign _8479 = ( n_n1074 ) | ( wire286 ) | ( wire316 ) ;
 assign _8489 = ( (~ i_7_) ) | ( (~ i_6_) ) | ( i_7_  &  i_6_  &  n_n4  &  n_n13 ) ;
 assign _8491 = ( n_n1021 ) | ( n_n953 ) | ( _473 ) | ( _8489 ) ;
 assign _8494 = ( o_20_ ) | ( wire292 ) | ( _302 ) | ( _8117 ) ;
 assign _8503 = ( i_1_  &  (~ i_2_)  &  (~ i_0_) ) ;
 assign _8505 = ( wire208 ) | ( n_n1010 ) | ( wire72  &  _8503 ) ;
 assign _8510 = ( n_n1238 ) | ( n_n1239 ) | ( n_n937 ) ;
 assign _8513 = ( wire3238 ) | ( wire3432 ) | ( _8510 ) ;
 assign _8515 = ( wire88 ) | ( n_n4  &  n_n11  &  _6944 ) ;
 assign _8519 = ( i_7_  &  i_6_  &  n_n7  &  n_n2 ) | ( (~ i_7_)  &  i_6_  &  n_n7  &  n_n2 ) ;
 assign _8530 = ( i_7_  &  i_6_  &  n_n0  &  n_n7 ) | ( (~ i_7_)  &  i_6_  &  n_n0  &  n_n7 ) ;
 assign _8533 = ( n_n573 ) | ( n_n990 ) | ( n_n574 ) ;
 assign _8535 = ( wire218 ) | ( wire279 ) | ( n_n1010 ) | ( _225 ) ;
 assign _8546 = ( wire3345 ) | ( wire238 ) | ( _8222 ) | ( _8535 ) ;
 assign _8549 = ( wire318 ) | ( wire3605 ) | ( wire319 ) | ( _8533 ) ;
 assign _8561 = ( i_7_  &  i_6_  &  n_n4  &  n_n10 ) | ( (~ i_7_)  &  i_6_  &  n_n4  &  n_n10 ) | ( i_7_  &  (~ i_6_)  &  n_n4  &  n_n10 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n4  &  n_n10 ) ;
 assign _8569 = ( n_n817 ) | ( n_n814 ) ;
 assign _8594 = ( wire254 ) | ( wire132 ) | ( n_n1275 ) ;
 assign _8610 = ( n_n1300 ) | ( n_n1258 ) | ( wire257 ) ;
 assign _8613 = ( wire77 ) | ( wire300 ) | ( wire247 ) | ( _7056 ) ;
 assign _8615 = ( n_n1021 ) | ( wire112 ) | ( _473 ) | ( _8108 ) ;
 assign _8616 = ( wire226 ) | ( _8610 ) | ( _8615 ) ;
 assign _8617 = ( wire3345 ) | ( wire3654 ) | ( _8222 ) | ( _8594 ) ;
 assign _8619 = ( wire3639 ) | ( wire189 ) | ( wire97 ) | ( _8569 ) ;
 assign _8622 = ( (~ i_1_)  &  i_2_  &  i_0_ ) ;
 assign _8626 = ( wire93 ) | ( wire466 ) | ( wire133 ) | ( _605 ) ;
 assign _8647 = ( wire77 ) | ( wire254 ) | ( n_n1028 ) | ( n_n1213 ) ;
 assign _8692 = ( o_10_ ) | ( wire197 ) | ( wire112 ) | ( n_n802 ) ;
 assign _8698 = ( n_n1121 ) | ( wire257 ) | ( wire133 ) ;
 assign _8700 = ( wire140 ) | ( wire284 ) | ( wire3719 ) | ( _8698 ) ;
 assign _8701 = ( n_n817 ) | ( n_n814 ) ;
 assign _8710 = ( wire154 ) | ( wire97 ) | ( wire3716 ) | ( _8701 ) ;
 assign _8711 = ( wire128 ) | ( n_n0  &  n_n7  &  _7798 ) ;
 assign _8716 = ( wire3296 ) | ( n_n609 ) | ( _8479 ) | ( _8711 ) ;
 assign _8718 = ( n_n660 ) | ( wire3725 ) | ( _8692 ) | ( _8700 ) ;
 assign _8720 = ( wire197 ) | ( wire154 ) ;
 assign _8722 = ( n_n1040 ) | ( n_n2  &  n_n11  &  _8137 ) ;
 assign _8726 = ( n_n817 ) | ( n_n814 ) ;
 assign _8729 = ( n_n1025 ) | ( wire128 ) | ( _177 ) | ( _540 ) ;
 assign _8730 = ( wire87 ) | ( wire97 ) | ( _7788 ) | ( _8726 ) ;
 assign _8733 = ( wire3745 ) | ( wire3355 ) | ( _8235 ) ;
 assign _8737 = ( o_9_ ) | ( n_n1302 ) | ( n_n1024 ) | ( n_n1301 ) ;
 assign _8738 = ( wire3218 ) | ( n_n1025 ) | ( _315 ) ;
 assign _8740 = ( n_n1021 ) | ( wire568 ) | ( _175 ) ;
 assign _8741 = ( n_n1020 ) | ( n_n1028 ) | ( wire162 ) | ( wire243 ) ;
 assign _8742 = ( _8737 ) | ( _8738 ) | ( _8740 ) | ( _8741 ) ;
 assign _8745 = ( wire108 ) | ( wire337 ) | ( wire3433 ) | ( _8194 ) ;
 assign _8759 = ( n_n468 ) | ( wire140 ) | ( wire284 ) | ( _7435 ) ;
 assign _8760 = ( wire3436 ) | ( _8745 ) | ( _8759 ) ;
 assign _8762 = ( n_n858 ) | ( n_n845 ) ;
 assign _8855 = ( o_11_ ) | ( wire128 ) | ( _540 ) | ( _583 ) ;
 assign _8860 = ( o_15_ ) | ( n_n1223 ) | ( n_n845 ) | ( wire414 ) ;
 assign _8875 = ( wire94 ) | ( n_n872 ) | ( wire564 ) | ( _7076 ) ;
 assign _8876 = ( n_n1009 ) | ( n_n19  &  n_n12  &  _7451 ) ;
 assign _8882 = ( wire152 ) | ( n_n673 ) | ( wire3283 ) | ( _8876 ) ;
 assign _8889 = ( wire248 ) | ( wire260 ) | ( _119 ) | ( _121 ) ;
 assign _8905 = ( wire3842 ) | ( wire3843 ) | ( wire3844 ) | ( _8882 ) ;
 assign _8906 = ( wire314 ) | ( wire95 ) | ( wire320 ) | ( _8860 ) ;
 assign _8910 = ( n_n1009 ) | ( wire134 ) | ( _113 ) | ( _115 ) ;
 assign _8915 = ( wire129 ) | ( wire107 ) | ( wire3900 ) ;
 assign _8923 = ( n_n1017 ) | ( wire76 ) | ( n_n814 ) ;
 assign _8927 = ( wire287 ) | ( n_n1268 ) | ( wire132 ) | ( n_n574 ) ;
 assign _8932 = ( wire222 ) | ( n_n5  &  n_n13 ) | ( n_n5  &  wire70 ) ;
 assign _8934 = ( wire3296 ) | ( wire337 ) | ( _8425 ) | ( _8711 ) ;
 assign _8941 = ( wire3358 ) | ( n_n1322 ) | ( _7830 ) | ( _8171 ) ;
 assign _8950 = ( n_n468 ) | ( wire140 ) | ( wire284 ) | ( _7435 ) ;
 assign _8951 = ( wire3436 ) | ( _8745 ) | ( _8950 ) ;
 assign _8952 = ( wire3921 ) | ( n_n895 ) | ( wire3441 ) | ( _8941 ) ;
 assign _8954 = ( wire331 ) | ( wire72  &  _8503 ) ;
 assign _8958 = ( n_n1017 ) | ( wire76 ) ;
 assign _8974 = ( i_7_  &  i_6_  &  n_n6  &  n_n11 ) | ( (~ i_7_)  &  i_6_  &  n_n6  &  n_n11 ) ;
 assign _8975 = ( i_7_  &  (~ i_6_)  &  n_n6  &  n_n12 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n6  &  n_n12 ) ;
 assign _8976 = ( wire134 ) | ( _115 ) | ( _8974 ) | ( _8975 ) ;
 assign _9005 = ( wire3638 ) | ( n_n809 ) ;
 assign _9008 = ( i_7_  &  (~ i_6_)  &  n_n7  &  n_n3 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n7  &  n_n3 ) ;
 assign _9009 = ( _9008 ) | ( wire277 ) ;
 assign _9011 = ( wire197 ) | ( wire154 ) | ( wire3975 ) | ( _9009 ) ;
 assign _9012 = ( n_n490 ) | ( wire462 ) | ( _7931 ) | ( _8222 ) ;
 assign _9019 = ( wire148 ) | ( wire150 ) | ( wire107 ) | ( _8188 ) ;
 assign _9021 = ( n_n476 ) | ( wire264 ) | ( wire3985 ) | ( _9019 ) ;
 assign _9032 = ( n_n1083 ) | ( wire236 ) | ( wire473 ) ;
 assign _9035 = ( n_n1253 ) | ( n_n3  &  n_n10  &  _7362 ) ;
 assign _9037 = ( n_n1022 ) | ( wire3716 ) | ( wire3997 ) | ( _9035 ) ;
 assign _9052 = ( wire197 ) | ( wire154 ) ;
 assign _9061 = ( wire85 ) | ( wire87 ) | ( _7256 ) | ( _7788 ) ;
 assign _9065 = ( wire3345 ) | ( wire77 ) | ( n_n1049 ) | ( _8222 ) ;
 assign _9068 = ( n_n1121 ) | ( wire133 ) | ( _605 ) ;
 assign _9071 = ( n_n1076 ) | ( n_n673 ) | ( wire3713 ) | ( _94 ) ;
 assign _9083 = ( (~ i_7_)  &  i_6_  &  n_n3  &  n_n12 ) | ( i_7_  &  (~ i_6_)  &  n_n3  &  n_n12 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n3  &  n_n12 ) ;
 assign _9087 = ( n_n858 ) | ( n_n845 ) ;
 assign _9088 = ( wire114 ) | ( wire3216 ) | ( _7160 ) | ( _9087 ) ;
 assign _9095 = ( n_n1017 ) | ( wire76 ) ;
 assign _9097 = ( _8737 ) | ( _8738 ) | ( _8740 ) | ( _8741 ) ;
 assign _9099 = ( (~ i_1_)  &  (~ i_2_)  &  (~ i_0_) ) ;
 assign _9104 = ( n_n990 ) | ( wire72  &  _9099 ) ;
 assign _9107 = ( wire3238 ) | ( wire3432 ) | ( _8510 ) ;
 assign _9116 = ( wire273 ) | ( n_n4  &  n_n10  &  _7024 ) ;
 assign _9120 = ( n_n961 ) | ( wire271 ) | ( _88 ) | ( _271 ) ;
 assign _9141 = ( n_n1137 ) | ( wire337 ) | ( _173 ) ;
 assign _9151 = ( i_7_  &  i_6_  &  n_n0  &  n_n11 ) | ( (~ i_7_)  &  i_6_  &  n_n0  &  n_n11 ) | ( i_7_  &  (~ i_6_)  &  n_n0  &  n_n11 ) ;
 assign _9153 = ( wire87 ) | ( wire4100 ) | ( _7788 ) ;
 assign _9162 = ( n_n476 ) | ( wire4117 ) ;
 assign _9187 = ( wire277 ) | ( wire112 ) | ( n_n802 ) | ( _420 ) ;
 assign _9191 = ( wire155 ) | ( wire3363 ) | ( _111 ) ;


endmodule

