module pdc_mapped (
	i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_14_, i_3_, 
	i_13_, i_4_, i_12_, i_1_, i_11_, i_2_, i_0_, i_15_, o_1_, o_19_, 
	o_2_, o_0_, o_29_, o_39_, o_38_, o_25_, o_12_, o_37_, o_26_, o_11_, 
	o_36_, o_27_, o_14_, o_35_, o_28_, o_13_, o_34_, o_21_, o_16_, o_33_, 
	o_22_, o_15_, o_32_, o_23_, o_18_, o_31_, o_24_, o_17_, o_30_, o_20_, 
	o_10_, o_9_, o_7_, o_8_, o_5_, o_6_, o_3_, o_4_);

input i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_14_, i_3_, i_13_, i_4_, i_12_, i_1_, i_11_, i_2_, i_0_, i_15_;

output o_1_, o_19_, o_2_, o_0_, o_29_, o_39_, o_38_, o_25_, o_12_, o_37_, o_26_, o_11_, o_36_, o_27_, o_14_, o_35_, o_28_, o_13_, o_34_, o_21_, o_16_, o_33_, o_22_, o_15_, o_32_, o_23_, o_18_, o_31_, o_24_, o_17_, o_30_, o_20_, o_10_, o_9_, o_7_, o_8_, o_5_, o_6_, o_3_, o_4_;

wire n_n5231, wire19373, wire19374, n_n3621, wire19592, wire19593, wire19601, wire19622, wire19648, n_n5792, n_n5794, wire19766, wire19822, wire19846, wire19847, n_n4718, wire19989, wire19990, n_n264, n_n153, n_n120, wire20002, wire20004, n_n5224, n_n2657, wire20115, wire20245, wire20355, n_n2789, n_n2795, wire20625, n_n4508, wire20648, n_n4186, wire20658, wire879, wire20665, n_n5797, wire20667, wire20671, wire20753, n_n5235, wire3945, wire20920, wire20924, n_n3089, n_n3094, wire21154, wire21178, n_n3892, n_n3890, wire21293, n_n2058, wire21620, wire21621, n_n1670, wire21904, wire22331, wire22334, wire2474, wire22594, wire22847, n_n260, n_n229, n_n165, n_n139, wire913, n_n151, n_n116, n_n5686, wire590, wire19306, wire19359, wire19365, wire48, wire503, n_n152, n_n4476, n_n220, wire54, n_n4477, wire394, wire927, wire929, wire507, n_n111, wire103, wire266, wire893, n_n208, n_n273, wire937, wire372, wire386, wire19380, n_n3424, n_n3642, wire19431, wire19435, n_n3625, n_n3382, wire19445, wire19446, wire19455, n_n3626, n_n3645, wire19472, wire19473, wire19480, n_n3627, wire19530, n_n4781, n_n3711, wire19544, wire19546, n_n3631, wire19553, wire19554, n_n3661, n_n3632, n_n284, n_n124, n_n123, wire289, wire364, wire535, wire777, n_n118, wire834, n_n281, wire914, wire907, wire939, n_n110, n_n106, n_n5678, n_n5671, wire396, wire880, n_n5677, n_n5672, wire582, wire5453, wire19613, wire19614, wire583, wire941, wire940, n_n272, wire19624, wire19625, wire19626, n_n4442, n_n4439, wire943, n_n231, wire19290, wire573, wire5389, wire19654, wire19655, n_n4203, n_n4846, n_n4842, wire19659, n_n4206, n_n1506, wire19677, n_n6, wire911, n_n228, wire75, n_n4807, n_n4808, n_n4809, wire541, n_n4223, wire585, wire5347, wire5348, n_n4224, n_n4307, wire19717, wire19718, n_n285, n_n1, n_n283, n_n2, n_n60, wire118, n_n2618, n_n206, wire72, n_n5769, n_n127, wire19835, n_n242, n_n279, n_n266, n_n265, n_n271, n_n268, wire273, n_n2550, wire5115, wire5116, wire19849, n_n2545, wire268, wire200, wire112, n_n155, n_n5796, n_n5, n_n4723, n_n4725, wire19980, wire19981, wire4935, n_n2772, n_n230, n_n130, n_n121, n_n132, wire1686, wire20007, wire1705, wire20008, wire949, wire905, wire948, n_n4416, n_n4418, wire20033, wire20034, n_n4549, n_n4544, wire20147, n_n4533, wire20166, wire20184, n_n4556, n_n4535, wire20240, n_n3900, n_n3899, n_n3901, n_n3918, n_n3919, wire20353, n_n4141, n_n4, wire912, wire95, n_n4015, n_n2793, wire20571, wire20614, n_n3727, n_n9, wire4264, n_n2840, wire4259, wire20616, wire20617, n_n2839, n_n128, n_n5682, n_n5676, wire20629, wire20630, wire826, wire4234, wire4235, wire4236, wire216, n_n255, wire894, wire20651, wire20652, n_n241, n_n54, n_n105, wire392, n_n177, n_n216, n_n45, wire559, wire902, n_n258, wire950, wire20662, wire926, wire19753, wire19754, wire19758, n_n4219, n_n4199, wire20718, n_n3361, n_n3360, wire20913, wire20914, n_n163, wire19294, n_n5693, n_n274, wire452, wire19296, wire758, wire923, wire20925, wire20926, n_n3140, n_n7424, n_n3, n_n8, n_n61, n_n4005, wire446, wire20946, wire20947, n_n3138, n_n3092, n_n3093, wire21131, n_n3107, n_n3108, wire21148, n_n133, wire21186, n_n3898, n_n3895, wire21220, n_n3914, n_n3915, n_n3897, n_n3913, wire3626, wire21276, n_n57, n_n56, n_n226, wire4059, wire4060, n_n2440, n_n257, wire208, wire199, wire955, n_n2073, n_n2108, wire21396, n_n145, wire21440, n_n2067, wire21508, n_n2081, n_n2080, n_n2063, n_n2085, n_n2083, n_n2064, wire21612, wire169, n_n126, n_n5660, n_n5659, wire581, wire21635, n_n1689, n_n1692, wire21881, wire21885, n_n1724, wire21896, n_n1693, n_n37, n_n83, wire154, wire64, n_n1111, wire2808, wire21999, wire22014, n_n1089, n_n240, n_n246, wire1345, wire22360, wire22361, n_n380, wire1347, wire1346, n_n381, wire2163, wire2169, wire22602, n_n741, n_n740, wire22827, n_n775, wire1837, wire22839, n_n282, n_n225, wire126, n_n189, wire6004, wire19279, wire19280, n_n5053, wire5936, wire19191, wire19192, n_n5061, wire5931, wire19194, wire19195, n_n5062, wire5922, wire5923, n_n5020, wire898, n_n99, n_n186, n_n222, wire863, n_n4970, wire906, wire153, wire901, wire908, wire88, n_n4926, wire5343, wire5344, n_n261, n_n263, n_n108, wire70, n_n4826, wire899, n_n256, wire66, n_n4828, wire900, wire73, n_n4823, wire19738, wire44, n_n65, wire584, n_n12, n_n70, wire79, wire5268, wire5269, wire19742, wire63, n_n4815, n_n11, n_n4821, wire137, n_n4814, n_n4816, wire60, n_n4834, wire166, n_n4961, wire224, n_n95, n_n49, n_n96, n_n4967, wire613, wire99, wire41, wire614, wire5033, n_n4287, wire904, wire389, wire708, wire4196, wire20675, n_n4211, wire180, wire617, wire254, wire673, wire674, wire20677, wire20678, n_n4210, n_n4892, wire113, n_n4898, n_n4895, wire132, wire5035, wire5031, wire878, n_n48, wire51, n_n53, n_n4179, wire903, wire40, n_n31, n_n4168, n_n197, wire89, n_n4094, n_n47, wire67, n_n104, n_n4174, wire407, n_n247, wire457, n_n4153, n_n4154, wire456, wire4593, wire20257, wire20385, n_n3964, n_n93, n_n46, n_n896, n_n76, n_n29, wire49, wire460, wire160, n_n252, wire409, n_n4920, n_n4907, n_n253, wire82, n_n15, wire635, wire42, wire636, wire21065, wire21070, wire539, wire639, wire3904, wire20950, n_n3172, n_n4605, wire20955, wire20956, n_n3118, n_n26, wire80, wire640, n_n80, wire3758, wire21136, wire453, n_n3259, wire245, n_n3260, wire61, n_n3772, n_n3257, wire20959, wire20962, n_n3113, n_n223, n_n2860, n_n3255, wire814, wire3884, wire71, wire68, wire496, n_n179, wire55, wire57, wire806, n_n10, n_n100, wire19578, n_n1359, wire84, n_n3525, n_n107, wire62, n_n204, n_n16, wire3358, n_n4671, wire252, wire329, wire21442, wire21443, n_n2169, n_n66, wire164, wire985, wire3354, wire21529, wire21533, wire333, wire3541, wire3542, n_n171, n_n74, wire21367, n_n147, n_n94, n_n280, n_n32, n_n4165, n_n42, wire81, wire69, n_n4624, wire85, n_n1412, n_n135, n_n41, wire347, n_n18, wire123, wire100, wire992, n_n4858, n_n4864, wire102, n_n4635, wire22106, n_n4870, wire78, n_n1497, n_n1130, n_n22, wire897, wire19407, n_n4852, n_n103, n_n1490, wire140, wire346, wire998, wire22119, n_n1095, n_n1240, wire22129, wire22130, n_n1242, n_n1243, wire22142, n_n1505, wire22148, wire22149, wire56, n_n1542, n_n3827, n_n1536, wire22157, n_n1135, wire2638, wire22169, wire22176, n_n1097, wire368, n_n88, n_n1066, n_n270, wire114, n_n275, wire120, wire459, wire22648, n_n855, wire19457, n_n3870, wire2091, wire2092, wire22654, n_n772, n_n254, wire301, wire461, wire2008, wire19577, wire670, wire2001, wire2002, n_n269, n_n227, n_n207, n_n84, n_n142, n_n136, wire896, n_n278, n_n259, n_n149, n_n122, n_n112, n_n212, n_n30, n_n221, n_n7, n_n144, n_n50, n_n267, n_n87, n_n34, n_n28, n_n75, n_n21, n_n17, n_n236, n_n40, n_n102, n_n33, n_n78, n_n200, n_n64, n_n150, n_n25, n_n24, n_n27, n_n20, n_n97, n_n52, n_n71, n_n69, n_n14, n_n63, n_n199, n_n92, n_n98, n_n38, n_n109, wire384, wire19205, wire19239, wire5910, wire19207, wire19208, n_n5063, wire165, n_n4839, wire53, n_n4960, n_n4954, n_n4953, n_n4955, wire671, wire20705, wire20706, wire20710, wire469, n_n4073, wire475, n_n4068, n_n4069, wire77, n_n1363, wire184, n_n3324, n_n6504, n_n1633, n_n4923, wire21073, wire21074, n_n3130, wire686, wire825, wire20973, wire20974, wire20975, n_n3167, wire278, wire1018, wire20984, n_n3117, n_n3242, wire557, wire3754, n_n3757, wire739, wire20931, wire20933, wire20934, wire20936, wire20938, n_n3519, n_n3520, n_n148, n_n81, wire470, n_n3019, n_n2986, n_n3524, wire185, wire3310, wire21560, wire21561, wire21562, n_n2148, n_n19, n_n2272, wire3491, wire21417, n_n2126, wire135, wire264, wire1031, wire1030, wire466, wire3533, wire3534, wire21374, n_n2104, wire411, wire3344, wire3345, n_n2137, wire21381, n_n2110, wire21387, wire3518, wire21390, wire476, wire104, wire228, wire21842, n_n58, wire667, wire696, wire21686, wire21687, n_n1757, n_n3581, wire143, wire306, wire22079, n_n1215, wire514, n_n1628, wire52, n_n2732, n_n1624, wire247, wire83, wire1044, wire175, wire579, wire764, wire2542, wire2543, wire699, wire22020, n_n1320, wire376, wire2686, wire22121, n_n4124, wire629, n_n62, wire631, n_n6879, wire679, wire2672, wire2673, wire2665, wire22134, wire22135, wire22136, wire223, wire168, wire128, wire22605, n_n203, n_n1058, wire20149, n_n3604, n_n3610, wire697, wire1061, wire22610, wire22611, n_n771, wire516, wire1062, wire1997, wire22725, wire22727, n_n825, wire675, wire310, wire1064, wire1063, wire1990, wire22731, wire22734, n_n762, n_n13, wire2436, wire2437, n_n458, wire1066, wire22372, n_n374, wire486, wire658, n_n707, wire2410, wire22384, n_n462, wire1069, wire22383, n_n346, n_n43, n_n82, n_n68, n_n113, n_n86, n_n79, n_n36, n_n44, n_n73, wire19265, wire19266, wire19267, wire1071, wire277, n_n4924, wire255, n_n4871, n_n4838, wire19896, n_n4730, wire1076, wire1079, wire632, wire5368, wire5369, n_n4330, wire5361, wire5363, wire19671, n_n4806, n_n101, wire65, n_n1341, wire4602, n_n3974, n_n4090, wire462, wire464, wire20330, wire20331, wire1089, wire20340, wire20341, n_n3506, wire4302, wire455, wire485, wire76, n_n3781, wire676, wire21006, n_n3184, wire96, wire712, wire4472, wire20397, wire20400, wire20987, n_n3116, n_n35, n_n4922, n_n4921, n_n4076, n_n3768, wire484, wire21303, n_n2439, wire21603, n_n4912, n_n4916, wire327, wire1094, wire191, wire1096, wire1095, wire167, wire210, wire235, wire399, wire1097, wire436, wire1102, wire641, wire3145, wire21690, wire21691, n_n1756, wire50, wire645, wire2596, wire2597, wire22203, n_n1286, wire2593, wire2594, wire2516, wire22280, n_n1255, n_n6848, wire479, wire656, wire22286, wire22287, n_n1137, wire2879, wire21914, n_n1157, wire1112, n_n1295, n_n1641, wire22190, wire22193, n_n1151, wire1113, wire22185, n_n1102, n_n1284, wire22219, wire22220, wire807, n_n4675, n_n4681, n_n1604, wire497, wire22227, wire22228, n_n1101, n_n1298, wire22236, n_n1152, wire874, n_n1154, n_n3881, wire784, n_n1103, wire647, wire22785, wire356, wire22613, n_n850, wire335, wire1121, wire1120, wire2138, wire22616, n_n4628, wire727, n_n431, wire22409, wire22412, wire2374, wire22414, wire22415, wire22416, n_n429, wire22400, wire22401, n_n343, wire2361, wire2356, wire2353, wire2354, n_n363, n_n438, wire22446, n_n443, wire22454, wire22457, wire809, wire22459, wire1128, wire22463, wire22464, n_n143, n_n39, n_n77, n_n67, wire1131, wire19213, wire1130, wire5893, wire19215, wire19216, wire19217, wire1132, wire190, n_n4941, n_n4942, wire157, wire728, wire729, n_n5685, wire4889, wire20020, wire20021, wire4882, wire20023, wire20027, wire794, n_n4394, n_n4381, n_n3850, wire5587, wire473, wire124, n_n4929, wire212, wire250, wire1141, wire4166, wire20712, n_n4279, wire4569, wire4570, wire20273, n_n3978, n_n1346, n_n884, wire21228, n_n3908, n_n3778, n_n3229, wire740, n_n1555, wire626, n_n3791, wire478, wire20387, wire736, wire20392, n_n2815, n_n2982, wire349, wire483, wire876, wire20996, n_n3097, n_n3099, n_n3101, wire21063, n_n3103, wire21122, wire4694, wire4695, n_n3864, wire780, n_n2702, wire654, wire1372, n_n2398, wire1150, n_n2724, wire1156, wire3340, wire21537, wire21538, n_n2133, wire388, wire747, wire21540, wire21541, n_n2132, wire391, wire21549, wire330, wire241, wire1159, wire21425, n_n2129, wire21431, wire21432, n_n2274, wire1163, wire2780, wire2781, wire22022, n_n1217, n_n4687, wire22213, wire22214, wire2503, wire750, n_n1433, wire1171, wire22034, wire22040, wire22041, n_n1120, n_n1476, wire2777, wire589, wire2525, wire22270, wire2521, wire22277, n_n3843, wire19385, wire662, n_n1584, wire706, wire406, n_n952, wire1984, wire22736, n_n819, wire930, n_n5673, n_n59, n_n90, wire6020, wire19269, wire19270, wire19271, wire1181, wire1187, wire1186, wire5885, wire19223, wire19230, n_n5007, wire936, wire198, wire760, wire119, wire761, wire762, wire5076, wire19878, wire763, n_n4183, n_n4770, n_n4160, wire1279, n_n1645, wire767, wire21098, wire21101, n_n3309, wire463, wire20999, wire21003, wire21004, n_n3124, wire3852, wire681, wire21013, wire21014, n_n3123, n_n3122, wire21035, n_n3128, wire21054, n_n3587, wire770, wire771, n_n3132, n_n3133, wire21116, wire653, wire548, wire773, wire774, wire20056, wire1194, wire20060, n_n2665, wire1196, wire1195, wire1198, wire3005, wire3198, wire21660, wire21665, n_n1697, wire690, wire270, wire3186, wire21657, wire21673, n_n1753, wire3159, wire21683, n_n1703, wire21697, n_n1704, wire21699, wire21700, wire21701, wire21702, n_n1752, wire21648, wire21649, n_n1356, wire22043, wire22044, n_n1208, n_n639, wire694, wire869, wire22053, wire22054, n_n1121, n_n876, wire850, wire22775, wire22776, n_n790, wire743, wire232, wire22336, wire1213, wire22338, wire2463, wire22348, wire22351, wire642, wire351, wire22352, wire1217, wire19341, wire19284, wire19285, n_n5051, wire1223, wire19288, n_n5017, wire1226, wire5874, wire5875, wire19882, n_n4633, wire705, wire1231, wire20719, wire20720, wire20721, wire20722, n_n4218, n_n4214, n_n4255, wire20729, wire20733, n_n1370, wire5591, wire5592, wire309, wire571, wire737, wire20300, wire20301, wire20304, wire5510, wire5514, wire5515, wire20155, n_n3598, wire3800, wire21083, n_n3209, wire628, wire21105, n_n4644, n_n4636, wire4745, wire20131, wire21019, wire21027, wire21028, n_n4632, wire487, wire742, wire931, wire20362, wire20364, n_n2876, n_n3731, n_n1597, wire3595, wire3588, wire21318, wire271, wire472, wire21723, wire21724, n_n1788, wire21713, wire21714, wire21718, wire21719, n_n1715, wire1250, wire1249, wire1248, wire21729, wire21730, n_n1792, wire158, wire1251, wire21728, wire21739, n_n1690, n_n1440, wire300, n_n1173, wire2740, wire22064, n_n1210, n_n6820, wire1253, wire22765, wire22766, wire1254, wire320, wire22335, n_n370, wire276, wire182, wire405, wire22477, wire1259, wire2304, wire2305, wire2296, wire22483, wire22487, wire877, wire2277, wire22495, wire22496, n_n464, wire688, wire358, wire1261, wire22493, wire22494, wire22504, wire5988, n_n5048, wire315, wire1265, wire1264, wire326, wire19260, wire19261, wire19263, n_n4911, n_n3736, n_n1339, n_n3579, n_n4674, wire3830, wire3831, wire4492, wire20366, wire20367, n_n2875, wire3316, wire3317, n_n2145, wire226, wire21832, n_n1785, wire1291, wire1290, wire1289, wire2566, wire22231, wire22232, wire687, wire22066, wire22067, n_n1212, wire374, wire434, wire799, wire22075, wire22076, n_n1123, wire20755, wire229, n_n5664, wire793, wire22240, wire22241, wire22242, wire1307, wire22512, wire22513, wire1311, wire2258, wire624, wire233, wire22522, n_n408, wire22524, wire22527, wire19909, n_n4736, wire481, n_n4913, n_n4259, n_n4915, n_n4914, wire721, wire5589, wire20121, n_n4256, wire101, wire5011, wire5552, wire465, wire5613, n_n3786, n_n3782, wire723, wire19384, wire19440, n_n4676, n_n4686, wire1322, wire3764, wire21108, wire21109, wire21110, n_n3221, wire1323, wire21046, wire21047, wire298, n_n5675, wire1327, wire3303, wire21565, wire21566, n_n2146, wire429, wire263, wire1329, wire1330, wire21770, wire21771, wire21772, n_n1774, wire3032, wire3033, wire1333, wire22187, wire22188, wire1334, n_n3884, wire580, wire22796, wire22797, n_n809, wire1340, wire1343, wire1344, wire22363, wire408, wire933, wire414, wire357, wire22340, wire22533, wire1354, wire1357, wire1355, wire22537, wire419, wire19604, wire20344, n_n4146, wire20253, wire20254, n_n3925, wire21250, wire3707, wire3708, wire21188, n_n3930, wire3702, wire21190, wire21191, n_n3929, wire4587, wire20259, wire20262, wire20271, n_n3980, wire20282, n_n3920, wire4558, wire20287, n_n3922, wire4552, wire20293, wire4530, wire20310, wire20319, wire59, wire19582, wire4131, wire20756, n_n3486, wire20764, wire20765, n_n3403, n_n3372, wire225, n_n2713, wire5506, wire370, wire130, wire4789, wire20775, wire20782, n_n3371, wire19936, wire19914, n_n3397, wire788, wire21077, wire21081, wire20374, wire20376, wire1371, wire20381, wire20382, wire21389, n_n2158, wire1378, wire1377, n_n4682, wire21445, wire21446, n_n2172, wire482, wire1379, wire3452, wire21449, wire21453, n_n2093, wire86, n_n4666, wire1383, wire21462, wire21463, wire21470, wire425, wire657, wire2939, wire21857, n_n1804, wire448, wire2745, wire22061, n_n1092, wire1491, wire21935, n_n1108, wire1492, wire21941, wire519, wire22625, wire22626, wire22646, n_n742, wire139, wire776, wire22662, wire22663, wire22670, n_n744, n_n5679, wire321, wire331, wire19319, wire19320, wire1400, wire546, wire634, wire21257, wire21258, wire4089, wire4090, n_n3406, wire3698, wire21193, n_n3932, wire21200, wire21201, n_n3904, n_n3806, wire5780, wire19381, n_n3408, wire20793, n_n3374, wire20798, wire19400, wire19401, wire633, wire20804, n_n3362, wire4391, wire20403, n_n2817, wire4470, wire533, wire20412, wire20484, n_n2804, wire20553, wire4319, wire3292, wire21574, n_n2140, wire3370, wire21516, wire21517, n_n2099, wire281, wire338, wire858, wire1413, wire242, wire1416, n_n2097, wire3419, wire21482, wire21483, n_n2180, wire1423, n_n3770, wire21963, wire1424, wire22000, wire22007, wire587, wire4565, wire20275, wire3660, wire3661, wire21236, n_n3709, wire882, wire4453, wire20429, wire20430, wire20452, wire20469, wire20495, wire4360, wire20516, wire20541, wire20542, wire19408, wire693, wire3277, wire21590, n_n2154, wire3368, wire1450, wire1451, wire823, wire22087, wire22088, n_n1124, wire22095, n_n1093, wire381, wire152, wire21281, wire21089, wire21090, wire20573, wire20574, wire20575, wire20576, wire1463, n_n2808, wire20435, wire4435, wire20437, wire20442, wire20583, n_n2806, wire792, wire3272, wire21593, n_n2155, wire21596, n_n3751, wire380, wire1474, wire20457, wire395, wire20562, wire829, wire21379, wire1485, wire21572, wire21551, wire1486, wire343, wire21930, wire2019, wire22710, n_n834, n_n560, wire5834, wire5835, wire5843, wire5844, n_n5009, wire4478, wire716, wire4344, wire20532, wire20533, wire3287, wire21579, n_n1598, wire704, n_n3523, wire21975, wire1514, n_n1591, wire144, n_n618, wire1517, wire5550, wire5244, wire5245, wire19865, n_n4773, n_n4680, wire468, wire21609, wire1528, wire369, wire1530, n_n4489, n_n4677, wire371, wire1545, wire20192, wire20117, wire4655, wire20199, wire20200, wire20209, wire1552, wire19485, n_n3638, wire19398, n_n3624, wire19405, wire5734, wire19413, n_n3550, wire20862, n_n3380, wire5569, wire20836, n_n3417, wire4071, wire4073, wire20809, wire5725, wire5726, n_n2598, n_n2579, wire2975, wire2976, wire21827, wire21828, n_n1781, n_n785, wire22546, wire22547, wire22548, n_n413, wire471, wire22556, wire22557, wire22558, n_n359, wire5238, wire5239, wire19900, wire1575, n_n4685, wire19387, wire19495, wire19489, wire19490, wire5720, wire20865, wire20866, n_n3379, wire4042, n_n3393, wire20501, wire20502, n_n2633, wire5711, wire812, wire19770, n_n2580, wire1593, wire21668, wire21834, wire1594, n_n1713, wire195, wire21748, wire21749, wire1597, wire375, wire240, wire21746, wire1596, wire857, wire1599, wire494, wire1600, wire21766, wire21767, wire21769, n_n1691, wire862, wire895, wire855, wire856, wire1606, wire22778, n_n750, wire22561, wire22562, wire22565, wire20134, wire20119, wire20122, wire5439, wire609, wire5721, wire19784, wire19778, wire19787, n_n2578, wire19793, n_n2572, wire19798, wire19802, n_n2582, wire1627, n_n1773, wire21783, wire21784, wire21792, n_n1709, wire21794, wire1630, wire21799, n_n1688, wire3000, wire21808, n_n1706, wire21813, wire21814, wire21817, wire21825, n_n1687, wire2960, wire2961, wire21847, n_n1711, wire21855, wire22675, wire22676, wire1637, wire22678, wire275, wire262, wire887, wire1640, wire1639, wire1638, wire145, wire22687, wire1641, wire22685, wire22686, wire22693, wire1649, wire1647, wire19931, wire19946, wire19959, wire19953, wire19967, wire672, n_n3803, wire20141, wire20142, wire20224, n_n4551, wire19537, n_n3708, wire20228, wire20232, wire20872, wire3989, wire20881, wire3985, wire20882, wire20888, wire20889, n_n3385, wire20508, wire227, wire1662, wire1661, wire1664, wire20068, wire20073, wire1668, wire21888, wire21889, wire426, wire134, wire544, wire1669, wire22792, wire22793, n_n755, wire22803, wire22804, wire22809, n_n756, wire22814, wire403, wire1673, wire22451, wire1678, wire1677, wire1676, wire292, wire1682, wire1680, wire1679, wire1687, wire5758, wire19393, wire20897, wire20904, wire20905, n_n3383, wire1696, wire21652, wire379, wire2011, wire22714, wire22717, wire22744, wire22763, wire22822, wire1703, wire1707, wire1706, wire5671, wire19458, n_n3686, wire1717, wire236, wire74, wire424, wire1730, wire1733, wire1737, wire22403, wire22404, wire1740, wire19465, wire19466, wire19467, wire19523, wire1747, wire1753, wire1752, wire1755, wire20075, wire20076, n_n2671, wire20094, n_n2673, wire20104, n_n2659, wire2994, wire3018, wire3019, wire21786, wire1773, wire1772, wire1771, wire1776, wire1777, wire22829, wire22830, wire20153, wire20157, wire1786, wire3578, wire21675, wire21676, wire21677, wire21678, wire622, wire1794, wire22341, wire22572, wire22573, wire22581, n_n341, wire1797, wire1796, wire19565, wire19566, wire1803, wire21864, wire21865, wire21874, wire21877, wire20096, wire3576, wire3577, n_n2431, wire441, wire1814, wire1813, wire1825, wire20176, wire1829, wire3720, wire21168, wire3558, wire21352, wire362, wire1835, wire161, wire22835, wire22833, wire1836, wire1849, wire47, wire19575, wire87, wire110, wire288, wire148, wire187, wire196, wire197, wire214, wire215, wire220, wire230, wire231, wire243, wire246, wire256, wire274, wire19238, wire19253, wire287, wire291, wire304, wire305, wire311, wire325, wire328, wire342, wire345, wire348, wire352, wire361, wire397, wire413, wire428, wire431, wire433, wire435, wire437, wire444, wire1874, wire1918, wire962, wire965, wire968, wire971, wire1074, wire1101, wire1135, wire1182, wire1199, wire1225, wire1317, wire1501, wire1619, wire1792, wire22841, wire238, wire505, wire22816, wire529, wire543, wire550, wire564, wire22795, wire608, wire22772, wire22769, wire1970, wire22752, wire1971, wire22746, wire1976, wire1977, wire22730, wire22719, wire2012, wire2022, wire2023, wire2030, wire2034, wire22696, wire2035, wire2041, wire2059, wire2067, wire22664, wire2072, wire2081, wire22657, wire2082, wire2089, wire22650, wire2103, wire2104, wire22631, wire2122, wire2128, wire2129, wire2162, wire22598, wire22597, wire2170, wire2173, wire2174, wire2176, wire2183, wire2196, wire2200, wire2205, wire2206, wire2225, wire2235, wire2237, wire2239, wire22535, wire2240, wire2246, wire22519, wire22515, wire22516, wire2260, wire2263, wire22506, wire2264, wire2267, wire2268, wire2269, wire2291, wire22475, wire22471, wire2306, wire2311, wire2333, wire2336, wire2344, wire22436, wire22429, wire2364, wire22407, wire22408, wire2378, wire2392, wire2393, wire2398, wire22387, wire2403, wire2425, wire22376, wire2426, wire2427, wire22374, wire2428, wire2472, wire2473, wire2478, wire2486, wire2491, wire2495, wire22290, wire2507, wire2508, wire2520, wire22275, wire22276, wire2532, wire2533, wire2534, wire22259, wire2545, wire2560, wire2561, wire2571, wire2572, wire2581, wire2583, wire22206, wire22210, wire22211, wire2601, wire2602, wire2623, wire22170, wire2631, wire22162, wire2637, wire22167, wire22168, wire2640, wire2652, wire22139, wire2659, wire2676, wire2703, wire2708, wire2709, wire2725, wire2726, wire22058, wire22059, wire2774, wire22033, wire22024, wire2784, wire22001, wire2813, wire2814, wire2822, wire21979, wire21980, wire2825, wire2827, wire21971, wire2830, wire2831, wire2839, wire21953, wire21954, wire2842, wire2845, wire2864, wire2874, wire21913, wire2883, wire2885, wire2888, wire2889, wire2893, wire21892, wire2917, wire2918, wire2919, wire2920, wire2927, wire2928, wire2929, wire2942, wire2943, wire2952, wire2973, wire2974, wire21821, wire21805, wire21807, wire3003, wire3004, wire21789, wire3012, wire21785, wire3043, wire3045, wire3056, wire3065, wire3072, wire3080, wire3098, wire3106, wire3109, wire3120, wire3178, wire3179, wire3187, wire3190, wire21658, wire3203, wire21650, wire3211, wire3213, wire3214, wire3219, wire21642, wire3220, wire3221, wire21639, wire21640, wire3222, wire3228, wire3232, wire21584, wire21576, wire3296, wire3297, wire3324, wire21536, wire3375, wire3376, wire3382, wire3393, wire3400, wire3401, wire3402, wire3409, wire3413, wire3416, wire3440, wire21457, wire21458, wire3441, wire3442, wire3447, wire3451, wire3469, wire3470, wire3480, wire3499, wire3500, wire3520, wire21383, wire3544, wire3550, wire3551, wire3562, wire3563, wire3565, wire3584, wire3585, wire3627, wire21266, wire3629, wire3642, wire3653, wire3662, wire3674, wire3680, wire3681, wire3682, wire3688, wire3689, wire3712, wire3725, wire3726, wire3733, wire3736, wire3778, wire3790, wire3791, wire3821, wire3837, wire3843, wire21009, wire3896, wire3924, wire3931, wire20917, wire3946, wire3967, wire3968, wire3975, wire3976, wire20874, wire3988, wire20875, wire4004, wire4005, wire4016, wire20839, wire20840, wire4036, wire4044, wire4056, wire4062, wire4081, wire4100, wire4117, wire4120, wire4159, wire4170, wire4183, wire4202, wire20637, wire20638, wire4248, wire4267, wire4276, wire4281, wire20585, wire4285, wire4313, wire4330, wire20512, wire20513, wire20514, wire4373, wire4380, wire4409, wire4417, wire4418, wire4423, wire4463, wire20365, wire4506, wire4520, wire4551, wire4573, wire4574, wire4617, wire4618, wire20213, wire4636, wire4641, wire4656, wire20180, wire4690, wire4691, wire4711, wire4727, wire4750, wire20107, wire4766, wire4790, wire20089, wire20090, wire4800, wire20086, wire20087, wire4805, wire4807, wire4808, wire4817, wire4844, wire4845, wire4849, wire4856, wire4869, wire4870, wire4871, wire4890, wire4892, wire4896, wire4899, wire4900, wire4902, wire4905, wire4928, wire4939, wire4947, wire4974, wire5002, wire5012, wire5013, wire5014, wire5023, wire5036, wire5047, wire5048, wire5054, wire5059, wire5091, wire5099, wire19848, wire5138, wire5144, wire5160, wire19814, wire5161, wire5184, wire5205, wire5215, wire5219, wire5228, wire5240, wire5241, wire5242, wire5243, wire5262, wire19713, wire19714, wire5299, wire5327, wire5328, wire19683, wire5357, wire5362, wire19668, wire5371, wire5372, wire5390, wire5400, wire5411, wire5412, wire5413, wire5426, wire5430, wire5441, wire5442, wire5445, wire19605, wire5472, wire5494, wire5509, wire19556, wire19548, wire5516, wire5517, wire5544, wire5564, wire5565, wire5577, wire5588, wire5590, wire5596, wire5606, wire19491, wire5617, wire5625, wire5626, wire5640, wire5642, wire5643, wire5650, wire5651, wire5656, wire19469, wire5657, wire5660, wire5661, wire5681, wire5699, wire5709, wire5743, wire5749, wire5754, wire5775, wire5778, wire5797, wire5812, wire5813, wire19350, wire5824, wire19344, wire19347, wire19348, wire19342, wire19237, wire5848, wire19334, wire5850, wire19332, wire5854, wire19329, wire19330, wire5861, wire5862, wire19244, wire5863, wire19313, wire5877, wire5878, wire5879, wire5880, wire19220, wire19221, wire19211, wire5900, wire19197, wire19198, wire19252, wire5953, wire5955, wire5973, wire5985, wire19291, wire5990, wire5999, wire6008, wire6014, wire19274, wire19275, wire6009, wire19212, wire19228, wire19233, wire19243, wire19250, wire19254, wire19255, wire19264, wire19278, wire19286, wire19287, wire19297, wire19299, wire19300, wire19301, wire19302, wire19303, wire19305, wire19307, wire19311, wire19318, wire19323, wire19326, wire19327, wire19331, wire19339, wire19345, wire19353, wire19354, wire19355, wire19363, wire19364, wire19369, wire19377, wire19379, wire19383, wire19394, wire19402, wire19422, wire19442, wire19443, wire19447, wire19452, wire19453, wire19460, wire19461, wire19470, wire19475, wire19478, wire19499, wire19502, wire19515, wire19516, wire19519, wire19520, wire19522, wire19526, wire19528, wire19534, wire19539, wire19541, wire19549, wire19550, wire19559, wire19568, wire19571, wire19588, wire19599, wire19609, wire19617, wire19619, wire19620, wire19628, wire19631, wire19632, wire19633, wire19636, wire19642, wire19644, wire19645, wire19665, wire19669, wire19696, wire19701, wire19703, wire19704, wire19705, wire19706, wire19707, wire19709, wire19710, wire19720, wire19724, wire19725, wire19728, wire19730, wire19732, wire19735, wire19747, wire19755, wire19757, wire19759, wire19761, wire19780, wire19791, wire19807, wire19808, wire19810, wire19812, wire19821, wire19825, wire19826, wire19830, wire19837, wire19842, wire19843, wire19854, wire19857, wire19859, wire19862, wire19867, wire19868, wire19872, wire19888, wire19904, wire19906, wire19916, wire19918, wire19919, wire19921, wire19925, wire19926, wire19927, wire19928, wire19938, wire19941, wire19943, wire19944, wire19952, wire19958, wire19965, wire19971, wire19973, wire19974, wire19977, wire19984, wire19986, wire19987, wire19996, wire19997, wire19999, wire20000, wire20011, wire20015, wire20016, wire20017, wire20028, wire20030, wire20031, wire20038, wire20041, wire20042, wire20045, wire20047, wire20048, wire20054, wire20055, wire20066, wire20070, wire20072, wire20081, wire20084, wire20088, wire20099, wire20100, wire20101, wire20108, wire20111, wire20113, wire20137, wire20174, wire20186, wire20188, wire20190, wire20191, wire20193, wire20203, wire20206, wire20212, wire20216, wire20227, wire20236, wire20238, wire20248, wire20264, wire20265, wire20268, wire20269, wire20277, wire20278, wire20279, wire20285, wire20299, wire20307, wire20323, wire20324, wire20325, wire20334, wire20336, wire20337, wire20343, wire20346, wire20347, wire20349, wire20350, wire20356, wire20369, wire20370, wire20371, wire20379, wire20390, wire20401, wire20404, wire20408, wire20409, wire20418, wire20419, wire20422, wire20424, wire20425, wire20434, wire20438, wire20444, wire20445, wire20449, wire20450, wire20455, wire20460, wire20461, wire20463, wire20474, wire20479, wire20480, wire20486, wire20492, wire20499, wire20506, wire20510, wire20519, wire20520, wire20522, wire20525, wire20527, wire20536, wire20537, wire20540, wire20549, wire20581, wire20590, wire20593, wire20600, wire20604, wire20606, wire20608, wire20609, wire20620, wire20622, wire20624, wire20633, wire20636, wire20641, wire20642, wire20643, wire20646, wire20655, wire20668, wire20682, wire20683, wire20686, wire20689, wire20692, wire20694, wire20695, wire20696, wire20699, wire20701, wire20703, wire20704, wire20711, wire20714, wire20716, wire20728, wire20737, wire20739, wire20742, wire20745, wire20746, wire20748, wire20751, wire20758, wire20759, wire20760, wire20767, wire20769, wire20772, wire20776, wire20779, wire20784, wire20800, wire20802, wire20814, wire20817, wire20820, wire20824, wire20826, wire20827, wire20831, wire20832, wire20833, wire20842, wire20847, wire20851, wire20853, wire20854, wire20856, wire20876, wire20883, wire20894, wire20895, wire20898, wire20899, wire20900, wire20907, wire20908, wire20909, wire20912, wire20942, wire20952, wire20967, wire20981, wire20982, wire20988, wire20989, wire20993, wire20994, wire20998, wire21010, wire21017, wire21021, wire21022, wire21023, wire21030, wire21042, wire21043, wire21049, wire21051, wire21057, wire21059, wire21061, wire21066, wire21072, wire21076, wire21085, wire21092, wire21093, wire21113, wire21114, wire21120, wire21125, wire21129, wire21143, wire21146, wire21151, wire21153, wire21157, wire21159, wire21160, wire21163, wire21164, wire21165, wire21169, wire21170, wire21173, wire21175, wire21180, wire21183, wire21195, wire21196, wire21197, wire21206, wire21208, wire21225, wire21233, wire21238, wire21248, wire21252, wire21253, wire21260, wire21261, wire21263, wire21268, wire21269, wire21271, wire21288, wire21298, wire21299, wire21329, wire21337, wire21356, wire21372, wire21385, wire21394, wire21403, wire21404, wire21408, wire21409, wire21415, wire21426, wire21427, wire21428, wire21434, wire21435, wire21438, wire21448, wire21455, wire21459, wire21466, wire21467, wire21474, wire21478, wire21479, wire21486, wire21487, wire21488, wire21490, wire21491, wire21493, wire21494, wire21497, wire21499, wire21500, wire21501, wire21505, wire21506, wire21521, wire21522, wire21525, wire21530, wire21531, wire21544, wire21545, wire21546, wire21569, wire21614, wire21626, wire21627, wire21628, wire21633, wire21647, wire21651, wire21655, wire21662, wire21663, wire21670, wire21671, wire21681, wire21694, wire21695, wire21709, wire21715, wire21716, wire21721, wire21726, wire21732, wire21733, wire21735, wire21737, wire21741, wire21742, wire21743, wire21744, wire21751, wire21752, wire21753, wire21756, wire21757, wire21759, wire21760, wire21761, wire21762, wire21764, wire21780, wire21781, wire21790, wire21811, wire21815, wire21844, wire21845, wire21849, wire21850, wire21853, wire21859, wire21860, wire21861, wire21862, wire21872, wire21884, wire21902, wire21910, wire21912, wire21918, wire21920, wire21922, wire21923, wire21925, wire21926, wire21927, wire21928, wire21933, wire21948, wire21950, wire21956, wire21962, wire21968, wire21969, wire21970, wire21973, wire21977, wire21981, wire21982, wire21987, wire21988, wire21991, wire21992, wire21993, wire22002, wire22005, wire22010, wire22012, wire22035, wire22039, wire22047, wire22048, wire22050, wire22052, wire22070, wire22071, wire22081, wire22082, wire22083, wire22084, wire22090, wire22093, wire22097, wire22101, wire22117, wire22124, wire22125, wire22126, wire22140, wire22154, wire22160, wire22164, wire22174, wire22181, wire22208, wire22217, wire22255, wire22262, wire22273, wire22282, wire22302, wire22308, wire22312, wire22314, wire22317, wire22322, wire22326, wire22327, wire22328, wire22330, wire22332, wire22337, wire22346, wire22356, wire22366, wire22369, wire22370, wire22378, wire22379, wire22380, wire22389, wire22395, wire22399, wire22443, wire22449, wire22456, wire22461, wire22489, wire22490, wire22491, wire22492, wire22502, wire22511, wire22518, wire22523, wire22532, wire22538, wire22539, wire22541, wire22543, wire22551, wire22552, wire22566, wire22567, wire22570, wire22571, wire22574, wire22575, wire22576, wire22578, wire22590, wire22593, wire22596, wire22600, wire22606, wire22618, wire22633, wire22635, wire22636, wire22637, wire22638, wire22639, wire22640, wire22642, wire22643, wire22651, wire22652, wire22658, wire22659, wire22665, wire22667, wire22668, wire22672, wire22680, wire22681, wire22683, wire22684, wire22689, wire22692, wire22695, wire22698, wire22700, wire22701, wire22703, wire22704, wire22708, wire22709, wire22712, wire22720, wire22732, wire22742, wire22780, wire22786, wire22787, wire22788, wire22801, wire22805, wire22806, wire22820, wire22837, wire22843, wire22844, _61, _92, _140, _143, _231, _235, _237, _290, _339, _350, _358, _361, _367, _370, _373, _379, _380, _382, _385, _399, _455, _492, _506, _560, _561, _562, _567, _605, _608, _614, _617, _632, _635, _654, _655, _675, _696, _699, _702, _703, _705, _706, _710, _713, _716, _719, _720, _721, _725, _726, _727, _728, _774, _788, _793, _796, _801, _808, _817, _822, _830, _833, _834, _848, _897, _899, _900, _945, _946, _995, _998, _1010, _1051, _1054, _1064, _1067, _1102, _1166, _1167, _1168, _1194, _1195, _1196, _1203, _1204, _1205, _1206, _1209, _1215, _1216, _1248, _1251, _1254, _1261, _1262, _1263, _1266, _1292, _1305, _1306, _1338, _1340, _1346, _1349, _1354, _1357, _1360, _1363, _1372, _1394, _1427, _1428, _1429, _1430, _1433, _1473, _1497, _1498, _1509, _1510, _1512, _1515, _1516, _1518, _1526, _1527, _1528, _1531, _1534, _1535, _1537, _1540, _1580, _1583, _1584, _1588, _1591, _1592, _1593, _1596, _1599, _1602, _1614, _1617, _1626, _1652, _1655, _1673, _1676, _1683, _1686, _1718, _1719, _1720, _1723, _1729, _1730, _1731, _1737, _1743, _1744, _1760, _1796, _1797, _1801, _1807, _1815, _1816, _1817, _1832, _1835, _1843, _1853, _1861, _1889, _1892, _1895, _1896, _1898, _1903, _1906, _1909, _1934, _1952, _1966, _1967, _1968, _1997, _1998, _2137, _2138, _2139, _2140, _2145, _2146, _2147, _2150, _2215, _2220, _2223, _2224, _2225, _2230, _2235, _2236, _2237, _2240, _2306, _2307, _2308, _2314, _2337, _2346, _2347, _2348, _2403, _2404, _2412, _2448, _2449, _2458, _2459, _2463, _2474, _2475, _2476, _2477, _2478, _2483, _2486, _2487, _2488, _2498, _2503, _2517, _2557, _2558, _2611, _2630, _2633, _2656, _2657, _2677, _2711, _2716, _2719, _2720, _2727, _2728, _2732, _2733, _2741, _2760, _2761, _2766, _2793, _2854, _2888, _2891, _2946, _2959, _2960, _2961, _2962, _2965, _2976, _2979, _2982, _2983, _2984, _2985, _2992, _2993, _3000, _3001, _3002, _3003, _3006, _3007, _3008, _3011, _3012, _3013, _3014, _3016, _3021, _3022, _3023, _3027, _3028, _3035, _3036, _3037, _3038, _3041, _3042, _3043, _3044, _3058, _3064, _3067, _3070, _3077, _3078, _3082, _3094, _3095, _3096, _3101, _3102, _3103, _3106, _3107, _3108, _3124, _3132, _3173, _3174, _3175, _3178, _3179, _3180, _3181, _3182, _3187, _3188, _3189, _3190, _3195, _3196, _3197, _3206, _3211, _3216, _3217, _3218, _3222, _3223, _3235, _3236, _3260, _3263, _3271, _3294, _3295, _3296, _3300, _3311, _3314, _3319, _3320, _3324, _3327, _3328, _3329, _3330, _3333, _3343, _3344, _3358, _3384, _3396, _3400, _3408, _3411, _3414, _3423, _3424, _3430, _3443, _3444, _3446, _3449, _3452, _3472, _3498, _3503, _3512, _3529, _3547, _3550, _3566, _3567, _3570, _3589, _3597, _3598, _3599, _3602, _3628, _3629, _3636, _3674, _3675, _3679, _3680, _3692, _3695, _3708, _3718, _3719, _3723, _3724, _3786, _3787, _3833, _3834, _3852, _3878, _3896, _3920, _3973, _3979, _3980, _3988, _3991, _4005, _4006, _4007, _4008, _4013, _4014, _4015, _4018, _4028, _4031, _4032, _4039, _4040, _4041, _4044, _4045, _4046, _4139, _4147, _4148, _4149, _4155, _4156, _4160, _4161, _4165, _4166, _4167, _4170, _4177, _4180, _4189, _4209, _4210, _4219, _4220, _4221, _4226, _4249, _4252, _4260, _4263, _4264, _4271, _4272, _4273, _4274, _4277, _4295, _4296, _4297, _4300, _4301, _4302, _4310, _4311, _4312, _4313, _4318, _4324, _4342, _4348, _4349, _4357, _4362, _4365, _4366, _4370, _4371, _4376, _4377, _4378, _4385, _4390, _4401, _4412, _4413, _4414, _4426, _4429, _4432, _4456, _4457, _4469, _4485, _4514, _4559, _4567, _4574, _4577, _4582, _4585, _4596, _4599, _4600, _4605, _4609, _4610, _4614, _4615, _4622, _4631, _4635, _4643, _4653, _4675, _4681, _4687, _4688, _4694, _4701, _4702, _4706, _4769, _4771, _4775, _4777, _4778, _4782, _4792, _4795, _4798, _4799, _4811, _4814, _4861, _4868, _4878, _4881, _4901, _4906, _4907, _4908, _4909, _4920, _4943, _4944, _4977, _5028, _5079, _5101, _5118, _5119, _5135, _5145, _5150, _5153, _5158, _5164, _5165, _5173, _5174, _5179, _5183, _5218, _5219, _5225, _5227, _5230, _5231, _5239, _5241, _5244, _5274, _5282, _5283, _5288, _5302, _5303, _5309, _5310, _5341, _5346, _5347, _5355, _5357, _5359, _5362, _5365, _5376, _5377, _5378, _5381, _5389, _5392, _5399, _5405, _5408, _5422, _5425, _5426, _5435, _5446, _5457, _5458, _5459, _5462, _5470, _5480, _5481, _5485, _5501, _5502, _5503, _5552, _5559, _5578, _5593, _5604, _5617, _5618, _5619, _5620, _5624, _5751, _5752, _5753, _5756, _5776, _5783, _5807, _5810, _5820, _5823, _5889, _5900, _5901, _5905, _5910, _5922, _5925, _5932, _5940, _5943, _5967, _5968, _5980, _5981, _5982, _5993, _5996, _6010, _6034, _6055, _6058, _6069, _6070, _6077, _6157, _6160, _6161, _6176, _6177, _6189, _6192, _6205, _6208, _6220, _6221, _6235, _6236, _6237, _6238, _6252, _6280, _6287, _6294, _6298, _6301, _6319, _6363, _6387, _6408, _6443, _6447, _6448, _6461, _6474, _6483, _6484, _6540, _6592, _6597, _6700, _6703, _6706, _6708, _6730, _6812, _6813, _6821, _6822, _6824, _6827, _6830, _6836, _6837, _6838, _6843, _6848, _6849, _6857, _6858, _6859, _6865, _6866, _6868, _6927, _6928, _6930, _6970, _6977, _6984, _6995, _6996, _6997, _6998, _34535, _34536, _34537, _34544, _34546, _34548, _34549, _34551, _34558, _34559, _34563, _34565, _34567, _34575, _34576, _34580, _34581, _34582, _34583, _34585, _34586, _34594, _34606, _34625, _34626, _34627, _34637, _34638, _34639, _34642, _34644, _34645, _34685, _34687, _34692, _34695, _34696, _34697, _34698, _34702, _34703, _34708, _34710, _34711, _34713, _34715, _34720, _34722, _34724, _34730, _34738, _34748, _34780, _34797, _34819, _34822, _34827, _34834, _34842, _34843, _34860, _34908, _34910, _34914, _34919, _34942, _34949, _34950, _34952, _34953, _34954, _34956, _34957, _34985, _34990, _35004, _35011, _35013, _35014, _35030, _35033, _35034, _35035, _35036, _35037, _35039, _35040, _35042, _35043, _35044, _35046, _35049, _35051, _35052, _35053, _35054, _35056, _35058, _35064, _35065, _35071, _35074, _35076, _35077, _35079, _35084, _35085, _35086, _35087, _35091, _35097, _35099, _35101, _35103, _35109, _35110, _35111, _35112, _35114, _35115, _35116, _35118, _35120, _35124, _35125, _35129, _35131, _35137, _35139, _35141, _35142, _35143, _35148, _35150, _35151, _35153, _35154, _35160, _35163, _35164, _35165, _35167, _35172, _35174, _35176, _35178, _35186, _35190, _35208, _35212, _35213, _35218, _35219, _35235, _35236, _35255, _35257, _35258, _35290, _35306, _35339, _35341, _35343, _35346, _35352, _35354, _35356, _35357, _35358, _35359, _35366, _35368, _35370, _35372, _35376, _35377, _35379, _35381, _35382, _35384, _35389, _35391, _35392, _35394, _35396, _35400, _35412, _35414, _35418, _35420, _35422, _35425, _35427, _35428, _35444, _35446, _35454, _35456, _35464, _35468, _35470, _35472, _35476, _35478, _35480, _35484, _35485, _35487, _35494, _35498, _35499, _35500, _35502, _35504, _35505, _35523, _35524, _35527, _35528, _35529, _35530, _35531, _35532, _35536, _35537, _35539, _35544, _35562, _35563, _35565, _35566, _35567, _35572, _35577, _35579, _35588, _35592, _35600, _35601, _35603, _35613, _35622, _35623, _35626, _35628, _35629, _35630, _35635, _35639, _35640, _35644, _35646, _35648, _35651, _35652, _35661, _35685, _35686, _35693, _35695, _35700, _35702, _35703, _35705, _35706, _35709, _35711, _35712, _35714, _35716, _35719, _35721, _35722, _35724, _35745, _35748, _35749, _35750, _35752, _35754, _35763, _35769, _35772, _35773, _35815, _35820, _35831, _35833, _35835, _35836, _35837, _35855, _35873, _35875, _35876, _35878, _35880, _35881, _35882, _35883, _35884, _35893, _35897, _35934, _35938, _35941, _35943, _35946, _35947, _35948, _35949, _35950, _35951, _35953, _35954, _35956, _35959, _35961, _35962, _35964, _35996, _35998, _35999, _36001, _36002, _36030, _36035, _36055, _36064, _36066, _36068, _36083, _36085, _36086, _36087, _36090, _36091, _36092, _36093, _36095, _36096, _36098, _36099, _36101, _36107, _36112, _36113, _36115, _36116, _36121, _36122, _36137, _36138, _36139, _36140, _36143, _36144, _36149, _36150, _36156, _36157, _36159, _36161, _36165, _36168, _36176, _36179, _36180, _36184, _36190, _36192, _36193, _36195, _36198, _36202, _36203, _36205, _36210, _36212, _36215, _36218, _36219, _36222, _36224, _36227, _36229, _36231, _36234, _36235, _36238, _36242, _36244, _36245, _36249, _36250, _36253, _36255, _36256, _36264, _36265, _36267, _36270, _36273, _36275, _36277, _36282, _36285, _36286, _36289, _36291, _36293, _36297, _36298, _36304, _36308, _36311, _36312, _36315, _36317, _36319, _36324, _36330, _36331, _36334, _36335, _36337, _36339, _36341, _36343, _36360, _36375, _36377, _36380, _36382, _36383, _36392, _36393, _36396, _36404, _36405, _36410, _36417, _36421, _36424, _36426, _36428, _36430, _36442, _36443, _36448, _36450, _36453, _36457, _36461, _36467, _36469, _36474, _36475, _36476, _36480, _36482, _36483, _36487, _36488, _36489, _36491, _36495, _36501, _36502, _36506, _36508, _36510, _36515, _36518, _36525, _36536, _36542, _36544, _36548, _36550, _36555, _36558, _36563, _36585, _36611, _36614, _36616, _36619, _36620, _36682, _36683, _36687, _36698, _36699, _36705, _36714, _36783, _36786, _36788, _36790, _36797, _36803, _36807, _36808, _36810, _36813, _36817, _36818, _36821, _36824, _36825, _36826, _36833, _36844, _36856, _36865, _36876, _36878, _36881, _36887, _36888, _36889, _36890, _36894, _36895, _36909, _36912, _36916, _36947, _36950, _36951, _36952, _36954, _36957, _36958, _36959, _36964, _36967, _36969, _36971, _36972, _36973, _36974, _36975, _36977, _36982, _36984, _36986, _36988, _36993, _36995, _37000, _37002, _37003, _37004, _37013, _37014, _37022, _37024, _37026, _37027, _37030, _37032, _37035, _37037, _37042, _37043, _37044, _37046, _37047, _37050, _37057, _37063, _37064, _37066, _37068, _37070, _37072, _37074, _37076, _37077, _37084, _37086, _37087, _37089, _37091, _37093, _37095, _37097, _37099, _37104, _37105, _37106, _37108, _37110, _37116, _37128, _37130, _37140, _37141, _37143, _37148, _37155, _37158, _37160, _37161, _37163, _37168, _37170, _37178, _37180, _37189, _37191, _37204, _37208, _37209, _37211, _37215, _37220, _37222, _37224, _37226, _37227, _37228, _37230, _37231, _37244, _37247, _37253, _37256, _37263, _37273, _37275, _37277, _37280, _37284, _37285, _37286, _37291, _37296, _37297, _37298, _37300, _37303, _37304, _37314, _37316, _37317, _37320, _37321, _37322, _37323, _37326, _37333, _37335, _37340, _37341, _37346, _37348, _37350, _37351, _37352, _37358, _37360, _37361, _37363, _37367, _37370, _37373, _37375, _37376, _37378, _37379, _37380, _37381, _37382, _37390, _37396, _37398, _37406, _37407, _37409, _37411, _37415, _37416, _37422, _37424, _37426, _37428, _37429, _37432, _37433, _37435, _37438, _37442, _37444, _37445, _37448, _37463, _37464, _37469, _37480, _37495, _37496, _37497, _37499, _37508, _37509, _37511, _37516, _37517, _37520, _37521, _37522, _37523, _37525, _37527, _37530, _37532, _37535, _37539, _37544, _37546, _37548, _37550, _37552, _37560, _37562, _37565, _37568, _37570, _37576, _37580, _37619, _37630, _37633, _37639, _37643, _37645, _37646, _37648, _37657, _37661, _37666, _37673, _37686, _37688, _37689, _37701, _37703, _37710, _37712, _37716, _37722, _37733, _37738, _37743, _37750, _37751, _37753, _37755, _37762, _37764, _37766, _37772, _37776, _37777, _37791, _37792, _37796, _37825, _37826, _37827, _37828, _37830, _37833, _37834, _37840, _37841, _37846, _37848, _37849, _37852, _37859, _37860, _37862, _37876, _37878, _37898, _37899, _37901, _37905, _37907, _37910, _37915, _37919, _37920, _37922, _37925, _37931, _37932, _37934, _37936, _37951, _37961, _37967, _37968, _37969, _37976, _37977, _37989, _37993, _37994, _38006, _38007, _38010, _38014, _38018, _38020, _38025, _38049, _38050, _38057, _38062, _38063, _38067, _38069, _38073, _38082, _38083, _38087, _38093, _38097, _38103, _38106, _38107, _38108, _38109, _38118, _38123, _38125, _38131, _38132, _38136, _38137, _38138, _38140, _38141, _38142, _38151, _38155, _38156, _38157, _38161, _38164, _38165, _38167, _38169, _38171, _38174, _38178, _38183, _38186, _38187, _38189, _38192, _38195, _38196, _38202, _38208, _38211, _38238, _38244, _38245, _38248, _38249, _38251, _38254, _38256, _38258, _38260, _38262, _38263, _38266, _38268, _38272, _38273, _38274, _38277, _38285, _38287, _38289, _38291, _38294, _38296, _38299, _38302, _38305, _38311, _38313, _38315, _38317, _38319, _38320, _38323, _38325, _38328, _38330, _38335, _38339, _38343, _38345, _38348, _38354, _38355, _38357, _38361, _38365, _38367, _38368, _38369, _38370, _38371, _38372, _38374, _38379, _38380, _38381, _38386, _38390, _38392, _38394, _38395, _38398, _38399, _38403, _38404, _38405, _38408, _38409, _38411, _38413, _38418, _38419, _38421, _38423, _38426, _38430, _38432, _38436, _38437, _38439, _38442, _38444, _38448, _38451, _38452, _38462, _38467, _38468, _38469, _38483, _38485, _38513, _38522, _38545, _38550, _38551, _38556, _38558, _38613, _38614, _38625, _38635, _38636, _38637, _38639, _38640, _38643, _38656, _38658, _38663, _38665, _38666, _38668, _38670, _38673, _38679, _38681, _38691, _38699, _38703, _38708, _38713, _38722, _38723, _38724, _38725, _38726, _38727, _38729, _38730, _38732, _38733, _38734, _38740, _38741, _38748, _38750, _38769, _38770, _38772, _38785, _38788, _38789, _38794, _38804, _38805, _38806, _38809, _38844, _38846, _38848, _38853, _38854, _38855, _38857, _38858, _38860, _38862, _38867, _38870, _38872, _38874, _38877, _38880, _38881, _38882, _38883, _38885, _38891, _38892, _38897, _38898, _38900, _38902, _38906, _38907, _38930, _38932, _38941, _38942, _38943, _38945, _38957, _38958, _38965, _38966, _38968, _38969, _38971, _38972, _38973, _38978, _38979, _38984, _38986, _39001, _39002, _39005, _39006, _39007, _39009, _39010, _39011, _39044, _39048, _39051, _39052, _39053, _39055, _39057, _39059, _39063, _39067, _39072, _39073, _39078, _39081, _39084, _39085, _39091, _39094, _39095, _39096, _39097, _39100, _39109, _39113, _39114, _39115, _39118, _39122, _39131, _39255, _39273, _39274, _39275, _39283, _39286, _39296, _39307, _39309, _39322, _39332, _39334, _39337, _39338, _39340, _39341, _39346, _39347, _39348, _39350, _39351, _39356, _39359, _39360, _39363, _39369, _39370, _39372, _39375, _39379, _39382, _39384, _39387, _39389, _39396, _39398, _39406, _39412, _39425, _39426, _39427, _39432, _39441, _39449, _39450, _39461, _39470, _39479, _39486, _39495, _39502, _39514, _39526, _39528, _39529, _39530, _39534, _39536, _39537, _39540, _39542, _39543, _39546, _39552, _39553, _39554, _39555, _39556, _39565, _39566, _39571, _39573, _39574, _39576, _39578, _39580, _39582, _39584, _39590, _39594, _39596, _39600, _39601, _39632, _39633, _39645, _39646, _39651, _39653, _39657, _39664, _39670, _39673, _39674, _39676, _39683, _39684, _39690, _39702, _39703, _39704, _39707, _39708, _39722, _39740, _39743, _39744, _39746, _39749, _39750, _39753, _39754, _39758, _39759, _39772, _39785, _39786, _39788, _39793, _39796, _39801, _39803, _39805, _39807, _39809, _39811, _39816, _39817, _39839, _39848, _39853, _39860, _39861, _39878, _39888, _39890, _39891, _39892, _39893, _39897, _39902, _39903, _39906, _39908, _39925, _39929, _39934, _39937, _39950, _39951, _39957, _39959, _39961, _39962, _40013, _40015, _40016, _40037, _40041, _40056, _40059, _40065, _40066, _40067, _40068, _40069, _40070, _40071, _40072, _40078, _40080, _40086, _40103, _40109, _40110, _40111, _40115, _40124, _40125, _40133, _40134, _40140, _40142, _40160, _40161, _40165, _40166, _40169, _40173, _40183, _40190, _40195, _40198, _40200, _40201, _40205, _40208, _40217, _40218, _40226, _40229, _40232, _40234, _40239, _40242, _40245, _40246, _40248, _40249, _40250, _40252, _40253, _40254, _40255, _40258, _40259, _40262, _40264, _40265, _40266, _40268, _40269, _40272, _40274, _40275, _40276, _40288, _40294, _40307, _40308, _40311, _40313, _40322, _40330, _40336, _40337, _40338, _40340, _40342, _40345, _40347, _40371, _40373, _40375, _40381, _40385, _40391, _40392, _40393, _40394, _40395, _40397, _40404, _40405, _40407, _40408, _40410, _40411, _40412, _40413, _40414, _40416, _40418, _40420, _40422, _40425, _40441, _40442, _40472, _40474, _40517, _40518, _40536, _40538, _40544, _40546, _40548, _40564, _40565, _40568, _40573, _40584, _40602, _40604, _40607, _40618, _40620, _40633, _40648, _40649, _40657, _40658, _40660, _40671, _40672, _40675, _40676, _40678, _40699, _40701, _40706, _40712, _40713, _40728, _40773, _40784, _40796, _40807, _40808, _40811, _40812, _40820, _40828, _40832, _40833, _40836, _40857, _40858, _40859;

assign o_1_ = ( wire590 ) | ( wire19306 ) | ( _34942 ) | ( _35011 ) ;
 assign o_19_ = ( n_n5231 ) | ( n_n3621 ) | ( wire19592 ) | ( wire19593 ) ;
 assign o_2_ = ( wire590 ) | ( wire19306 ) | ( _34942 ) | ( _35750 ) ;
 assign o_0_ = ( wire19622 ) | ( wire590 ) | ( wire19306 ) | ( _34942 ) ;
 assign o_29_ = ( wire19648 ) | ( wire590 ) | ( wire19306 ) | ( _34942 ) ;
 assign o_39_ = ( wire590 ) | ( wire19306 ) | ( _34942 ) | ( _35875 ) ;
 assign o_38_ = ( wire590 ) | ( wire19306 ) | ( _34942 ) | ( _35878 ) ;
 assign o_25_ = ( n_n5231 ) | ( wire19766 ) | ( n_n4307 ) | ( _36068 ) ;
 assign o_12_ = ( wire19822 ) | ( wire590 ) | ( wire19306 ) | ( _34942 ) ;
 assign o_37_ = ( wire590 ) | ( wire19306 ) | ( _34942 ) | ( _36335 ) ;
 assign o_26_ = ( wire590 ) | ( wire19306 ) | ( _34942 ) | ( _36375 ) ;
 assign o_11_ = ( wire590 ) | ( wire19306 ) | ( _34942 ) | ( _36393 ) ;
 assign o_36_ = ( n_n5231 ) | ( n_n4718 ) | ( wire19989 ) | ( wire19990 ) ;
 assign o_27_ = ( wire590 ) | ( wire19306 ) | ( _5079 ) | ( _34942 ) ;
 assign o_14_ = ( wire590 ) | ( wire19306 ) | ( _34942 ) | ( _36611 ) ;
 assign o_35_ = ( wire590 ) | ( wire19306 ) | ( _34942 ) | ( _36620 ) ;
 assign o_28_ = ( n_n5224 ) | ( wire590 ) | ( wire19306 ) | ( _34942 ) ;
 assign o_13_ = ( n_n5231 ) | ( wire20115 ) | ( _36865 ) ;
 assign o_34_ = ( n_n5231 ) | ( wire20245 ) | ( n_n4535 ) | ( _36950 ) ;
 assign o_21_ = ( wire20355 ) | ( wire590 ) | ( wire19306 ) | ( _34942 ) ;
 assign o_16_ = ( n_n5231 ) | ( n_n2789 ) | ( n_n2795 ) | ( wire20625 ) ;
 assign o_33_ = ( wire590 ) | ( wire19306 ) | ( _34942 ) | ( _37633 ) ;
 assign o_22_ = ( wire590 ) | ( wire19306 ) | ( _34942 ) | ( _37639 ) ;
 assign o_15_ = ( wire590 ) | ( wire19306 ) | ( _37643 ) | ( _37648 ) ;
 assign o_32_ = ( wire590 ) | ( wire19306 ) | ( _34942 ) | ( _37657 ) ;
 assign o_23_ = ( n_n5231 ) | ( wire20753 ) | ( n_n4199 ) | ( _37703 ) ;
 assign o_18_ = ( n_n5235 ) | ( wire590 ) | ( wire19306 ) | ( _34942 ) ;
 assign o_31_ = ( wire590 ) | ( wire19306 ) | ( _34942 ) | ( _37967 ) ;
 assign o_24_ = ( wire20924 ) | ( wire590 ) | ( wire19306 ) | ( _34942 ) ;
 assign o_17_ = ( n_n5231 ) | ( n_n3089 ) | ( n_n3094 ) | ( wire21154 ) ;
 assign o_30_ = ( wire590 ) | ( wire19306 ) | ( _34942 ) | ( _38245 ) ;
 assign o_20_ = ( n_n5231 ) | ( n_n3892 ) | ( n_n3890 ) | ( wire21293 ) ;
 assign o_10_ = ( n_n5231 ) | ( _38468 ) | ( _38469 ) ;
 assign o_9_ = ( n_n5231 ) | ( n_n2058 ) | ( wire21620 ) | ( wire21621 ) ;
 assign o_7_ = ( wire590 ) | ( wire19306 ) | ( _34942 ) | ( _38932 ) ;
 assign o_8_ = ( wire21881 ) | ( _39346 ) | ( _39384 ) ;
 assign o_5_ = ( n_n5231 ) | ( wire22331 ) | ( wire22334 ) ;
 assign o_6_ = ( wire2474 ) | ( wire590 ) | ( wire19306 ) | ( _37643 ) ;
 assign o_3_ = ( _40392 ) | ( _40393 ) | ( _40395 ) | ( _40442 ) ;
 assign o_4_ = ( wire22827 ) | ( _40811 ) | ( _40859 ) ;
 assign n_n5231 = ( wire590 ) | ( wire19306 ) | ( _34942 ) ;
 assign wire19373 = ( n_n4476 ) | ( wire893 ) | ( wire19363 ) | ( wire19364 ) ;
 assign wire19374 = ( n_n4477 ) | ( wire507 ) | ( wire5797 ) | ( wire19369 ) ;
 assign n_n3621 = ( wire19489 ) | ( wire19490 ) | ( _35131 ) | ( _35341 ) ;
 assign wire19592 = ( n_n3625 ) | ( n_n3626 ) | ( n_n3624 ) | ( wire19422 ) ;
 assign wire19593 = ( n_n3627 ) | ( n_n3631 ) | ( n_n3632 ) | ( wire19588 ) ;
 assign wire19601 = ( wire535 ) | ( wire19599 ) | ( _5905 ) | ( _5910 ) ;
 assign wire19622 = ( wire19619 ) | ( wire19620 ) | ( _35815 ) ;
 assign wire19648 = ( n_n4442 ) | ( n_n4439 ) | ( wire19644 ) | ( wire19645 ) ;
 assign n_n5792 = ( i_5_  &  i_3_  &  n_n165  &  _35831 ) ;
 assign n_n5794 = ( i_5_  &  i_3_  &  n_n165  &  _35833 ) ;
 assign wire19766 = ( n_n4203 ) | ( wire19757 ) | ( _36234 ) | ( _36235 ) ;
 assign wire19822 = ( n_n2572 ) | ( wire19812 ) | ( _36312 ) ;
 assign wire19846 = ( n_n3550 ) | ( wire19842 ) | ( n_n207  &  wire1813 ) ;
 assign wire19847 = ( wire887 ) | ( wire19843 ) | ( n_n227  &  wire1814 ) ;
 assign n_n4718 = ( n_n4723 ) | ( n_n4725 ) | ( wire19980 ) | ( wire19981 ) ;
 assign wire19989 = ( wire19888 ) | ( _36487 ) | ( _36488 ) | ( _36508 ) ;
 assign wire19990 = ( n_n4736 ) | ( n_n3397 ) | ( _36558 ) ;
 assign n_n264 = ( i_5_  &  (~ i_3_)  &  (~ i_4_) ) ;
 assign n_n153 = ( i_7_  &  i_6_ ) ;
 assign n_n120 = ( i_1_  &  (~ i_2_)  &  i_0_ ) ;
 assign wire20002 = ( wire777 ) | ( n_n5675 ) | ( wire4928 ) | ( wire19999 ) ;
 assign wire20004 = ( wire879 ) | ( n_n2772 ) | ( wire19996 ) | ( wire19997 ) ;
 assign n_n5224 = ( n_n4416 ) | ( n_n4418 ) | ( wire20033 ) | ( wire20034 ) ;
 assign n_n2657 = ( wire20094 ) | ( wire20084 ) | ( wire20088 ) | ( _36797 ) ;
 assign wire20115 = ( n_n2659 ) | ( wire20054 ) | ( wire20055 ) | ( wire20113 ) ;
 assign wire20245 = ( n_n4533 ) | ( wire20166 ) | ( _37077 ) | ( _37108 ) ;
 assign wire20355 = ( n_n3900 ) | ( n_n3899 ) | ( n_n3901 ) | ( n_n4141 ) ;
 assign n_n2789 = ( n_n2793 ) | ( wire20571 ) | ( wire20484 ) | ( _37352 ) ;
 assign n_n2795 = ( wire20614 ) | ( wire4267 ) | ( _4018 ) | ( _37544 ) ;
 assign wire20625 = ( n_n2808 ) | ( n_n2806 ) | ( wire20590 ) | ( wire20624 ) ;
 assign n_n4508 = ( wire826 ) | ( wire4234 ) | ( wire4235 ) | ( wire4236 ) ;
 assign wire20648 = ( wire20636 ) | ( wire20646 ) | ( _37630 ) ;
 assign n_n4186 = ( wire372 ) | ( wire894 ) | ( wire20651 ) | ( wire20652 ) ;
 assign wire20658 = ( wire392 ) | ( wire20655 ) | ( n_n241  &  n_n104 ) ;
 assign wire879 = ( i_7_  &  i_6_  &  wire929 ) | ( (~ i_7_)  &  i_6_  &  wire929 ) | ( i_7_  &  (~ i_6_)  &  wire929 ) | ( (~ i_7_)  &  i_6_  &  wire936 ) | ( i_7_  &  (~ i_6_)  &  wire936 ) | ( (~ i_7_)  &  (~ i_6_)  &  wire936 ) ;
 assign wire20665 = ( _37645 ) | ( _37646 ) ;
 assign n_n5797 = ( i_5_  &  i_3_  &  n_n165  &  _35820 ) ;
 assign wire20667 = ( n_n153  &  n_n260  &  n_n165 ) | ( n_n153  &  n_n165  &  n_n284 ) ;
 assign wire20671 = ( n_n5796 ) | ( wire4202 ) | ( wire20668 ) ;
 assign wire20753 = ( wire20751 ) | ( _37733 ) ;
 assign n_n5235 = ( n_n3361 ) | ( n_n3360 ) | ( wire20913 ) | ( wire20914 ) ;
 assign wire3945 = ( _3570 ) | ( (~ i_9_)  &  (~ i_10_)  &  wire20917 ) ;
 assign wire20920 = ( n_n5693 ) | ( wire452 ) | ( wire5441 ) | ( wire5442 ) ;
 assign wire20924 = ( _3566 ) | ( _3567 ) | ( wire396  &  _37968 ) ;
 assign n_n3089 = ( n_n3092 ) | ( n_n3093 ) | ( wire21131 ) ;
 assign n_n3094 = ( n_n3107 ) | ( n_n3108 ) | ( wire21148 ) ;
 assign wire21154 = ( wire20931 ) | ( wire21153 ) | ( _38183 ) | ( _38202 ) ;
 assign wire21178 = ( n_n4476 ) | ( n_n4477 ) | ( wire3712 ) | ( wire21175 ) ;
 assign n_n3892 = ( n_n3900 ) | ( n_n3899 ) | ( wire20319 ) | ( _37231 ) ;
 assign n_n3890 = ( n_n3895 ) | ( n_n3904 ) | ( _38319 ) | ( _38320 ) ;
 assign wire21293 = ( n_n3898 ) | ( n_n3897 ) | ( n_n3913 ) | ( _38374 ) ;
 assign n_n2058 = ( n_n2067 ) | ( _38635 ) | ( _38636 ) | ( _38637 ) ;
 assign wire21620 = ( n_n2073 ) | ( wire21396 ) | ( _38670 ) | ( _38734 ) ;
 assign wire21621 = ( n_n2063 ) | ( n_n2064 ) | ( _38902 ) ;
 assign n_n1670 = ( _2448 ) | ( _2449 ) | ( wire1825  &  _38906 ) ;
 assign wire21904 = ( wire21885 ) | ( n_n1693 ) | ( wire21902 ) | ( _39356 ) ;
 assign wire22331 = ( n_n1089 ) | ( wire21927 ) | ( wire21928 ) | ( wire21950 ) ;
 assign wire22334 = ( wire22326 ) | ( wire22327 ) | ( wire22328 ) | ( wire22332 ) ;
 assign wire2474 = ( i_3_  &  (~ i_1_)  &  i_2_  &  (~ i_0_) ) | ( i_3_  &  (~ i_1_)  &  (~ i_2_)  &  (~ i_0_) ) ;
 assign wire22594 = ( wire22338 ) | ( wire22593 ) | ( _40404 ) | ( _40441 ) ;
 assign wire22847 = ( _40857 ) | ( _40858 ) ;
 assign n_n260 = ( (~ i_5_)  &  (~ i_3_)  &  i_4_ ) ;
 assign n_n229 = ( (~ i_7_)  &  (~ i_8_)  &  i_6_ ) ;
 assign n_n165 = ( i_1_  &  (~ i_2_)  &  (~ i_0_) ) ;
 assign n_n139 = ( n_n260  &  n_n229  &  n_n165 ) ;
 assign wire913 = ( (~ i_9_)  &  i_10_  &  (~ i_11_)  &  (~ i_15_) ) ;
 assign n_n151 = ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  wire913 ) ;
 assign n_n116 = ( (~ i_1_)  &  (~ i_2_)  &  i_0_ ) ;
 assign n_n5686 = ( (~ i_7_)  &  (~ i_6_)  &  n_n260  &  n_n116 ) ;
 assign wire590 = ( wire19341 ) | ( wire19323 ) | ( _34606 ) | ( _34685 ) ;
 assign wire19306 = ( n_n5007 ) | ( n_n5048 ) | ( wire19303 ) | ( wire19305 ) ;
 assign wire19359 = ( i_1_  &  i_2_ ) | ( i_2_  &  (~ i_0_) ) | ( i_3_  &  i_1_  &  (~ i_2_)  &  i_0_ ) | ( i_3_  &  (~ i_1_)  &  (~ i_2_)  &  (~ i_0_) ) ;
 assign wire19365 = ( wire826 ) | ( n_n281  &  wire914  &  wire1474 ) ;
 assign wire48 = ( i_15_  &  n_n281  &  n_n242 ) | ( (~ i_15_)  &  n_n242  &  n_n279 ) ;
 assign wire503 = ( i_7_  &  (~ i_6_)  &  n_n260  &  n_n165 ) ;
 assign n_n152 = ( n_n260  &  n_n165  &  n_n283 ) ;
 assign n_n4476 = ( wire503 ) | ( wire48  &  n_n152 ) ;
 assign n_n220 = ( (~ i_14_)  &  i_13_  &  (~ i_12_) ) ;
 assign wire54 = ( n_n247  &  _34949 ) | ( n_n247  &  _34950 ) ;
 assign n_n4477 = ( n_n152  &  wire54 ) | ( wire913  &  n_n152  &  n_n220 ) ;
 assign wire394 = ( i_7_  &  i_6_  &  n_n260  &  n_n165 ) ;
 assign wire927 = ( (~ i_1_)  &  (~ i_2_)  &  i_0_  &  _34990 ) ;
 assign wire929 = ( (~ i_1_)  &  (~ i_2_)  &  i_0_  &  _34985 ) ;
 assign wire507 = ( i_7_  &  i_6_  &  wire927 ) | ( (~ i_7_)  &  i_6_  &  wire927 ) | ( i_7_  &  (~ i_6_)  &  wire927 ) | ( (~ i_7_)  &  i_6_  &  wire929 ) | ( i_7_  &  (~ i_6_)  &  wire929 ) | ( (~ i_7_)  &  (~ i_6_)  &  wire929 ) ;
 assign n_n111 = ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  wire914 ) ;
 assign wire103 = ( n_n259  &  _34953 ) | ( n_n259  &  _34954 ) ;
 assign wire266 = ( (~ i_9_)  &  (~ i_10_) ) | ( n_n220  &  wire905 ) ;
 assign wire893 = ( n_n152  &  n_n111 ) | ( n_n152  &  wire103 ) | ( n_n152  &  wire266 ) ;
 assign n_n208 = ( (~ i_7_)  &  i_8_  &  i_6_ ) ;
 assign n_n273 = ( (~ i_7_)  &  i_8_  &  (~ i_6_) ) ;
 assign wire937 = ( n_n260  &  n_n165  &  n_n208 ) | ( n_n260  &  n_n165  &  n_n273 ) ;
 assign wire372 = ( n_n177  &  n_n200 ) | ( n_n189  &  n_n101 ) ;
 assign wire386 = ( n_n177  &  n_n45 ) | ( n_n189  &  n_n102 ) ;
 assign wire19380 = ( wire392 ) | ( wire19377 ) | ( n_n255  &  n_n31 ) ;
 assign n_n3424 = ( wire5720 ) | ( _35346 ) ;
 assign n_n3642 = ( n_n3778 ) | ( wire812 ) | ( _6319 ) | ( _35354 ) ;
 assign wire19431 = ( n_n3757 ) | ( wire5709 ) | ( _35359 ) ;
 assign wire19435 = ( n_n2598 ) | ( wire5699 ) | ( _6294 ) | ( _35372 ) ;
 assign n_n3625 = ( n_n3424 ) | ( n_n3642 ) | ( wire19431 ) | ( wire19435 ) ;
 assign n_n3382 = ( wire19440 ) | ( _6287 ) | ( _35379 ) | ( _35384 ) ;
 assign wire19445 = ( n_n3727 ) | ( wire409 ) | ( wire546 ) | ( wire19443 ) ;
 assign wire19446 = ( wire5681 ) | ( wire19442 ) | ( _35414 ) ;
 assign wire19455 = ( wire694 ) | ( wire544 ) | ( wire19452 ) | ( wire19453 ) ;
 assign n_n3626 = ( n_n3382 ) | ( wire19445 ) | ( wire19446 ) | ( wire19455 ) ;
 assign n_n3645 = ( wire19465 ) | ( wire19466 ) | ( wire19467 ) ;
 assign wire19472 = ( wire5651 ) | ( wire19470 ) ;
 assign wire19473 = ( n_n3806 ) | ( wire5650 ) | ( wire5656 ) | ( wire5657 ) ;
 assign wire19480 = ( n_n3686 ) | ( wire5643 ) | ( wire19475 ) | ( wire19478 ) ;
 assign n_n3627 = ( n_n3645 ) | ( wire19472 ) | ( wire19473 ) | ( wire19480 ) ;
 assign wire19530 = ( wire19528 ) | ( _35257 ) | ( _35258 ) | ( _35339 ) ;
 assign n_n4781 = ( wire5552 ) | ( wire5550 ) | ( n_n57  &  wire44 ) ;
 assign n_n3711 = ( _6077 ) | ( _35565 ) ;
 assign wire19544 = ( n_n3709 ) | ( n_n4680 ) | ( n_n4677 ) | ( wire19534 ) ;
 assign wire19546 = ( n_n3708 ) | ( wire19541 ) | ( _35588 ) ;
 assign n_n3631 = ( n_n4781 ) | ( n_n3711 ) | ( wire19544 ) | ( wire19546 ) ;
 assign wire19553 = ( wire471 ) | ( wire19549 ) | ( wire19550 ) ;
 assign wire19554 = ( n_n1641 ) | ( wire5516 ) | ( wire5517 ) ;
 assign n_n3661 = ( wire19553 ) | ( wire19554 ) | ( _5967 ) | ( _5968 ) ;
 assign n_n3632 = ( wire19565 ) | ( wire19566 ) | ( _35613 ) | ( _35640 ) ;
 assign n_n284 = ( (~ i_5_)  &  (~ i_3_)  &  (~ i_4_) ) ;
 assign n_n124 = ( n_n229  &  n_n165  &  n_n284 ) ;
 assign n_n123 = ( n_n165  &  n_n208  &  n_n284 ) ;
 assign wire289 = ( i_7_  &  i_6_ ) | ( (~ i_7_)  &  i_6_ ) | ( i_7_  &  (~ i_6_) ) ;
 assign wire364 = ( i_7_  &  i_6_  &  n_n165  &  n_n284 ) ;
 assign wire535 = ( i_7_  &  i_6_  &  n_n264  &  n_n116 ) | ( i_7_  &  (~ i_6_)  &  n_n264  &  n_n116 ) ;
 assign wire777 = ( (~ i_7_)  &  i_6_  &  n_n264  &  n_n116 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n264  &  n_n116 ) ;
 assign n_n118 = ( (~ i_1_)  &  i_2_  &  i_0_ ) ;
 assign wire834 = ( (~ i_7_)  &  (~ i_6_)  &  n_n264  &  n_n118 ) ;
 assign n_n281 = ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_) ) ;
 assign wire914 = ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  (~ i_15_) ) ;
 assign wire907 = ( (~ i_9_)  &  (~ i_10_)  &  (~ i_11_)  &  (~ i_15_) ) ;
 assign wire939 = ( wire913  &  n_n281 ) | ( n_n281  &  wire914 ) | ( n_n281  &  wire907 ) ;
 assign n_n110 = ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  wire913 ) ;
 assign n_n106 = ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  wire907 ) ;
 assign n_n5678 = ( (~ i_7_)  &  (~ i_6_)  &  n_n116  &  n_n284 ) ;
 assign n_n5671 = ( i_7_  &  i_6_  &  n_n264  &  n_n116 ) ;
 assign wire396 = ( n_n165  &  n_n208  &  n_n284 ) | ( n_n165  &  n_n273  &  n_n284 ) ;
 assign wire880 = ( i_7_  &  i_6_  &  n_n116  &  n_n284 ) | ( i_7_  &  (~ i_6_)  &  n_n116  &  n_n284 ) ;
 assign n_n5677 = ( (~ i_7_)  &  i_6_  &  n_n116  &  n_n284 ) ;
 assign n_n5672 = ( i_7_  &  (~ i_6_)  &  n_n264  &  n_n116 ) ;
 assign wire582 = ( wire777 ) | ( wire880 ) | ( n_n5677 ) | ( n_n5672 ) ;
 assign wire5453 = ( i_7_  &  i_6_  &  n_n264  &  n_n118 ) | ( (~ i_7_)  &  i_6_  &  n_n264  &  n_n118 ) | ( i_7_  &  (~ i_6_)  &  n_n264  &  n_n118 ) ;
 assign wire19613 = ( n_n264  &  n_n118  &  n_n155 ) | ( n_n284  &  n_n118  &  n_n155 ) ;
 assign wire19614 = ( i_7_  &  i_6_  &  n_n284  &  n_n118 ) | ( (~ i_7_)  &  i_6_  &  n_n284  &  n_n118 ) | ( i_7_  &  (~ i_6_)  &  n_n284  &  n_n118 ) ;
 assign wire583 = ( wire5453 ) | ( wire19613 ) | ( wire19614 ) ;
 assign wire941 = ( n_n165  &  n_n208  &  n_n284 ) | ( n_n165  &  n_n273  &  n_n284 ) ;
 assign wire940 = ( wire913  &  n_n281 ) | ( n_n281  &  wire914 ) ;
 assign n_n272 = ( i_7_  &  (~ i_6_) ) ;
 assign wire19624 = ( n_n5693 ) | ( n_n220  &  wire914  &  n_n130 ) ;
 assign wire19625 = ( n_n5797 ) | ( wire5441 ) | ( wire5442 ) ;
 assign wire19626 = ( wire5439 ) | ( wire54  &  n_n128 ) | ( n_n111  &  n_n128 ) ;
 assign n_n4442 = ( wire19624 ) | ( wire19625 ) | ( wire19626 ) ;
 assign n_n4439 = ( n_n5797 ) | ( _35837 ) | ( n_n139  &  wire54 ) ;
 assign wire943 = ( i_5_  &  (~ i_3_)  &  i_4_  &  n_n118 ) | ( (~ i_5_)  &  (~ i_3_)  &  i_4_  &  n_n118 ) | ( i_5_  &  (~ i_3_)  &  (~ i_4_)  &  n_n118 ) ;
 assign n_n231 = ( (~ i_7_)  &  i_6_ ) ;
 assign wire19290 = ( i_5_  &  i_3_ ) ;
 assign wire573 = ( n_n5  &  wire70 ) | ( n_n6  &  n_n12 ) ;
 assign wire5389 = ( n_n5  &  wire101 ) | ( n_n220  &  n_n5  &  wire901 ) ;
 assign wire19654 = ( wire5390 ) | ( wire5400 ) | ( n_n5  &  wire1874 ) ;
 assign wire19655 = ( n_n4815 ) | ( n_n4821 ) | ( n_n4814 ) | ( n_n4816 ) ;
 assign n_n4203 = ( wire573 ) | ( wire5389 ) | ( wire19654 ) | ( wire19655 ) ;
 assign n_n4846 = ( n_n5  &  wire49 ) | ( n_n6  &  n_n22 ) ;
 assign n_n4842 = ( n_n5  &  n_n76 ) | ( n_n6  &  wire82 ) ;
 assign wire19659 = ( _5501 ) | ( _5502 ) ;
 assign n_n4206 = ( _5501 ) | ( _5502 ) | ( _36198 ) ;
 assign n_n1506 = ( n_n5  &  n_n42 ) | ( n_n6  &  wire81 ) ;
 assign wire19677 = ( wire5357 ) | ( wire5371 ) | ( wire5372 ) | ( wire19665 ) ;
 assign n_n6 = ( n_n285  &  n_n230  &  n_n261 ) ;
 assign wire911 = ( (~ i_9_)  &  i_10_  &  (~ i_11_)  &  i_15_ ) ;
 assign n_n228 = ( i_14_  &  i_13_  &  i_12_ ) ;
 assign wire75 = ( i_15_  &  n_n220  &  n_n242 ) | ( (~ i_15_)  &  n_n242  &  n_n258 ) ;
 assign n_n4807 = ( n_n6  &  wire75 ) | ( n_n6  &  wire911  &  n_n228 ) ;
 assign n_n4808 = ( wire75  &  n_n5 ) | ( wire913  &  n_n281  &  n_n5 ) ;
 assign n_n4809 = ( n_n6  &  wire72 ) | ( n_n206  &  n_n5 ) ;
 assign wire541 = ( n_n6  &  wire118 ) | ( n_n60  &  n_n5 ) ;
 assign n_n4223 = ( n_n4808 ) | ( n_n4809 ) | ( wire541 ) ;
 assign wire585 = ( n_n5  &  wire132 ) | ( n_n6  &  n_n59 ) ;
 assign wire5347 = ( n_n6  &  wire50 ) | ( n_n281  &  n_n6  &  wire903 ) ;
 assign wire5348 = ( n_n5  &  wire63 ) | ( n_n228  &  n_n5  &  wire902 ) ;
 assign n_n4224 = ( wire585 ) | ( wire5347 ) | ( wire5348 ) ;
 assign n_n4307 = ( wire5328 ) | ( wire19696 ) | ( _35959 ) | ( _35962 ) ;
 assign wire19717 = ( _5751 ) | ( _5752 ) | ( _35996 ) ;
 assign wire19718 = ( wire19703 ) | ( wire19704 ) | ( wire19709 ) | ( wire19710 ) ;
 assign n_n285 = ( (~ i_1_)  &  (~ i_2_)  &  (~ i_0_) ) ;
 assign n_n1 = ( n_n260  &  n_n273  &  n_n285 ) ;
 assign n_n283 = ( (~ i_7_)  &  (~ i_8_)  &  (~ i_6_) ) ;
 assign n_n2 = ( n_n260  &  n_n285  &  n_n283 ) ;
 assign n_n60 = ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  wire908 ) ;
 assign wire118 = ( n_n259  &  _35950 ) | ( n_n259  &  _35951 ) ;
 assign n_n2618 = ( n_n2  &  n_n60 ) | ( n_n1  &  wire118 ) ;
 assign n_n206 = ( i_14_  &  i_13_  &  i_12_  &  wire911 ) ;
 assign wire72 = ( n_n259  &  _34638 ) | ( n_n259  &  _34639 ) ;
 assign n_n5769 = ( i_7_  &  (~ i_6_)  &  n_n165  &  n_n284 ) ;
 assign n_n127 = ( n_n165  &  n_n284  &  n_n283 ) ;
 assign wire19835 = ( wire5138 ) | ( _5346 ) | ( _5347 ) ;
 assign n_n242 = ( (~ i_9_)  &  i_10_  &  (~ i_11_) ) ;
 assign n_n279 = ( i_14_  &  (~ i_13_)  &  (~ i_12_) ) ;
 assign n_n266 = ( i_7_  &  i_8_  &  i_6_ ) ;
 assign n_n265 = ( n_n284  &  n_n285  &  n_n266 ) ;
 assign n_n271 = ( i_7_  &  (~ i_8_)  &  i_6_ ) ;
 assign n_n268 = ( n_n284  &  n_n285  &  n_n271 ) ;
 assign wire273 = ( (~ i_14_)  &  i_13_  &  i_12_  &  wire912 ) | ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire912 ) | ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  wire912 ) ;
 assign n_n2550 = ( _5302 ) | ( n_n268  &  wire273 ) ;
 assign wire5115 = ( n_n265  &  wire101 ) | ( n_n281  &  wire907  &  n_n265 ) ;
 assign wire5116 = ( n_n268  &  wire95 ) | ( n_n268  &  n_n11 ) | ( n_n268  &  wire19848 ) ;
 assign wire19849 = ( n_n268  &  n_n148 ) | ( n_n265  &  n_n62 ) ;
 assign n_n2545 = ( wire5115 ) | ( wire5116 ) | ( wire19849 ) ;
 assign wire268 = ( (~ i_14_)  &  i_13_  &  i_12_  &  wire907 ) | ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire907 ) | ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  wire907 ) ;
 assign wire200 = ( (~ i_14_)  &  i_13_  &  i_12_  &  wire901 ) | ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire901 ) | ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  wire901 ) ;
 assign wire112 = ( i_14_  &  i_13_  &  i_12_  &  wire907 ) | ( i_14_  &  i_13_  &  (~ i_12_)  &  wire907 ) | ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire907 ) ;
 assign n_n155 = ( (~ i_7_)  &  (~ i_6_) ) ;
 assign n_n5796 = ( (~ i_7_)  &  (~ i_6_)  &  n_n165  &  _36410 ) ;
 assign n_n5 = ( n_n285  &  n_n230  &  n_n263 ) ;
 assign n_n4723 = ( wire19936 ) | ( wire19946 ) | ( _36404 ) | ( _36417 ) ;
 assign n_n4725 = ( wire19959 ) | ( wire19967 ) | ( _36424 ) | ( _36450 ) ;
 assign wire19980 = ( n_n4954 ) | ( n_n4953 ) | ( wire672 ) | ( _36457 ) ;
 assign wire19981 = ( wire19926 ) | ( wire19927 ) | ( wire19973 ) | ( wire19974 ) ;
 assign wire4935 = ( i_7_  &  i_6_  &  n_n118  &  n_n230 ) ;
 assign n_n2772 = ( wire5453 ) | ( wire19613 ) | ( wire19614 ) | ( wire4935 ) ;
 assign n_n230 = ( i_5_  &  (~ i_3_)  &  i_4_ ) ;
 assign n_n130 = ( n_n229  &  n_n165  &  n_n230 ) ;
 assign n_n121 = ( n_n264  &  n_n165  &  n_n271 ) ;
 assign n_n132 = ( n_n165  &  n_n283  &  n_n230 ) ;
 assign wire1686 = ( wire913  &  n_n220 ) | ( n_n220  &  wire914 ) | ( n_n220  &  wire905 ) ;
 assign wire20007 = ( n_n111  &  n_n127 ) | ( n_n127  &  n_n108 ) | ( n_n108  &  n_n122 ) ;
 assign wire1705 = ( wire913  &  n_n220 ) | ( n_n220  &  wire914 ) ;
 assign wire20008 = ( n_n110  &  n_n127 ) | ( n_n139  &  wire1703 ) ;
 assign wire949 = ( wire913  &  n_n220 ) | ( n_n220  &  wire914 ) ;
 assign wire905 = ( i_9_  &  i_10_  &  (~ i_11_)  &  (~ i_15_) ) ;
 assign wire948 = ( wire913  &  n_n220 ) | ( n_n220  &  wire905 ) ;
 assign n_n4416 = ( wire4889 ) | ( wire20020 ) | ( wire20021 ) ;
 assign n_n4418 = ( wire4882 ) | ( wire20023 ) | ( wire20027 ) ;
 assign wire20033 = ( wire4902 ) | ( wire20015 ) | ( wire20030 ) | ( wire20031 ) ;
 assign wire20034 = ( wire4896 ) | ( wire4899 ) | ( wire20016 ) | ( wire20017 ) ;
 assign n_n4549 = ( n_n4256 ) | ( wire5011 ) | ( wire20122 ) | ( _36959 ) ;
 assign n_n4544 = ( wire20141 ) | ( wire20142 ) | ( _4675 ) | ( _37004 ) ;
 assign wire20147 = ( wire4745 ) | ( wire20131 ) | ( _37030 ) ;
 assign n_n4533 = ( n_n4544 ) | ( wire20147 ) | ( wire20134 ) | ( _37002 ) ;
 assign wire20166 = ( n_n1490 ) | ( n_n4628 ) | ( _37076 ) ;
 assign wire20184 = ( n_n4806 ) | ( wire4690 ) | ( _4559 ) | ( _37104 ) ;
 assign n_n4556 = ( n_n4681 ) | ( _4777 ) | ( _4778 ) | ( _36894 ) ;
 assign n_n4535 = ( n_n3709 ) | ( n_n4551 ) | ( wire20228 ) | ( wire20232 ) ;
 assign wire20240 = ( wire20216 ) | ( wire20238 ) | ( _36947 ) ;
 assign n_n3900 = ( n_n3925 ) | ( wire20262 ) | ( wire20271 ) | ( _37140 ) ;
 assign n_n3899 = ( n_n3920 ) | ( n_n3922 ) | ( wire4552 ) | ( wire20293 ) ;
 assign n_n3901 = ( _4365 ) | ( _4366 ) | ( _37230 ) | ( _37231 ) ;
 assign n_n3918 = ( n_n3974 ) | ( wire20330 ) | ( wire20331 ) ;
 assign n_n3919 = ( n_n4153 ) | ( n_n4154 ) | ( wire20340 ) | ( wire20341 ) ;
 assign wire20353 = ( wire298 ) | ( n_n4146 ) | ( wire20349 ) | ( wire20350 ) ;
 assign n_n4141 = ( n_n3918 ) | ( n_n3919 ) | ( wire20353 ) ;
 assign n_n4 = ( n_n208  &  n_n284  &  n_n285 ) ;
 assign wire912 = ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  i_15_ ) ;
 assign wire95 = ( n_n247  &  _36179 ) | ( n_n247  &  _36180 ) ;
 assign n_n4015 = ( n_n4  &  wire95 ) | ( n_n228  &  n_n4  &  wire912 ) ;
 assign n_n2793 = ( n_n2804 ) | ( wire20553 ) | ( _37378 ) | ( _37379 ) ;
 assign wire20571 = ( n_n2815 ) | ( n_n2817 ) | ( wire20412 ) | ( _37523 ) ;
 assign wire20614 = ( wire4276 ) | ( wire4281 ) | ( wire20600 ) | ( wire20606 ) ;
 assign n_n3727 = ( n_n60  &  n_n4 ) | ( n_n4  &  n_n8 ) | ( n_n4  &  n_n61 ) ;
 assign n_n9 = ( i_14_  &  i_13_  &  i_12_  &  wire902 ) ;
 assign wire4264 = ( n_n4  &  wire113 ) | ( n_n4  &  wire50 ) | ( n_n4  &  n_n59 ) ;
 assign n_n2840 = ( n_n3727 ) | ( wire4264 ) | ( n_n4  &  n_n9 ) ;
 assign wire4259 = ( n_n151  &  n_n4 ) | ( wire75  &  n_n4 ) | ( n_n206  &  n_n4 ) ;
 assign wire20616 = ( n_n4  &  _37580 ) | ( n_n4  &  wire899  &  _37091 ) ;
 assign wire20617 = ( n_n4  &  n_n145 ) | ( n_n4  &  n_n7 ) | ( n_n4  &  n_n144 ) ;
 assign n_n2839 = ( wire4259 ) | ( wire20616 ) | ( wire20617 ) ;
 assign n_n128 = ( n_n165  &  n_n271  &  n_n230 ) ;
 assign n_n5682 = ( (~ i_7_)  &  (~ i_6_)  &  n_n116  &  n_n230 ) ;
 assign n_n5676 = ( i_7_  &  (~ i_6_)  &  n_n116  &  n_n284 ) ;
 assign wire20629 = ( n_n121  &  wire216 ) | ( n_n132  &  n_n107 ) ;
 assign wire20630 = ( n_n122  &  wire1707 ) | ( n_n130  &  wire1706 ) ;
 assign wire826 = ( n_n260  &  n_n229  &  n_n165  &  n_n163 ) ;
 assign wire4234 = ( n_n132  &  wire216 ) | ( wire216  &  wire20637 ) | ( wire216  &  wire20638 ) ;
 assign wire4235 = ( n_n281  &  wire899  &  wire20637 ) | ( n_n281  &  wire899  &  wire20638 ) ;
 assign wire4236 = ( n_n260  &  n_n165  &  n_n283  &  n_n163 ) ;
 assign wire216 = ( n_n281  &  wire911 ) | ( n_n281  &  wire912 ) ;
 assign n_n255 = ( n_n260  &  n_n285  &  n_n271 ) ;
 assign wire894 = ( wire914  &  n_n279  &  n_n189 ) ;
 assign wire20651 = ( n_n177  &  n_n112 ) | ( n_n189  &  n_n109 ) ;
 assign wire20652 = ( n_n189  &  n_n102 ) | ( n_n177  &  n_n35 ) ;
 assign n_n241 = ( n_n260  &  n_n285  &  n_n266 ) ;
 assign n_n54 = ( i_14_  &  (~ i_13_)  &  i_12_  &  wire898 ) ;
 assign n_n105 = ( i_14_  &  (~ i_13_)  &  i_12_  &  wire900 ) ;
 assign wire392 = ( n_n255  &  n_n54 ) | ( n_n241  &  n_n105 ) ;
 assign n_n177 = ( n_n273  &  n_n285  &  n_n230 ) ;
 assign n_n216 = ( i_14_  &  (~ i_13_)  &  i_12_  &  wire911 ) ;
 assign n_n45 = ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire906 ) ;
 assign wire559 = ( n_n241  &  n_n216 ) | ( n_n177  &  n_n45 ) ;
 assign wire902 = ( i_9_  &  (~ i_10_)  &  i_11_  &  i_15_ ) ;
 assign n_n258 = ( i_14_  &  (~ i_13_)  &  i_12_ ) ;
 assign wire950 = ( wire912  &  n_n258 ) | ( wire902  &  n_n258 ) ;
 assign wire20662 = ( i_1_  &  i_2_  &  i_0_ ) | ( i_3_  &  i_1_  &  (~ i_2_)  &  i_0_ ) ;
 assign wire926 = ( i_2_  &  (~ i_0_) ) ;
 assign wire19753 = ( n_n4858 ) | ( n_n4864 ) | ( _5485 ) ;
 assign wire19754 = ( wire5244 ) | ( wire5228 ) | ( _36231 ) ;
 assign wire19758 = ( wire5238 ) | ( wire5242 ) | ( _36219 ) | ( _36222 ) ;
 assign n_n4219 = ( wire20705 ) | ( wire20706 ) | ( wire20710 ) ;
 assign n_n4199 = ( n_n4214 ) | ( n_n4255 ) | ( wire20729 ) | ( wire20733 ) ;
 assign wire20718 = ( n_n4279 ) | ( wire20703 ) | ( wire20704 ) | ( wire20716 ) ;
 assign n_n3361 = ( n_n3372 ) | ( n_n3371 ) | ( n_n3397 ) | ( _37777 ) ;
 assign n_n3360 = ( n_n3393 ) | ( wire20856 ) | ( _37846 ) | ( _37848 ) ;
 assign wire20913 = ( n_n3380 ) | ( n_n3379 ) | ( wire20872 ) | ( _37898 ) ;
 assign wire20914 = ( n_n3362 ) | ( wire20817 ) | ( wire20912 ) | ( _37934 ) ;
 assign n_n163 = ( (~ i_9_)  &  (~ i_10_) ) ;
 assign wire19294 = ( (~ i_5_)  &  i_3_  &  i_4_ ) ;
 assign n_n5693 = ( n_n165  &  n_n273  &  n_n163  &  wire19294 ) ;
 assign n_n274 = ( (~ i_9_)  &  i_10_ ) ;
 assign wire452 = ( n_n165  &  n_n283  &  wire19294  &  n_n274 ) ;
 assign wire19296 = ( (~ i_5_)  &  i_3_  &  (~ i_4_) ) ;
 assign wire758 = ( n_n165  &  n_n283  &  n_n274  &  wire19296 ) ;
 assign wire923 = ( i_9_  &  (~ i_10_) ) ;
 assign wire20925 = ( n_n3  &  n_n66 ) | ( n_n4  &  n_n148 ) ;
 assign wire20926 = ( n_n3  &  wire160 ) | ( n_n3  &  n_n252 ) | ( n_n3  &  n_n14 ) ;
 assign n_n3140 = ( n_n4015 ) | ( wire20925 ) | ( wire20926 ) ;
 assign n_n7424 = ( n_n228  &  n_n4  &  wire902 ) ;
 assign n_n3 = ( n_n229  &  n_n284  &  n_n285 ) ;
 assign n_n8 = ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  wire902 ) ;
 assign n_n61 = ( i_14_  &  (~ i_13_)  &  i_12_  &  wire908 ) ;
 assign n_n4005 = ( wire72  &  n_n3 ) | ( wire905  &  n_n258  &  n_n3 ) ;
 assign wire446 = ( n_n4  &  _37497 ) | ( n_n4  &  wire899  &  _35953 ) ;
 assign wire20946 = ( n_n4  &  _38195 ) | ( n_n4  &  wire899  &  _37091 ) ;
 assign wire20947 = ( n_n3  &  _38196 ) | ( n_n3  &  wire899  &  _37091 ) ;
 assign n_n3138 = ( n_n4005 ) | ( wire446 ) | ( wire20946 ) | ( wire20947 ) ;
 assign n_n3092 = ( n_n3099 ) | ( n_n3101 ) | ( wire21063 ) ;
 assign n_n3093 = ( n_n3103 ) | ( wire21122 ) | ( wire21116 ) | ( _38082 ) ;
 assign wire21131 = ( n_n3113 ) | ( n_n3097 ) | ( wire21129 ) | ( _38109 ) ;
 assign n_n3107 = ( wire3758 ) | ( wire21136 ) | ( _3973 ) | ( _37570 ) ;
 assign n_n3108 = ( wire3754 ) | ( _3324 ) | ( _38164 ) | ( _38165 ) ;
 assign wire21148 = ( wire21146 ) | ( _3319 ) | ( _3320 ) | ( _38174 ) ;
 assign n_n133 = ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  wire911 ) ;
 assign wire21186 = ( wire4302 ) | ( wire21183 ) | ( _3132 ) | ( _38325 ) ;
 assign n_n3898 = ( n_n3918 ) | ( n_n3919 ) | ( wire21186 ) ;
 assign n_n3895 = ( n_n3908 ) | ( wire3660 ) | ( wire3661 ) | ( wire21236 ) ;
 assign wire21220 = ( wire716 ) | ( wire3674 ) | ( wire3682 ) | ( wire21208 ) ;
 assign n_n3914 = ( n_n3964 ) | ( wire21250 ) | ( _3124 ) | ( _38330 ) ;
 assign n_n3915 = ( wire736 ) | ( wire21257 ) | ( wire21258 ) ;
 assign n_n3897 = ( n_n3914 ) | ( n_n3915 ) | ( wire21263 ) | ( _38343 ) ;
 assign n_n3913 = ( _3101 ) | ( _3102 ) | ( _38354 ) ;
 assign wire3626 = ( _3094 ) | ( _3095 ) | ( _3096 ) ;
 assign wire21276 = ( wire3627 ) | ( wire3629 ) | ( wire21268 ) | ( wire21269 ) ;
 assign n_n57 = ( n_n285  &  n_n266  &  n_n230 ) ;
 assign n_n56 = ( n_n285  &  n_n271  &  n_n230 ) ;
 assign n_n226 = ( i_14_  &  i_13_  &  i_12_  &  wire899 ) ;
 assign wire4059 = ( n_n151  &  n_n56 ) | ( wire75  &  n_n56 ) | ( n_n206  &  n_n56 ) ;
 assign wire4060 = ( n_n57  &  wire225 ) | ( n_n57  &  wire130 ) ;
 assign n_n2440 = ( wire4059 ) | ( wire4060 ) | ( n_n56  &  n_n226 ) ;
 assign n_n257 = ( i_14_  &  (~ i_13_)  &  i_12_  &  wire905 ) ;
 assign wire208 = ( n_n270  &  _35527 ) | ( n_n270  &  _35528 ) ;
 assign wire199 = ( n_n270  &  _35523 ) | ( n_n270  &  _35524 ) ;
 assign wire955 = ( wire72 ) | ( n_n257 ) | ( wire208 ) | ( wire199 ) ;
 assign n_n2073 = ( n_n2110 ) | ( wire21387 ) | ( _2760 ) | ( _2761 ) ;
 assign n_n2108 = ( wire3518 ) | ( wire21390 ) | ( n_n3  &  n_n186 ) ;
 assign wire21396 = ( n_n2104 ) | ( wire21394 ) | ( _38668 ) ;
 assign n_n145 = ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  wire905 ) ;
 assign wire21440 = ( n_n2126 ) | ( wire3470 ) | ( wire21435 ) | ( wire21438 ) ;
 assign n_n2067 = ( n_n2093 ) | ( wire21462 ) | ( wire21463 ) | ( wire21470 ) ;
 assign wire21508 = ( n_n2158 ) | ( wire21493 ) | ( wire21494 ) | ( wire21499 ) ;
 assign n_n2081 = ( wire3358 ) | ( wire21533 ) | ( _2611 ) | ( _38785 ) ;
 assign n_n2080 = ( n_n2133 ) | ( n_n2132 ) | ( wire21549 ) ;
 assign n_n2063 = ( n_n2081 ) | ( n_n2080 ) | ( n_n2137 ) | ( _38809 ) ;
 assign n_n2085 = ( n_n2148 ) | ( n_n2146 ) | ( wire21572 ) ;
 assign n_n2083 = ( n_n2140 ) | ( _2517 ) | ( _38846 ) | ( _38848 ) ;
 assign n_n2064 = ( n_n2085 ) | ( n_n2083 ) | ( n_n2145 ) | ( _38858 ) ;
 assign wire21612 = ( n_n2154 ) | ( _2458 ) | ( _2459 ) | ( _38898 ) ;
 assign wire169 = ( i_8_  &  n_n284  &  n_n231  &  n_n285 ) | ( (~ i_8_)  &  n_n284  &  n_n231  &  n_n285 ) ;
 assign n_n126 = ( n_n165  &  n_n273  &  n_n284 ) ;
 assign n_n5660 = ( (~ i_7_)  &  (~ i_6_)  &  n_n284  &  n_n118 ) ;
 assign n_n5659 = ( (~ i_7_)  &  i_6_  &  n_n284  &  n_n118 ) ;
 assign wire581 = ( (~ i_7_)  &  i_6_  &  n_n116  &  n_n284 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n116  &  n_n284 ) ;
 assign wire21635 = ( n_n4  &  n_n76 ) | ( n_n4  &  n_n25 ) | ( n_n4  &  n_n27 ) ;
 assign n_n1689 = ( n_n1713 ) | ( n_n1711 ) | ( wire21855 ) ;
 assign n_n1692 = ( wire21864 ) | ( wire21865 ) | ( wire21874 ) | ( wire21877 ) ;
 assign wire21881 = ( n_n1690 ) | ( n_n1691 ) | ( n_n1688 ) | ( n_n1687 ) ;
 assign wire21885 = ( wire2917 ) | ( wire2918 ) | ( wire21884 ) ;
 assign n_n1724 = ( wire21888 ) | ( wire21889 ) | ( _39363 ) ;
 assign wire21896 = ( n_n4  &  n_n144 ) | ( n_n4  &  n_n150 ) | ( n_n3  &  n_n150 ) ;
 assign n_n1693 = ( n_n1724 ) | ( _1861 ) | ( _39370 ) | ( _39372 ) ;
 assign n_n37 = ( i_14_  &  i_13_  &  (~ i_12_)  &  wire901 ) ;
 assign n_n83 = ( i_14_  &  i_13_  &  (~ i_12_)  &  wire907 ) ;
 assign wire154 = ( n_n282  &  _39005 ) | ( n_n282  &  _39006 ) ;
 assign wire64 = ( (~ i_14_)  &  i_13_  &  i_12_  &  wire901 ) | ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire901 ) ;
 assign n_n1111 = ( wire22007 ) | ( _1832 ) | ( _39387 ) | ( _39389 ) ;
 assign wire2808 = ( _1815 ) | ( _1816 ) ;
 assign wire21999 = ( wire823 ) | ( _1807 ) | ( n_n265  &  wire437 ) ;
 assign wire22014 = ( n_n1173 ) | ( wire22012 ) | ( _1796 ) | ( _1797 ) ;
 assign n_n1089 = ( n_n1111 ) | ( wire2808 ) | ( wire21999 ) | ( wire22014 ) ;
 assign n_n240 = ( i_14_  &  (~ i_13_)  &  i_12_  &  wire913 ) ;
 assign n_n246 = ( i_14_  &  (~ i_13_)  &  i_12_  &  wire914 ) ;
 assign wire1345 = ( i_8_  &  n_n284  &  n_n231  &  n_n285 ) | ( (~ i_8_)  &  n_n284  &  n_n231  &  n_n285 ) ;
 assign wire22360 = ( n_n4  &  n_n258  &  wire906 ) | ( n_n4  &  n_n258  &  wire908 ) ;
 assign wire22361 = ( n_n3  &  n_n252 ) | ( n_n4  &  wire1344 ) | ( n_n3  &  wire1344 ) ;
 assign n_n380 = ( wire22360 ) | ( wire22361 ) | ( n_n246  &  wire1345 ) ;
 assign wire1347 = ( n_n109 ) | ( wire143 ) | ( wire306 ) | ( wire22363 ) ;
 assign wire1346 = ( wire913  &  n_n256 ) | ( n_n258  &  wire904 ) ;
 assign n_n381 = ( n_n3  &  wire1347 ) | ( n_n4  &  wire1346 ) ;
 assign wire2163 = ( _92 ) | ( n_n3  &  wire22598 ) ;
 assign wire2169 = ( n_n4  &  wire19457 ) | ( n_n4  &  n_n25 ) | ( n_n4  &  wire22597 ) ;
 assign wire22602 = ( n_n876 ) | ( wire2162 ) | ( wire22600 ) ;
 assign n_n741 = ( n_n834 ) | ( wire2011 ) | ( wire22714 ) | ( wire22717 ) ;
 assign n_n740 = ( n_n762 ) | ( wire22744 ) | ( _40517 ) | ( _40518 ) ;
 assign wire22827 = ( n_n744 ) | ( wire22693 ) | ( _40807 ) | ( _40808 ) ;
 assign n_n775 = ( wire22829 ) | ( wire22830 ) | ( _40836 ) ;
 assign wire1837 = ( n_n203 ) | ( wire20149 ) | ( wire161 ) | ( wire22835 ) ;
 assign wire22839 = ( wire505 ) | ( wire22837 ) | ( n_n3  &  wire1836 ) ;
 assign n_n282 = ( (~ i_9_)  &  (~ i_10_)  &  (~ i_11_) ) ;
 assign n_n225 = ( (~ i_14_)  &  i_13_  &  i_12_ ) ;
 assign wire126 = ( i_15_  &  n_n282  &  n_n225 ) | ( (~ i_15_)  &  n_n282  &  n_n225 ) ;
 assign n_n189 = ( n_n285  &  n_n283  &  n_n230 ) ;
 assign wire6004 = ( i_9_  &  i_10_  &  i_12_  &  i_11_ ) | ( i_9_  &  (~ i_10_)  &  i_12_  &  i_11_ ) ;
 assign wire19279 = ( n_n279  &  wire902 ) | ( n_n253  &  n_n278 ) ;
 assign wire19280 = ( n_n279  &  wire912 ) | ( wire197  &  wire962 ) ;
 assign n_n5053 = ( n_n189  &  wire6004 ) | ( n_n189  &  wire19279 ) | ( n_n189  &  wire19280 ) ;
 assign wire5936 = ( (~ i_12_)  &  _34738 ) | ( i_13_  &  i_12_  &  _34738 ) | ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  _34738 ) ;
 assign wire19191 = ( wire913  &  n_n258 ) | ( n_n258  &  wire903 ) ;
 assign wire19192 = ( n_n267  &  wire965 ) | ( n_n267  &  _34730 ) ;
 assign n_n5061 = ( n_n241  &  wire5936 ) | ( n_n241  &  wire19191 ) | ( n_n241  &  wire19192 ) ;
 assign wire5931 = ( (~ i_12_)  &  _34748 ) | ( i_13_  &  i_12_  &  _34748 ) | ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  _34748 ) ;
 assign wire19194 = ( (~ i_9_) ) | ( wire914  &  n_n258 ) ;
 assign wire19195 = ( n_n258  &  wire908 ) | ( n_n247  &  wire968 ) ;
 assign n_n5062 = ( n_n255  &  wire5931 ) | ( n_n255  &  wire19194 ) | ( n_n255  &  wire19195 ) ;
 assign wire5922 = ( n_n241  &  wire19197 ) | ( n_n241  &  wire19198 ) ;
 assign wire5923 = ( (~ i_7_)  &  i_6_  &  n_n260  &  n_n285 ) ;
 assign n_n5020 = ( n_n5061 ) | ( n_n5062 ) | ( wire5922 ) | ( wire5923 ) ;
 assign wire898 = ( i_9_  &  i_10_  &  i_11_  &  i_15_ ) ;
 assign n_n99 = ( i_14_  &  i_13_  &  (~ i_12_)  &  wire898 ) ;
 assign n_n186 = ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire898 ) ;
 assign n_n222 = ( i_14_  &  i_13_  &  (~ i_12_) ) ;
 assign wire863 = ( n_n258  &  n_n57  &  wire898 ) | ( n_n57  &  wire898  &  n_n222 ) ;
 assign n_n4970 = ( n_n54  &  n_n57 ) | ( n_n57  &  n_n99 ) | ( n_n57  &  n_n186 ) ;
 assign wire906 = ( (~ i_9_)  &  i_10_  &  i_11_  &  (~ i_15_) ) ;
 assign wire153 = ( (~ i_14_)  &  i_13_  &  i_12_  &  wire906 ) | ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire906 ) | ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  wire906 ) ;
 assign wire901 = ( (~ i_9_)  &  (~ i_10_)  &  (~ i_11_)  &  i_15_ ) ;
 assign wire908 = ( i_9_  &  (~ i_10_)  &  i_11_  &  (~ i_15_) ) ;
 assign wire88 = ( n_n270  &  _35064 ) | ( n_n270  &  _35065 ) ;
 assign n_n4926 = ( n_n56  &  wire88 ) | ( n_n56  &  n_n222  &  wire908 ) ;
 assign wire5343 = ( n_n56  &  wire70 ) | ( n_n56  &  n_n14 ) | ( n_n56  &  wire256 ) ;
 assign wire5344 = ( n_n57  &  wire73 ) | ( n_n57  &  n_n65 ) | ( n_n57  &  n_n12 ) ;
 assign n_n261 = ( i_7_  &  i_8_  &  (~ i_6_) ) ;
 assign n_n263 = ( i_7_  &  (~ i_8_)  &  (~ i_6_) ) ;
 assign n_n108 = ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  wire905 ) ;
 assign wire70 = ( n_n253  &  _35084 ) | ( n_n253  &  _35085 ) ;
 assign n_n4826 = ( n_n5  &  n_n108 ) | ( n_n6  &  wire70 ) ;
 assign wire899 = ( i_9_  &  i_10_  &  (~ i_11_)  &  i_15_ ) ;
 assign n_n256 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_ ) ;
 assign wire66 = ( n_n259  &  _36143 ) | ( n_n259  &  _36144 ) ;
 assign n_n4828 = ( n_n5  &  wire66 ) | ( n_n5  &  wire899  &  n_n256 ) ;
 assign wire900 = ( (~ i_9_)  &  i_10_  &  i_11_  &  i_15_ ) ;
 assign wire73 = ( n_n267  &  _35086 ) | ( n_n267  &  _35087 ) ;
 assign n_n4823 = ( n_n6  &  wire73 ) | ( n_n6  &  n_n228  &  wire900 ) ;
 assign wire19738 = ( i_15_  &  n_n281  &  n_n242 ) | ( (~ i_15_)  &  n_n242  &  n_n225 ) ;
 assign wire44 = ( n_n253  &  _35042 ) | ( n_n253  &  _35043 ) ;
 assign n_n65 = ( i_14_  &  i_13_  &  i_12_  &  wire900 ) ;
 assign wire584 = ( n_n6  &  wire44 ) | ( n_n5  &  n_n65 ) ;
 assign n_n12 = ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  wire906 ) ;
 assign n_n70 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire905 ) ;
 assign wire79 = ( n_n259  &  _36138 ) | ( n_n259  &  _36139 ) ;
 assign wire5268 = ( n_n5  &  wire82 ) | ( n_n5  &  wire42 ) | ( n_n5  &  n_n223 ) ;
 assign wire5269 = ( wire913  &  n_n220  &  n_n6 ) ;
 assign wire19742 = ( n_n4826 ) | ( n_n4828 ) | ( n_n4823 ) | ( wire584 ) ;
 assign wire63 = ( n_n270  &  _35034 ) | ( n_n270  &  _35035 ) ;
 assign n_n4815 = ( n_n6  &  wire63 ) | ( n_n6  &  n_n228  &  wire902 ) ;
 assign n_n11 = ( i_14_  &  i_13_  &  i_12_  &  wire912 ) ;
 assign n_n4821 = ( n_n5  &  wire44 ) | ( n_n6  &  n_n11 ) ;
 assign wire137 = ( n_n275  &  _35053 ) | ( n_n275  &  _35054 ) ;
 assign n_n4814 = ( n_n6  &  n_n60 ) | ( n_n5  &  wire137 ) ;
 assign n_n4816 = ( n_n5  &  wire95 ) | ( n_n281  &  wire914  &  n_n5 ) ;
 assign wire60 = ( i_15_  &  n_n242  &  n_n258 ) | ( i_15_  &  n_n242  &  n_n222 ) ;
 assign n_n4834 = ( n_n110  &  n_n5 ) | ( n_n6  &  wire60 ) ;
 assign wire166 = ( i_14_  &  i_13_  &  i_12_  &  wire906 ) | ( i_14_  &  i_13_  &  (~ i_12_)  &  wire906 ) | ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire906 ) ;
 assign n_n4961 = ( n_n285  &  n_n266  &  n_n230  &  wire166 ) ;
 assign wire224 = ( i_14_  &  (~ i_13_)  &  i_12_  &  wire900 ) | ( i_14_  &  i_13_  &  (~ i_12_)  &  wire900 ) | ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire900 ) ;
 assign n_n95 = ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  wire904 ) ;
 assign n_n49 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire904 ) ;
 assign n_n96 = ( (~ i_14_)  &  i_13_  &  i_12_  &  wire904 ) ;
 assign n_n4967 = ( n_n57  &  n_n95 ) | ( n_n57  &  n_n49 ) | ( n_n57  &  n_n96 ) ;
 assign wire613 = ( n_n56  &  wire153 ) | ( n_n57  &  wire224 ) ;
 assign wire99 = ( (~ i_14_)  &  i_13_  &  i_12_  &  wire898 ) | ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire898 ) | ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  wire898 ) ;
 assign wire41 = ( i_14_  &  i_13_  &  i_12_  &  wire904 ) | ( i_14_  &  i_13_  &  (~ i_12_)  &  wire904 ) | ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire904 ) ;
 assign wire614 = ( n_n57  &  wire99 ) | ( n_n57  &  wire41 ) ;
 assign wire5033 = ( n_n151  &  n_n57 ) | ( wire75  &  n_n57 ) | ( n_n206  &  n_n57 ) ;
 assign n_n4287 = ( n_n5796 ) | ( wire72  &  n_n56 ) ;
 assign wire904 = ( i_9_  &  i_10_  &  i_11_  &  (~ i_15_) ) ;
 assign wire389 = ( n_n220  &  n_n6  &  wire904 ) | ( n_n6  &  n_n256  &  wire904 ) ;
 assign wire708 = ( n_n5  &  wire224 ) | ( n_n6  &  n_n96 ) ;
 assign wire4196 = ( n_n285  &  n_n230  &  n_n261  &  wire99 ) ;
 assign wire20675 = ( n_n4287 ) | ( wire389 ) | ( wire632 ) | ( wire5613 ) ;
 assign n_n4211 = ( wire20675 ) | ( _37722 ) ;
 assign wire180 = ( (~ i_14_)  &  i_13_  &  i_12_  &  wire900 ) | ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire900 ) | ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  wire900 ) ;
 assign wire617 = ( n_n6  &  wire166 ) | ( n_n6  &  wire180 ) ;
 assign wire254 = ( i_14_  &  (~ i_13_)  &  i_12_  &  wire898 ) | ( i_14_  &  i_13_  &  (~ i_12_)  &  wire898 ) | ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire898 ) ;
 assign wire673 = ( n_n5  &  wire41 ) | ( n_n5  &  wire254 ) ;
 assign wire674 = ( n_n5  &  wire153 ) | ( n_n5  &  wire180 ) ;
 assign wire20677 = ( n_n6  &  wire153 ) | ( n_n6  &  wire224 ) ;
 assign wire20678 = ( n_n6  &  wire166 ) | ( n_n5  &  wire166 ) | ( n_n6  &  wire180 ) ;
 assign n_n4210 = ( wire673 ) | ( wire674 ) | ( wire20677 ) | ( wire20678 ) ;
 assign n_n4892 = ( n_n56  &  wire63 ) | ( n_n228  &  wire902  &  n_n56 ) ;
 assign wire113 = ( n_n282  &  _35883 ) | ( n_n282  &  _35884 ) ;
 assign n_n4898 = ( n_n56  &  n_n11 ) | ( n_n57  &  wire113 ) ;
 assign n_n4895 = ( n_n60  &  n_n57 ) | ( n_n56  &  wire137 ) ;
 assign wire132 = ( n_n275  &  _35051 ) | ( n_n275  &  _35052 ) ;
 assign wire5035 = ( n_n57  &  n_n7 ) | ( n_n57  &  wire50 ) | ( n_n57  &  n_n59 ) ;
 assign wire5031 = ( wire118  &  n_n57 ) | ( wire72  &  n_n57 ) ;
 assign wire878 = ( _36510 ) | ( wire118  &  n_n57 ) | ( wire72  &  n_n57 ) ;
 assign n_n48 = ( n_n264  &  n_n285  &  n_n283 ) ;
 assign wire51 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire906 ) | ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  wire906 ) ;
 assign n_n53 = ( n_n264  &  n_n273  &  n_n285 ) ;
 assign n_n4179 = ( n_n48  &  wire51 ) | ( n_n105  &  n_n53 ) ;
 assign wire903 = ( (~ i_9_)  &  (~ i_10_)  &  i_11_  &  (~ i_15_) ) ;
 assign wire40 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire903 ) | ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  wire903 ) ;
 assign n_n31 = ( i_14_  &  (~ i_13_)  &  i_12_  &  wire902 ) ;
 assign n_n4168 = ( n_n53  &  wire40 ) | ( n_n48  &  n_n31 ) ;
 assign n_n197 = ( i_14_  &  (~ i_13_)  &  i_12_  &  wire899 ) ;
 assign wire89 = ( n_n282  &  _36112 ) | ( n_n282  &  _36113 ) ;
 assign n_n4094 = ( n_n53  &  wire89 ) | ( n_n222  &  wire901  &  n_n53 ) ;
 assign n_n47 = ( i_14_  &  i_13_  &  (~ i_12_)  &  wire900 ) ;
 assign wire67 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire914 ) | ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  wire914 ) ;
 assign n_n104 = ( i_14_  &  (~ i_13_)  &  i_12_  &  wire901 ) ;
 assign n_n4174 = ( n_n53  &  wire67 ) | ( n_n48  &  n_n104 ) ;
 assign wire407 = ( n_n264  &  n_n285  &  n_n282  &  n_n261 ) ;
 assign n_n247 = ( i_9_  &  (~ i_10_)  &  (~ i_11_) ) ;
 assign wire457 = ( n_n264  &  n_n285  &  n_n263  &  n_n247 ) ;
 assign n_n4153 = ( wire407 ) | ( wire457 ) | ( n_n53  &  n_n104 ) ;
 assign n_n4154 = ( wire72  &  n_n48 ) | ( wire905  &  n_n258  &  n_n48 ) ;
 assign wire456 = ( n_n220  &  wire905  &  n_n53 ) | ( wire905  &  n_n256  &  n_n53 ) ;
 assign wire4593 = ( wire66  &  n_n53 ) | ( wire905  &  n_n222  &  n_n53 ) ;
 assign wire20257 = ( n_n53  &  n_n107 ) | ( n_n53  &  n_n20 ) | ( n_n53  &  n_n19 ) ;
 assign wire20385 = ( n_n61  &  n_n53 ) | ( n_n108  &  n_n53 ) | ( n_n70  &  n_n53 ) ;
 assign n_n3964 = ( wire4593 ) | ( wire20257 ) | ( wire20385 ) ;
 assign n_n93 = ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire900 ) ;
 assign n_n46 = ( i_14_  &  i_13_  &  i_12_  &  wire906 ) ;
 assign n_n896 = ( n_n4  &  n_n47 ) | ( n_n4  &  n_n93 ) | ( n_n4  &  n_n46 ) ;
 assign n_n76 = ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  wire908 ) ;
 assign n_n29 = ( i_14_  &  i_13_  &  (~ i_12_)  &  wire908 ) ;
 assign wire49 = ( i_14_  &  (~ i_13_)  &  i_12_  &  wire902 ) | ( i_14_  &  i_13_  &  (~ i_12_)  &  wire902 ) ;
 assign wire460 = ( n_n57  &  wire88 ) | ( n_n57  &  n_n29 ) | ( n_n57  &  wire49 ) ;
 assign wire160 = ( n_n247  &  _35880 ) | ( n_n247  &  _35881 ) ;
 assign n_n252 = ( i_14_  &  (~ i_13_)  &  i_12_  &  wire904 ) ;
 assign wire409 = ( n_n3  &  _35389 ) | ( n_n3  &  wire904  &  _35391 ) ;
 assign n_n4920 = ( n_n57  &  wire79 ) | ( wire905  &  n_n57  &  n_n256 ) ;
 assign n_n4907 = ( n_n56  &  n_n108 ) | ( n_n57  &  wire70 ) ;
 assign n_n253 = ( i_9_  &  i_10_  &  i_11_ ) ;
 assign wire82 = ( i_14_  &  (~ i_13_)  &  i_12_  &  wire899 ) | ( i_14_  &  i_13_  &  (~ i_12_)  &  wire899 ) ;
 assign n_n15 = ( i_14_  &  i_13_  &  i_12_  &  wire898 ) ;
 assign wire635 = ( n_n56  &  wire44 ) | ( n_n56  &  n_n252 ) | ( n_n56  &  n_n15 ) ;
 assign wire42 = ( i_14_  &  i_13_  &  i_12_  &  wire905 ) | ( i_14_  &  i_13_  &  (~ i_12_)  &  wire905 ) ;
 assign wire636 = ( n_n56  &  wire42 ) | ( n_n279  &  n_n56  &  wire899 ) ;
 assign wire21065 = ( n_n57  &  n_n108 ) | ( n_n56  &  wire82 ) ;
 assign wire21070 = ( n_n4920 ) | ( n_n4907 ) | ( wire21066 ) ;
 assign wire539 = ( n_n281  &  n_n5  &  wire904 ) ;
 assign wire639 = ( n_n5  &  wire70 ) | ( n_n220  &  n_n5  &  wire898 ) ;
 assign wire3904 = ( n_n6  &  wire160 ) | ( n_n6  &  wire184 ) ;
 assign wire20950 = ( n_n5  &  _38123 ) | ( n_n5  &  wire904  &  _35427 ) ;
 assign n_n3172 = ( wire639 ) | ( wire3904 ) | ( wire20950 ) ;
 assign n_n4605 = ( n_n6  &  wire72 ) | ( n_n6  &  wire905  &  n_n258 ) ;
 assign wire20955 = ( n_n4605 ) | ( wire20952 ) | ( n_n5  &  wire208 ) ;
 assign wire20956 = ( n_n4815 ) | ( n_n4816 ) | ( wire3896 ) ;
 assign n_n3118 = ( n_n3172 ) | ( wire20955 ) | ( wire20956 ) ;
 assign n_n26 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire908 ) ;
 assign wire80 = ( n_n270  &  _35076 ) | ( n_n270  &  _35077 ) ;
 assign wire640 = ( n_n4  &  n_n76 ) | ( n_n4  &  n_n26 ) | ( n_n4  &  wire80 ) ;
 assign n_n80 = ( i_14_  &  i_13_  &  (~ i_12_)  &  wire902 ) ;
 assign wire3758 = ( _3343 ) | ( n_n3  &  _38155 ) | ( n_n3  &  _38156 ) ;
 assign wire21136 = ( wire640 ) | ( wire485 ) | ( n_n3  &  n_n76 ) ;
 assign wire453 = ( n_n247  &  _36098 ) | ( n_n247  &  _36099 ) ;
 assign n_n3259 = ( n_n1  &  wire453 ) | ( wire914  &  n_n1  &  n_n256 ) ;
 assign wire245 = ( n_n247  &  _36092 ) | ( n_n247  &  _36093 ) ;
 assign n_n3260 = ( n_n1  &  wire245 ) | ( n_n1  &  wire912  &  n_n225 ) ;
 assign wire61 = ( (~ i_14_)  &  i_13_  &  i_12_  &  wire902 ) | ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire902 ) ;
 assign n_n3772 = ( n_n1  &  wire61 ) | ( n_n1  &  n_n279  &  wire908 ) ;
 assign n_n3257 = ( n_n2  &  wire245 ) | ( n_n2  &  wire912  &  n_n225 ) ;
 assign wire20959 = ( n_n111  &  n_n1 ) | ( n_n1  &  wire453 ) | ( n_n1  &  n_n38 ) ;
 assign wire20962 = ( n_n3260 ) | ( n_n3772 ) | ( wire395 ) | ( wire5219 ) ;
 assign n_n3113 = ( wire20962 ) | ( _38103 ) ;
 assign n_n223 = ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire899 ) ;
 assign n_n2860 = ( _5435 ) | ( n_n1  &  wire42 ) | ( n_n1  &  n_n223 ) ;
 assign n_n3255 = ( n_n2  &  n_n76 ) | ( n_n1  &  wire82 ) ;
 assign wire814 = ( n_n1  &  n_n76 ) | ( n_n1  &  n_n26 ) | ( n_n1  &  wire80 ) ;
 assign wire3884 = ( n_n2  &  wire88 ) | ( n_n2  &  n_n29 ) | ( n_n2  &  wire49 ) ;
 assign wire71 = ( n_n253  &  _35150 ) | ( n_n253  &  _35151 ) ;
 assign wire68 = ( i_14_  &  (~ i_13_)  &  i_12_  &  wire898 ) | ( i_14_  &  i_13_  &  (~ i_12_)  &  wire898 ) ;
 assign wire496 = ( n_n2  &  n_n95 ) | ( n_n2  &  n_n49 ) | ( n_n2  &  wire71 ) ;
 assign n_n179 = ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire912 ) ;
 assign wire55 = ( n_n247  &  _36001 ) | ( n_n247  &  _36002 ) ;
 assign wire57 = ( n_n247  &  _35998 ) | ( n_n247  &  _35999 ) ;
 assign wire806 = ( n_n1  &  n_n179 ) | ( n_n1  &  wire55 ) | ( n_n1  &  wire57 ) ;
 assign n_n10 = ( i_14_  &  (~ i_13_)  &  i_12_  &  wire907 ) ;
 assign n_n100 = ( n_n260  &  n_n285  &  n_n261 ) ;
 assign wire19578 = ( n_n267  &  _35702 ) | ( n_n267  &  _35703 ) ;
 assign n_n1359 = ( n_n4  &  wire19578 ) | ( n_n4  &  n_n222  &  wire906 ) ;
 assign wire84 = ( (~ i_14_)  &  i_13_  &  i_12_  &  wire911 ) | ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire911 ) ;
 assign n_n3525 = ( n_n1  &  wire84 ) | ( wire913  &  n_n1  &  n_n279 ) ;
 assign n_n107 = ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  wire899 ) ;
 assign wire62 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire913 ) | ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  wire913 ) ;
 assign n_n204 = ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire911 ) ;
 assign n_n16 = ( (~ i_14_)  &  i_13_  &  i_12_  &  wire913 ) ;
 assign wire3358 = ( n_n5  &  wire62 ) | ( n_n279  &  n_n5  &  wire899 ) ;
 assign n_n4671 = ( n_n57  &  wire453 ) | ( wire914  &  n_n57  &  n_n256 ) ;
 assign wire252 = ( i_15_  &  n_n279  &  n_n282 ) | ( (~ i_15_)  &  n_n279  &  n_n282 ) ;
 assign wire329 = ( i_15_  &  n_n279  &  n_n247 ) | ( (~ i_15_)  &  n_n279  &  n_n247 ) ;
 assign wire21442 = ( n_n111  &  n_n57 ) | ( n_n56  &  n_n95 ) ;
 assign wire21443 = ( n_n56  &  wire252 ) | ( n_n57  &  wire329 ) ;
 assign n_n2169 = ( n_n4671 ) | ( wire21442 ) | ( wire21443 ) ;
 assign n_n66 = ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  wire904 ) ;
 assign wire164 = ( i_8_  &  n_n272  &  n_n285  &  n_n230 ) | ( (~ i_8_)  &  n_n272  &  n_n285  &  n_n230 ) ;
 assign wire985 = ( n_n281  &  wire914 ) | ( n_n281  &  wire903 ) ;
 assign wire3354 = ( n_n5  &  wire79 ) | ( n_n5  &  n_n109 ) | ( n_n5  &  wire83 ) ;
 assign wire21529 = ( n_n6  &  n_n12 ) | ( n_n5  &  n_n12 ) | ( n_n6  &  n_n66 ) | ( n_n5  &  n_n66 ) ;
 assign wire21533 = ( wire21530 ) | ( wire21531 ) | ( n_n106  &  wire164 ) ;
 assign wire333 = ( n_n220  &  wire905  &  n_n4 ) | ( wire905  &  n_n4  &  n_n256 ) ;
 assign wire3541 = ( wire48  &  n_n3 ) | ( n_n3  &  n_n204 ) | ( n_n3  &  n_n16 ) ;
 assign wire3542 = ( n_n4  &  wire79 ) | ( n_n279  &  wire905  &  n_n4 ) ;
 assign n_n171 = ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire897 ) ;
 assign n_n74 = ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  wire897 ) ;
 assign wire21367 = ( (~ i_14_)  &  i_13_  &  i_12_  &  wire903 ) | ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire903 ) ;
 assign n_n147 = ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  wire912 ) ;
 assign n_n94 = ( n_n260  &  n_n285  &  n_n263 ) ;
 assign n_n280 = ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  wire901 ) ;
 assign n_n32 = ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  wire907 ) ;
 assign n_n4165 = ( n_n216  &  n_n53 ) | ( n_n48  &  wire62 ) ;
 assign n_n42 = ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  wire906 ) ;
 assign wire81 = ( i_14_  &  (~ i_13_)  &  i_12_  &  wire900 ) | ( i_14_  &  i_13_  &  (~ i_12_)  &  wire900 ) ;
 assign wire69 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire908 ) | ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  wire908 ) ;
 assign n_n4624 = ( n_n6  &  n_n197 ) | ( n_n5  &  wire69 ) ;
 assign wire85 = ( i_14_  &  (~ i_13_)  &  i_12_  &  wire901 ) | ( i_14_  &  i_13_  &  (~ i_12_)  &  wire901 ) ;
 assign n_n1412 = ( n_n2  &  n_n32 ) | ( n_n1  &  wire85 ) ;
 assign n_n135 = ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  wire912 ) ;
 assign n_n41 = ( i_14_  &  (~ i_13_)  &  i_12_  &  wire912 ) ;
 assign wire347 = ( (~ i_15_)  &  n_n228  &  n_n247 ) | ( i_15_  &  n_n222  &  n_n247 ) | ( (~ i_15_)  &  n_n222  &  n_n247 ) ;
 assign n_n18 = ( i_14_  &  i_13_  &  i_12_  &  wire913 ) ;
 assign wire123 = ( i_14_  &  i_13_  &  i_12_  &  wire905 ) | ( i_14_  &  i_13_  &  (~ i_12_)  &  wire905 ) | ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire905 ) ;
 assign wire100 = ( (~ i_14_)  &  i_13_  &  i_12_  &  wire899 ) | ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire899 ) | ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  wire899 ) ;
 assign wire992 = ( wire60 ) | ( n_n18 ) | ( wire123 ) | ( wire100 ) ;
 assign n_n4858 = ( n_n111  &  n_n5 ) | ( n_n6  &  wire49 ) ;
 assign n_n4864 = ( n_n6  &  wire64 ) | ( wire907  &  n_n6  &  n_n279 ) ;
 assign wire102 = ( n_n247  &  _36974 ) | ( n_n247  &  _36975 ) ;
 assign n_n4635 = ( n_n5  &  wire102 ) | ( wire914  &  n_n279  &  n_n5 ) ;
 assign wire22106 = ( wire2703 ) | ( n_n5  &  wire102 ) | ( n_n5  &  n_n113 ) ;
 assign n_n4870 = ( n_n111  &  n_n6 ) | ( n_n5  &  wire85 ) ;
 assign wire78 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire907 ) | ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  wire907 ) ;
 assign n_n1497 = ( n_n6  &  n_n104 ) | ( n_n5  &  wire78 ) ;
 assign n_n1130 = ( n_n4870 ) | ( n_n1497 ) | ( _1588 ) | ( _39600 ) ;
 assign n_n22 = ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  wire903 ) ;
 assign wire897 = ( (~ i_9_)  &  (~ i_10_)  &  i_11_  &  i_15_ ) ;
 assign wire19407 = ( n_n275  &  _35114 ) | ( n_n275  &  _35115 ) ;
 assign n_n4852 = ( n_n5  &  wire19407 ) | ( n_n5  &  n_n256  &  wire897 ) ;
 assign n_n103 = ( i_14_  &  (~ i_13_)  &  i_12_  &  wire897 ) ;
 assign n_n1490 = ( n_n6  &  wire69 ) | ( n_n5  &  n_n103 ) ;
 assign wire140 = ( i_14_  &  i_13_  &  i_12_  &  wire908 ) | ( i_14_  &  i_13_  &  (~ i_12_)  &  wire908 ) | ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire908 ) ;
 assign wire346 = ( (~ i_15_)  &  n_n228  &  n_n275 ) | ( i_15_  &  n_n222  &  n_n275 ) | ( (~ i_15_)  &  n_n222  &  n_n275 ) ;
 assign wire998 = ( wire40 ) | ( n_n74 ) | ( wire140 ) | ( wire346 ) ;
 assign wire22119 = ( wire22117 ) | ( _1580 ) | ( _1583 ) | ( _1584 ) ;
 assign n_n1095 = ( wire22106 ) | ( n_n1130 ) | ( wire22119 ) | ( _39594 ) ;
 assign n_n1240 = ( wire461 ) | ( wire376 ) | ( wire2686 ) | ( wire22121 ) ;
 assign wire22129 = ( wire631 ) | ( wire22124 ) | ( wire22126 ) ;
 assign wire22130 = ( n_n4124 ) | ( wire2676 ) | ( wire22125 ) ;
 assign n_n1242 = ( n_n6879 ) | ( wire679 ) | ( wire2672 ) | ( wire2673 ) ;
 assign n_n1243 = ( wire2665 ) | ( wire22134 ) | ( wire22135 ) | ( wire22136 ) ;
 assign wire22142 = ( n_n4153 ) | ( wire2659 ) | ( wire22140 ) ;
 assign n_n1505 = ( n_n5  &  n_n54 ) | ( n_n6  &  wire51 ) ;
 assign wire22148 = ( n_n1506 ) | ( wire389 ) | ( n_n1505 ) ;
 assign wire22149 = ( wire2652 ) | ( _1534 ) | ( _1535 ) ;
 assign wire56 = ( i_14_  &  (~ i_13_)  &  i_12_  &  wire897 ) | ( i_14_  &  i_13_  &  (~ i_12_)  &  wire897 ) ;
 assign n_n1542 = ( n_n48  &  n_n22 ) | ( n_n53  &  wire56 ) ;
 assign n_n3827 = ( n_n48  &  wire61 ) | ( n_n279  &  wire908  &  n_n48 ) ;
 assign n_n1536 = ( wire60  &  n_n48 ) | ( n_n108  &  n_n53 ) ;
 assign wire22157 = ( wire624 ) | ( wire22154 ) | ( n_n48  &  wire69 ) ;
 assign n_n1135 = ( wire22157 ) | ( _1497 ) | ( _1498 ) | ( _39676 ) ;
 assign wire2638 = ( n_n48  &  wire22167 ) | ( n_n48  &  wire22168 ) ;
 assign wire22169 = ( n_n3581 ) | ( wire2637 ) | ( wire2640 ) | ( wire22160 ) ;
 assign wire22176 = ( n_n4168 ) | ( n_n1542 ) | ( wire2631 ) | ( wire22174 ) ;
 assign n_n1097 = ( n_n1135 ) | ( wire2638 ) | ( wire22169 ) | ( wire22176 ) ;
 assign wire368 = ( n_n247  &  _37013 ) | ( n_n247  &  _37014 ) ;
 assign n_n88 = ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  _36683 ) ;
 assign n_n1066 = ( n_n94  &  wire368 ) | ( n_n247  &  n_n94  &  _36683 ) ;
 assign n_n270 = ( i_9_  &  (~ i_10_)  &  i_11_ ) ;
 assign wire114 = ( i_15_  &  n_n225  &  n_n270 ) | ( (~ i_15_)  &  n_n225  &  n_n270 ) ;
 assign n_n275 = ( (~ i_9_)  &  (~ i_10_)  &  i_11_ ) ;
 assign wire120 = ( i_15_  &  n_n225  &  n_n275 ) | ( (~ i_15_)  &  n_n225  &  n_n275 ) ;
 assign wire459 = ( wire88  &  n_n94 ) | ( n_n31  &  n_n94 ) | ( n_n80  &  n_n94 ) ;
 assign wire22648 = ( n_n100  &  wire120 ) | ( n_n258  &  wire899  &  n_n100 ) ;
 assign n_n855 = ( wire459 ) | ( wire22648 ) | ( n_n94  &  wire114 ) ;
 assign wire19457 = ( n_n275  &  _35536 ) | ( n_n275  &  _35537 ) ;
 assign n_n3870 = ( n_n100  &  wire19457 ) | ( n_n222  &  n_n100  &  wire897 ) ;
 assign wire2091 = ( wire88  &  n_n100 ) | ( n_n80  &  n_n100 ) | ( n_n100  &  wire114 ) ;
 assign wire2092 = ( n_n94  &  wire19457 ) | ( n_n94  &  n_n25 ) | ( n_n94  &  wire22650 ) ;
 assign wire22654 = ( n_n3870 ) | ( wire22651 ) | ( wire22652 ) ;
 assign n_n772 = ( n_n855 ) | ( wire2091 ) | ( wire2092 ) | ( wire22654 ) ;
 assign n_n254 = ( i_13_  &  i_12_ ) ;
 assign wire301 = ( (~ i_14_)  &  i_15_  &  n_n282  &  n_n254 ) | ( i_14_  &  (~ i_15_)  &  n_n282  &  n_n254 ) | ( (~ i_14_)  &  (~ i_15_)  &  n_n282  &  n_n254 ) ;
 assign wire461 = ( n_n48  &  _38010 ) | ( n_n48  &  n_n247  &  _36683 ) ;
 assign wire2008 = ( n_n48  &  wire304 ) | ( n_n279  &  wire912  &  n_n48 ) ;
 assign wire19577 = ( i_14_  &  i_13_  &  (~ i_12_)  &  wire900 ) | ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire900 ) ;
 assign wire670 = ( n_n6  &  n_n105 ) | ( n_n6  &  n_n46 ) | ( n_n6  &  wire19577 ) ;
 assign wire2001 = ( n_n6  &  n_n99 ) | ( n_n6  &  wire96 ) | ( n_n6  &  wire134 ) ;
 assign wire2002 = ( n_n5  &  n_n46 ) | ( n_n5  &  wire19577 ) | ( n_n5  &  wire22719 ) ;
 assign n_n269 = ( i_9_  &  i_10_ ) ;
 assign n_n227 = ( n_n229  &  n_n285  &  n_n230 ) ;
 assign n_n207 = ( n_n208  &  n_n285  &  n_n230 ) ;
 assign n_n84 = ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire901 ) ;
 assign n_n142 = ( n_n260  &  n_n165  &  n_n273 ) ;
 assign n_n136 = ( n_n260  &  n_n165  &  n_n208 ) ;
 assign wire896 = ( i_5_  &  (~ i_3_)  &  i_4_  &  _34695 ) ;
 assign n_n278 = ( i_13_  &  (~ i_12_) ) ;
 assign n_n259 = ( i_9_  &  i_10_  &  (~ i_11_) ) ;
 assign n_n149 = ( (~ i_9_)  &  i_10_  &  i_12_  &  (~ i_11_) ) ;
 assign n_n122 = ( n_n264  &  n_n229  &  n_n165 ) ;
 assign n_n112 = ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire913 ) ;
 assign n_n212 = ( i_14_  &  i_13_  &  i_12_  &  wire903 ) ;
 assign n_n30 = ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire902 ) ;
 assign n_n221 = ( i_14_  &  i_13_  &  (~ i_12_)  &  wire899 ) ;
 assign n_n7 = ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  wire903 ) ;
 assign n_n144 = ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  wire899 ) ;
 assign n_n50 = ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  wire898 ) ;
 assign n_n267 = ( (~ i_9_)  &  i_10_  &  i_11_ ) ;
 assign n_n87 = ( i_14_  &  i_13_  &  i_12_  &  wire914 ) ;
 assign n_n34 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire901 ) ;
 assign n_n28 = ( (~ i_14_)  &  i_13_  &  i_12_  &  wire902 ) ;
 assign n_n75 = ( (~ i_14_)  &  i_13_  &  i_12_  &  wire897 ) ;
 assign n_n21 = ( i_14_  &  i_13_  &  i_12_  &  wire905 ) ;
 assign n_n17 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire911 ) ;
 assign n_n236 = ( i_14_  &  (~ i_13_)  &  i_12_  &  wire903 ) ;
 assign n_n40 = ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  _40255 ) ;
 assign n_n102 = ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire904 ) ;
 assign n_n33 = ( (~ i_14_)  &  i_13_  &  i_12_  &  wire907 ) ;
 assign n_n78 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire902 ) ;
 assign n_n200 = ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire903 ) ;
 assign n_n64 = ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  wire900 ) ;
 assign n_n150 = ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  wire911 ) ;
 assign n_n25 = ( i_14_  &  i_13_  &  (~ i_12_)  &  wire897 ) ;
 assign n_n24 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire897 ) ;
 assign n_n27 = ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  wire902 ) ;
 assign n_n20 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire899 ) ;
 assign n_n97 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire898 ) ;
 assign n_n52 = ( i_14_  &  i_13_  &  (~ i_12_)  &  wire904 ) ;
 assign n_n71 = ( (~ i_14_)  &  i_13_  &  i_12_  &  wire899 ) ;
 assign n_n69 = ( i_14_  &  i_13_  &  (~ i_12_)  &  _39255 ) ;
 assign n_n14 = ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  wire898 ) ;
 assign n_n63 = ( i_14_  &  i_13_  &  i_12_  &  wire901 ) ;
 assign n_n199 = ( i_14_  &  i_13_  &  (~ i_12_)  &  wire903 ) ;
 assign n_n92 = ( i_14_  &  i_13_  &  (~ i_12_)  &  wire906 ) ;
 assign n_n98 = ( i_14_  &  i_13_  &  i_12_  &  wire904 ) ;
 assign n_n38 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire914 ) ;
 assign n_n109 = ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire905 ) ;
 assign wire384 = ( n_n282  &  wire152 ) | ( n_n282  &  _34642 ) ;
 assign wire19205 = ( i_9_ ) | ( (~ i_9_)  &  i_10_ ) | ( (~ i_9_)  &  (~ i_10_)  &  i_11_ ) | ( (~ i_9_)  &  (~ i_10_)  &  i_12_  &  (~ i_11_) ) ;
 assign wire19239 = ( n_n270 ) | ( n_n281  &  wire905 ) ;
 assign wire5910 = ( (~ i_1_)  &  (~ i_2_)  &  (~ i_0_)  &  _34797 ) ;
 assign wire19207 = ( wire905  &  n_n258 ) | ( n_n258  &  wire904 ) ;
 assign wire19208 = ( i_11_  &  n_n256  &  n_n269 ) | ( (~ i_11_)  &  n_n256  &  n_n269 ) | ( i_11_  &  n_n269  &  wire288 ) | ( (~ i_11_)  &  n_n269  &  wire288 ) ;
 assign n_n5063 = ( wire5910 ) | ( n_n255  &  wire19207 ) | ( n_n255  &  wire19208 ) ;
 assign wire165 = ( (~ i_14_)  &  i_13_  &  i_12_  &  wire902 ) | ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire902 ) | ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  wire902 ) ;
 assign n_n4839 = ( n_n6  &  wire79 ) | ( n_n6  &  wire905  &  n_n256 ) ;
 assign wire53 = ( i_14_  &  i_13_  &  i_12_  &  wire903 ) | ( i_14_  &  i_13_  &  (~ i_12_)  &  wire903 ) ;
 assign n_n4960 = ( n_n285  &  n_n266  &  n_n230  &  wire180 ) ;
 assign n_n4954 = ( n_n57  &  wire55 ) | ( n_n279  &  wire912  &  n_n57 ) ;
 assign n_n4953 = ( n_n57  &  wire57 ) | ( wire914  &  n_n279  &  n_n57 ) ;
 assign n_n4955 = ( n_n56  &  n_n95 ) | ( n_n56  &  n_n49 ) | ( n_n56  &  n_n96 ) ;
 assign wire671 = ( n_n56  &  wire99 ) | ( n_n56  &  wire41 ) ;
 assign wire20705 = ( n_n57  &  wire153 ) | ( n_n56  &  wire254 ) ;
 assign wire20706 = ( wire273  &  n_n57 ) | ( n_n57  &  wire180 ) ;
 assign wire20710 = ( n_n4954 ) | ( n_n4953 ) | ( n_n4955 ) | ( wire671 ) ;
 assign wire469 = ( n_n259  &  _37043 ) | ( n_n259  &  _37044 ) ;
 assign n_n4073 = ( n_n53  &  wire469 ) | ( n_n222  &  wire899  &  n_n53 ) ;
 assign wire475 = ( n_n53  &  _37840 ) | ( wire899  &  n_n53  &  _35953 ) ;
 assign n_n4068 = ( n_n9  &  n_n53 ) | ( n_n145  &  n_n53 ) | ( n_n53  &  n_n144 ) ;
 assign n_n4069 = ( n_n60  &  n_n53 ) | ( n_n8  &  n_n53 ) | ( n_n226  &  n_n53 ) ;
 assign wire77 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire904 ) | ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  wire904 ) ;
 assign n_n1363 = ( n_n105  &  n_n3 ) | ( n_n4  &  wire77 ) ;
 assign wire184 = ( n_n247  &  _34581 ) | ( n_n247  &  _34582 ) ;
 assign n_n3324 = ( n_n9  &  n_n57 ) | ( n_n56  &  wire184 ) ;
 assign n_n6504 = ( wire912  &  n_n258  &  n_n48 ) ;
 assign n_n1633 = ( n_n197  &  n_n100 ) | ( n_n94  &  wire69 ) ;
 assign n_n4923 = ( n_n56  &  n_n76 ) | ( n_n57  &  wire82 ) ;
 assign wire21073 = ( n_n4923 ) | ( n_n4924 ) | ( wire5544 ) ;
 assign wire21074 = ( n_n4922 ) | ( n_n4921 ) | ( wire21072 ) ;
 assign n_n3130 = ( wire21073 ) | ( wire21074 ) | ( _4160 ) | ( _4161 ) ;
 assign wire686 = ( wire912  &  n_n225  &  n_n94 ) | ( wire912  &  n_n256  &  n_n94 ) ;
 assign wire825 = ( n_n247  &  _35998  &  _38131 ) | ( n_n247  &  _35999  &  _38131 ) ;
 assign wire20973 = ( n_n4  &  n_n31 ) | ( n_n147  &  n_n94 ) ;
 assign wire20974 = ( n_n94  &  _38132 ) | ( n_n247  &  n_n94  &  _36683 ) ;
 assign wire20975 = ( n_n11  &  n_n94 ) | ( n_n94  &  n_n86 ) | ( n_n94  &  n_n39 ) ;
 assign n_n3167 = ( wire825 ) | ( wire20973 ) | ( wire20974 ) | ( wire20975 ) ;
 assign wire278 = ( i_8_  &  n_n231  &  n_n285  &  n_n230 ) | ( (~ i_8_)  &  n_n231  &  n_n285  &  n_n230 ) ;
 assign wire1018 = ( n_n228  &  wire902 ) | ( wire905  &  n_n258 ) ;
 assign wire20984 = ( wire20981 ) | ( wire20982 ) | ( wire278  &  wire1018 ) ;
 assign n_n3117 = ( n_n3167 ) | ( wire20984 ) | ( _3358 ) | ( _38142 ) ;
 assign n_n3242 = ( n_n4  &  wire245 ) | ( n_n4  &  wire912  &  n_n225 ) ;
 assign wire557 = ( n_n3  &  n_n95 ) | ( n_n3  &  n_n49 ) | ( n_n3  &  wire71 ) ;
 assign wire3754 = ( _3327 ) | ( _3328 ) | ( _3329 ) ;
 assign n_n3757 = ( n_n1  &  wire63 ) | ( n_n281  &  n_n1  &  wire908 ) ;
 assign wire739 = ( n_n228  &  n_n2  &  wire899 ) ;
 assign wire20931 = ( n_n2618 ) | ( n_n3757 ) | ( wire739 ) | ( wire3931 ) ;
 assign wire20933 = ( n_n4  &  n_n95 ) | ( n_n268  &  n_n148 ) ;
 assign wire20934 = ( n_n4  &  wire68 ) | ( n_n3  &  wire68 ) ;
 assign wire20936 = ( wire3924 ) | ( _3300 ) ;
 assign wire20938 = ( n_n1  &  n_n108 ) | ( n_n2  &  wire82 ) ;
 assign n_n3519 = ( n_n2  &  n_n108 ) | ( n_n1  &  wire70 ) ;
 assign n_n3520 = ( n_n2  &  wire79 ) | ( n_n2  &  wire905  &  n_n256 ) ;
 assign n_n148 = ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  wire914 ) ;
 assign n_n81 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire907 ) ;
 assign wire470 = ( n_n53  &  _37110 ) | ( wire907  &  n_n53  &  _36856 ) ;
 assign n_n3019 = ( n_n53  &  n_n280 ) | ( n_n53  &  n_n33 ) | ( n_n53  &  n_n81 ) ;
 assign n_n2986 = ( n_n4  &  wire79 ) | ( n_n4  &  wire899  &  n_n256 ) ;
 assign n_n3524 = ( n_n1  &  wire19738 ) | ( wire913  &  n_n1  &  n_n256 ) ;
 assign wire185 = ( i_8_  &  n_n264  &  n_n285  &  n_n155 ) | ( (~ i_8_)  &  n_n264  &  n_n285  &  n_n155 ) ;
 assign wire3310 = ( n_n281  &  wire907  &  wire185 ) ;
 assign wire21560 = ( n_n281  &  wire905  &  n_n53 ) | ( n_n281  &  wire908  &  n_n53 ) ;
 assign wire21561 = ( n_n281  &  wire914  &  n_n48 ) | ( n_n281  &  wire914  &  n_n53 ) ;
 assign wire21562 = ( n_n60  &  n_n48 ) | ( n_n48  &  n_n7 ) | ( n_n53  &  n_n7 ) ;
 assign n_n2148 = ( wire3310 ) | ( wire21560 ) | ( wire21561 ) | ( wire21562 ) ;
 assign n_n19 = ( (~ i_14_)  &  i_13_  &  i_12_  &  wire905 ) ;
 assign n_n2272 = ( n_n108  &  n_n53 ) | ( n_n70  &  n_n53 ) | ( n_n53  &  n_n19 ) ;
 assign wire3491 = ( n_n2  &  n_n84 ) | ( n_n2  &  n_n35 ) | ( n_n2  &  wire86 ) ;
 assign wire21417 = ( n_n281  &  wire905  &  n_n53 ) | ( n_n281  &  wire908  &  n_n53 ) ;
 assign n_n2126 = ( n_n2272 ) | ( wire3491 ) | ( wire21417 ) ;
 assign wire135 = ( i_8_  &  n_n260  &  n_n285  &  n_n155 ) | ( (~ i_8_)  &  n_n260  &  n_n285  &  n_n155 ) ;
 assign wire264 = ( i_15_  &  n_n279  &  n_n275 ) | ( (~ i_15_)  &  n_n279  &  n_n275 ) ;
 assign wire1031 = ( n_n281  &  wire905 ) | ( n_n281  &  wire908 ) ;
 assign wire1030 = ( wire913  &  n_n281 ) | ( n_n281  &  wire903 ) ;
 assign wire466 = ( n_n220  &  n_n4  &  wire908 ) | ( n_n4  &  wire908  &  n_n256 ) ;
 assign wire3533 = ( n_n3  &  wire67 ) | ( n_n279  &  n_n3  &  wire897 ) ;
 assign wire3534 = ( n_n4  &  wire80 ) | ( n_n279  &  n_n4  &  wire908 ) ;
 assign wire21374 = ( n_n4  &  n_n76 ) | ( n_n4  &  n_n26 ) | ( n_n4  &  n_n30 ) ;
 assign n_n2104 = ( wire3533 ) | ( wire3534 ) | ( wire21374 ) ;
 assign wire411 = ( n_n220  &  n_n6  &  wire905 ) | ( n_n6  &  wire905  &  n_n256 ) ;
 assign wire3344 = ( wire48  &  n_n5 ) | ( n_n5  &  n_n204 ) | ( n_n5  &  n_n16 ) ;
 assign wire3345 = ( n_n6  &  wire79 ) | ( n_n6  &  n_n279  &  wire905 ) ;
 assign n_n2137 = ( wire411 ) | ( wire3344 ) | ( wire3345 ) ;
 assign wire21381 = ( n_n4  &  n_n186 ) | ( n_n268  &  n_n148 ) ;
 assign n_n2110 = ( wire21381 ) | ( _2766 ) | ( n_n265  &  _38639 ) ;
 assign wire21387 = ( wire3520 ) | ( wire21385 ) | ( n_n268  &  n_n22 ) ;
 assign wire3518 = ( n_n4  &  wire51 ) | ( n_n4  &  n_n90 ) | ( n_n4  &  wire21389 ) ;
 assign wire21390 = ( n_n3  &  wire51 ) | ( n_n4  &  n_n93 ) ;
 assign wire476 = ( n_n220  &  n_n3  &  wire904 ) | ( n_n3  &  n_n256  &  wire904 ) ;
 assign wire104 = ( n_n275  &  _35629 ) | ( n_n275  &  _35630 ) ;
 assign wire228 = ( n_n275  &  _39072 ) | ( n_n275  &  _39073 ) ;
 assign wire21842 = ( n_n53  &  n_n76 ) | ( n_n53  &  n_n25 ) | ( n_n53  &  n_n27 ) ;
 assign n_n58 = ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  wire897 ) ;
 assign wire667 = ( n_n247  &  n_n94  &  _39057 ) | ( n_n247  &  n_n94  &  _39059 ) ;
 assign wire696 = ( n_n281  &  wire911  &  n_n94 ) | ( wire911  &  n_n225  &  n_n94 ) ;
 assign wire21686 = ( n_n94  &  _39063 ) | ( n_n222  &  n_n94  &  _36699 ) ;
 assign wire21687 = ( n_n94  &  n_n58 ) | ( n_n94  &  n_n86 ) | ( n_n94  &  n_n39 ) ;
 assign n_n1757 = ( wire667 ) | ( wire696 ) | ( wire21686 ) | ( wire21687 ) ;
 assign n_n3581 = ( n_n53  &  wire84 ) | ( wire913  &  n_n279  &  n_n53 ) ;
 assign wire143 = ( n_n259  &  _38136 ) | ( n_n259  &  _38137 ) ;
 assign wire306 = ( n_n259  &  _38140 ) | ( n_n259  &  _38141 ) ;
 assign wire22079 = ( n_n70  &  n_n227 ) | ( n_n257  &  n_n207 ) ;
 assign n_n1215 = ( wire22079 ) | ( _1292 ) | ( n_n207  &  _39860 ) ;
 assign wire514 = ( (~ i_15_)  &  n_n242  &  n_n279 ) | ( (~ i_15_)  &  n_n242  &  n_n222 ) ;
 assign n_n1628 = ( n_n94  &  wire514 ) | ( wire911  &  n_n225  &  n_n94 ) ;
 assign wire52 = ( (~ i_15_)  &  n_n228  &  n_n242 ) | ( (~ i_15_)  &  n_n242  &  n_n222 ) ;
 assign n_n2732 = ( n_n100  &  wire52 ) | ( wire913  &  n_n279  &  n_n100 ) ;
 assign n_n1624 = ( n_n100  &  wire62 ) | ( n_n197  &  n_n94 ) ;
 assign wire247 = ( (~ i_14_)  &  i_13_  &  i_12_  &  wire911 ) | ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire911 ) | ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  wire911 ) ;
 assign wire83 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire905 ) | ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  wire905 ) ;
 assign wire1044 = ( wire60 ) | ( n_n107 ) | ( wire247 ) | ( wire83 ) ;
 assign wire175 = ( i_15_  &  n_n256  &  n_n253 ) | ( (~ i_15_)  &  n_n256  &  n_n253 ) ;
 assign wire579 = ( n_n264  &  n_n285  &  n_n242  &  n_n261 ) ;
 assign wire764 = ( n_n264  &  n_n285  &  n_n263  &  n_n259 ) ;
 assign wire2542 = ( n_n56  &  n_n240 ) | ( n_n56  &  wire63 ) | ( n_n56  &  wire50 ) ;
 assign wire2543 = ( n_n57  &  wire223 ) | ( n_n57  &  wire22259 ) ;
 assign wire699 = ( n_n6  &  wire66 ) | ( n_n6  &  wire899  &  n_n256 ) ;
 assign wire22020 = ( n_n4834 ) | ( wire411 ) | ( wire2784 ) ;
 assign n_n1320 = ( n_n110  &  n_n4 ) | ( n_n3  &  wire82 ) ;
 assign wire376 = ( n_n220  &  wire907  &  n_n53 ) | ( wire907  &  n_n256  &  n_n53 ) ;
 assign wire2686 = ( wire64  &  n_n53 ) | ( wire907  &  n_n279  &  n_n53 ) ;
 assign wire22121 = ( n_n53  &  n_n280 ) | ( n_n48  &  n_n87 ) ;
 assign n_n4124 = ( n_n48  &  wire102 ) | ( wire914  &  n_n279  &  n_n48 ) ;
 assign wire629 = ( n_n281  &  wire912  &  n_n48 ) | ( wire912  &  n_n256  &  n_n48 ) ;
 assign n_n62 = ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  wire901 ) ;
 assign wire631 = ( n_n48  &  n_n147 ) | ( n_n53  &  n_n62 ) ;
 assign n_n6879 = ( wire905  &  n_n258  &  n_n53 ) ;
 assign wire679 = ( n_n8  &  n_n48 ) | ( n_n53  &  n_n144 ) ;
 assign wire2672 = ( wire75  &  n_n48 ) | ( n_n258  &  wire908  &  n_n48 ) ;
 assign wire2673 = ( n_n53  &  wire50 ) | ( wire913  &  n_n258  &  n_n53 ) ;
 assign wire2665 = ( n_n275  &  _35036  &  _39632 ) | ( n_n275  &  _35037  &  _39632 ) ;
 assign wire22134 = ( n_n53  &  _39633 ) | ( wire908  &  n_n53  &  _35046 ) ;
 assign wire22135 = ( n_n246  &  n_n48 ) | ( n_n53  &  n_n10 ) ;
 assign wire22136 = ( n_n48  &  n_n147 ) | ( n_n48  &  n_n62 ) | ( n_n53  &  n_n62 ) ;
 assign wire223 = ( n_n259  &  _39426 ) | ( n_n259  &  _39427 ) ;
 assign wire168 = ( i_8_  &  n_n260  &  n_n272  &  n_n285 ) | ( (~ i_8_)  &  n_n260  &  n_n272  &  n_n285 ) ;
 assign wire128 = ( i_15_  &  n_n225  &  n_n259 ) | ( (~ i_15_)  &  n_n225  &  n_n259 ) ;
 assign wire22605 = ( n_n65  &  n_n100 ) | ( n_n15  &  n_n100 ) | ( n_n65  &  n_n94 ) ;
 assign n_n203 = ( i_14_  &  i_13_  &  (~ i_12_)  &  _36699 ) ;
 assign n_n1058 = ( n_n204  &  n_n94 ) | ( n_n94  &  n_n18 ) | ( n_n94  &  n_n203 ) ;
 assign wire20149 = ( (~ i_15_)  &  n_n228  &  n_n242 ) | ( i_15_  &  n_n242  &  n_n279 ) ;
 assign n_n3604 = ( n_n100  &  wire20149 ) | ( n_n222  &  n_n100  &  _36699 ) ;
 assign n_n3610 = ( n_n100  &  wire469 ) | ( n_n222  &  wire899  &  n_n100 ) ;
 assign wire697 = ( wire913  &  n_n225  &  n_n94 ) | ( wire911  &  n_n225  &  n_n94 ) ;
 assign wire1061 = ( i_15_  &  n_n242  &  n_n225 ) | ( (~ i_15_)  &  n_n242  &  n_n225 ) | ( i_15_  &  n_n225  &  n_n259 ) | ( (~ i_15_)  &  n_n225  &  n_n259 ) ;
 assign wire22610 = ( wire697 ) | ( n_n216  &  n_n100 ) | ( n_n100  &  wire1061 ) ;
 assign wire22611 = ( n_n1058 ) | ( n_n3604 ) | ( n_n3610 ) | ( wire22606 ) ;
 assign n_n771 = ( wire22605 ) | ( wire22610 ) | ( wire22611 ) | ( _290 ) ;
 assign wire516 = ( n_n258  &  wire901  &  n_n53 ) | ( n_n222  &  wire901  &  n_n53 ) ;
 assign wire1062 = ( n_n279  &  wire901 ) | ( n_n228  &  wire897 ) ;
 assign wire1997 = ( n_n228  &  wire902  &  n_n48 ) ;
 assign wire22725 = ( n_n228  &  wire899  &  n_n48 ) | ( n_n228  &  wire899  &  n_n53 ) ;
 assign wire22727 = ( n_n206  &  n_n48 ) | ( n_n206  &  n_n53 ) | ( n_n53  &  wire1062 ) ;
 assign n_n825 = ( wire516 ) | ( wire1997 ) | ( wire22725 ) | ( wire22727 ) ;
 assign wire675 = ( n_n228  &  wire898  &  n_n48 ) ;
 assign wire310 = ( n_n228  &  wire912 ) | ( n_n228  &  wire897 ) ;
 assign wire1064 = ( n_n221 ) | ( wire469 ) | ( wire128 ) | ( wire310 ) ;
 assign wire1063 = ( n_n228  &  wire901 ) | ( n_n228  &  wire900 ) ;
 assign wire1990 = ( n_n53  &  wire161 ) | ( n_n53  &  wire22730 ) ;
 assign wire22731 = ( n_n9  &  n_n53 ) | ( n_n48  &  n_n15 ) ;
 assign wire22734 = ( wire22732 ) | ( n_n48  &  wire1064 ) ;
 assign n_n762 = ( n_n825 ) | ( wire1990 ) | ( wire22731 ) | ( wire22734 ) ;
 assign n_n13 = ( i_14_  &  (~ i_13_)  &  i_12_  &  wire906 ) ;
 assign wire2436 = ( n_n100  &  wire110 ) | ( n_n258  &  wire904  &  n_n100 ) ;
 assign wire2437 = ( n_n94  &  wire123 ) | ( n_n94  &  wire187 ) ;
 assign n_n458 = ( wire2436 ) | ( wire2437 ) | ( n_n197  &  n_n94 ) ;
 assign wire1066 = ( wire914  &  n_n258 ) | ( n_n258  &  wire908 ) ;
 assign wire22372 = ( n_n2732 ) | ( wire22369 ) | ( wire22370 ) ;
 assign n_n374 = ( n_n458 ) | ( wire22372 ) | ( _995 ) | ( _40115 ) ;
 assign wire486 = ( i_14_  &  i_13_  &  i_12_  &  wire904 ) | ( i_14_  &  i_13_  &  (~ i_12_)  &  wire904 ) ;
 assign wire658 = ( n_n256  &  wire903  &  n_n94 ) | ( n_n256  &  n_n94  &  wire897 ) ;
 assign n_n707 = ( n_n94  &  n_n212 ) | ( n_n94  &  n_n200 ) | ( n_n94  &  n_n199 ) ;
 assign wire2410 = ( n_n100  &  n_n270  &  _40140 ) | ( n_n100  &  n_n270  &  _40142 ) ;
 assign wire22384 = ( n_n258  &  n_n100  &  wire897 ) | ( n_n258  &  n_n94  &  wire897 ) ;
 assign n_n462 = ( wire658 ) | ( n_n707 ) | ( wire2410 ) | ( wire22384 ) ;
 assign wire1069 = ( i_15_  &  n_n258  &  n_n270 ) | ( i_15_  &  n_n256  &  n_n270 ) | ( (~ i_15_)  &  n_n256  &  n_n270 ) ;
 assign wire22383 = ( wire2425 ) | ( wire2426 ) | ( wire2427 ) | ( wire2428 ) ;
 assign n_n346 = ( n_n374 ) | ( n_n462 ) | ( _40160 ) | ( _40161 ) ;
 assign n_n43 = ( (~ i_14_)  &  i_13_  &  i_12_  &  wire906 ) ;
 assign n_n82 = ( (~ i_14_)  &  i_13_  &  i_12_  &  wire901 ) ;
 assign n_n68 = ( (~ i_14_)  &  i_13_  &  i_12_  &  wire911 ) ;
 assign n_n113 = ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire914 ) ;
 assign n_n86 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire912 ) ;
 assign n_n79 = ( i_14_  &  i_13_  &  i_12_  &  wire908 ) ;
 assign n_n36 = ( i_14_  &  i_13_  &  i_12_  &  wire907 ) ;
 assign n_n44 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire900 ) ;
 assign n_n73 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire903 ) ;
 assign wire19265 = ( n_n225  &  n_n270 ) | ( n_n220  &  n_n275 ) ;
 assign wire19266 = ( wire19264 ) | ( n_n258  &  wire899 ) ;
 assign wire19267 = ( n_n228  &  wire908 ) | ( n_n259  &  wire148 ) ;
 assign wire1071 = ( wire19265 ) | ( wire19266 ) | ( wire19267 ) ;
 assign wire277 = ( i_14_  &  (~ i_13_)  &  i_12_  &  wire901 ) | ( i_14_  &  i_13_  &  (~ i_12_)  &  wire901 ) | ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire901 ) ;
 assign n_n4924 = ( n_n56  &  wire80 ) | ( n_n56  &  wire908  &  n_n256 ) ;
 assign wire255 = ( (~ i_14_)  &  i_13_  &  i_12_  &  wire904 ) | ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire904 ) | ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  wire904 ) ;
 assign n_n4871 = ( n_n285  &  n_n230  &  n_n263  &  wire255 ) ;
 assign n_n4838 = ( n_n6  &  n_n108 ) | ( n_n5  &  wire60 ) ;
 assign wire19896 = ( n_n4842 ) | ( n_n4839 ) | ( wire5054 ) ;
 assign n_n4730 = ( wire19896 ) | ( _5164 ) | ( _5165 ) | ( _36495 ) ;
 assign wire1076 = ( n_n229  &  n_n165  &  n_n284 ) | ( n_n165  &  n_n284  &  n_n283 ) ;
 assign wire1079 = ( n_n264  &  n_n229  &  n_n165 ) | ( n_n264  &  n_n165  &  n_n271 ) ;
 assign wire632 = ( n_n6  &  n_n258  &  wire898 ) | ( n_n6  &  wire898  &  n_n222 ) ;
 assign wire5368 = ( wire118  &  n_n56 ) | ( n_n56  &  n_n145 ) | ( n_n56  &  n_n144 ) ;
 assign wire5369 = ( n_n6  &  wire96 ) | ( n_n6  &  n_n222  &  wire904 ) ;
 assign n_n4330 = ( wire632 ) | ( wire5368 ) | ( wire5369 ) ;
 assign wire5361 = ( n_n6  &  wire71 ) | ( n_n6  &  n_n102 ) | ( n_n6  &  wire807 ) ;
 assign wire5363 = ( n_n151  &  n_n57 ) | ( wire75  &  n_n57 ) | ( n_n57  &  wire19668 ) ;
 assign wire19671 = ( wire5362 ) | ( wire19669 ) | ( n_n5  &  wire81 ) ;
 assign n_n4806 = ( n_n151  &  n_n6 ) | ( wire118  &  n_n5 ) ;
 assign n_n101 = ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire908 ) ;
 assign wire65 = ( i_14_  &  i_13_  &  (~ i_12_)  &  wire908 ) | ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire908 ) ;
 assign n_n1341 = ( n_n4  &  wire65 ) | ( n_n4  &  wire902  &  n_n225 ) ;
 assign wire4602 = ( n_n53  &  n_n34 ) | ( n_n53  &  n_n82 ) | ( n_n53  &  wire47 ) ;
 assign n_n3974 = ( n_n6504 ) | ( wire470 ) | ( wire376 ) | ( wire4602 ) ;
 assign n_n4090 = ( n_n48  &  wire368 ) | ( n_n48  &  n_n247  &  _36683 ) ;
 assign wire462 = ( n_n220  &  wire914  &  n_n48 ) | ( wire914  &  n_n256  &  n_n48 ) ;
 assign wire464 = ( n_n48  &  _37116 ) | ( wire914  &  n_n48  &  _36977 ) ;
 assign wire20330 = ( wire631 ) | ( wire462 ) | ( wire464 ) | ( wire20323 ) ;
 assign wire20331 = ( n_n4124 ) | ( n_n4090 ) | ( wire20324 ) | ( wire20325 ) ;
 assign wire1089 = ( wire75 ) | ( n_n206 ) | ( wire208 ) | ( wire199 ) ;
 assign wire20340 = ( wire4520 ) | ( wire20334 ) | ( wire20337 ) ;
 assign wire20341 = ( n_n4094 ) | ( wire20336 ) | ( n_n48  &  wire1089 ) ;
 assign n_n3506 = ( n_n4  &  wire42 ) | ( n_n279  &  n_n4  &  wire899 ) ;
 assign wire4302 = ( n_n4  &  wire66 ) | ( n_n4  &  wire79 ) | ( n_n4  &  n_n20 ) ;
 assign wire455 = ( n_n4  &  n_n258  &  wire900 ) | ( n_n4  &  n_n222  &  wire900 ) ;
 assign wire485 = ( n_n4  &  n_n258  &  wire899 ) | ( n_n4  &  n_n222  &  wire899 ) ;
 assign wire76 = ( i_14_  &  i_13_  &  i_12_  &  wire906 ) | ( i_14_  &  i_13_  &  (~ i_12_)  &  wire906 ) ;
 assign n_n3781 = ( n_n1  &  wire76 ) | ( n_n1  &  n_n279  &  wire900 ) ;
 assign wire676 = ( n_n53  &  _37326 ) | ( wire899  &  n_n53  &  _37091 ) ;
 assign wire21006 = ( n_n48  &  _38025 ) | ( wire899  &  n_n48  &  _37091 ) ;
 assign n_n3184 = ( n_n4154 ) | ( wire475 ) | ( wire676 ) | ( wire21006 ) ;
 assign wire96 = ( n_n253  &  _35142 ) | ( n_n253  &  _35143 ) ;
 assign wire712 = ( n_n54  &  n_n3 ) | ( n_n3  &  n_n99 ) | ( n_n3  &  wire96 ) ;
 assign wire4472 = ( n_n4  &  wire80 ) | ( n_n4  &  wire902  &  n_n256 ) ;
 assign wire20397 = ( n_n4  &  n_n197 ) | ( n_n4  &  n_n76 ) | ( n_n4  &  n_n26 ) ;
 assign wire20400 = ( n_n1341 ) | ( n_n884 ) | ( n_n876 ) | ( wire4478 ) ;
 assign wire20987 = ( wire333 ) | ( n_n2986 ) | ( wire712 ) ;
 assign n_n3116 = ( wire4472 ) | ( wire20397 ) | ( wire20400 ) | ( wire20987 ) ;
 assign n_n35 = ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire907 ) ;
 assign n_n4922 = ( n_n57  &  wire42 ) | ( n_n279  &  n_n57  &  wire899 ) ;
 assign n_n4921 = ( n_n57  &  wire66 ) | ( n_n57  &  wire899  &  n_n256 ) ;
 assign n_n4076 = ( n_n53  &  wire65 ) | ( wire902  &  n_n225  &  n_n53 ) ;
 assign n_n3768 = ( n_n1  &  wire19407 ) | ( n_n1  &  n_n256  &  wire897 ) ;
 assign wire484 = ( n_n220  &  n_n57  &  wire904 ) | ( n_n57  &  n_n256  &  wire904 ) ;
 assign wire21303 = ( wire372 ) | ( wire386 ) | ( wire894 ) | ( wire484 ) ;
 assign n_n2439 = ( wire21303 ) | ( _3064 ) | ( _38379 ) | ( _38386 ) ;
 assign wire21603 = ( n_n12  &  n_n48 ) | ( n_n12  &  n_n53 ) | ( n_n53  &  n_n66 ) ;
 assign n_n4912 = ( n_n57  &  wire19738 ) | ( wire913  &  n_n57  &  n_n256 ) ;
 assign n_n4916 = ( n_n56  &  wire19738 ) | ( wire913  &  n_n56  &  n_n256 ) ;
 assign wire327 = ( i_15_  &  n_n242  &  n_n279 ) | ( (~ i_15_)  &  n_n242  &  n_n279 ) ;
 assign wire1094 = ( i_8_  &  n_n153  &  n_n285  &  n_n230 ) | ( (~ i_8_)  &  n_n153  &  n_n285  &  n_n230 ) ;
 assign wire191 = ( i_8_  &  n_n153  &  n_n285  &  n_n230 ) | ( (~ i_8_)  &  n_n153  &  n_n285  &  n_n230 ) ;
 assign wire1096 = ( n_n281  &  wire906 ) | ( n_n281  &  wire904 ) ;
 assign wire1095 = ( n_n281  &  wire914 ) | ( n_n281  &  wire906 ) | ( n_n281  &  wire904 ) ;
 assign wire167 = ( (~ i_14_)  &  i_13_  &  i_12_  &  wire908 ) | ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire908 ) | ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  wire908 ) ;
 assign wire210 = ( (~ i_14_)  &  i_13_  &  i_12_  &  wire913 ) | ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire913 ) | ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  wire913 ) ;
 assign wire235 = ( i_15_  &  n_n281  &  n_n270 ) | ( i_15_  &  n_n279  &  n_n270 ) | ( (~ i_15_)  &  n_n279  &  n_n270 ) ;
 assign wire399 = ( i_15_  &  n_n281  &  n_n242 ) | ( i_15_  &  n_n242  &  n_n279 ) | ( (~ i_15_)  &  n_n242  &  n_n279 ) ;
 assign wire1097 = ( wire167 ) | ( wire210 ) | ( wire235 ) | ( wire399 ) ;
 assign wire436 = ( i_15_  &  n_n281  &  n_n282 ) | ( i_15_  &  n_n279  &  n_n282 ) | ( (~ i_15_)  &  n_n279  &  n_n282 ) ;
 assign wire1102 = ( wire268 ) | ( wire167 ) | ( wire235 ) | ( wire436 ) ;
 assign wire641 = ( n_n4  &  _39067 ) | ( n_n4  &  wire902  &  _39044 ) ;
 assign wire3145 = ( n_n4  &  wire61 ) | ( n_n4  &  n_n222  &  wire908 ) ;
 assign wire21690 = ( n_n4  &  n_n80 ) | ( n_n147  &  n_n94 ) ;
 assign wire21691 = ( n_n4  &  n_n221 ) | ( n_n94  &  n_n150 ) ;
 assign n_n1756 = ( wire641 ) | ( wire3145 ) | ( wire21690 ) | ( wire21691 ) ;
 assign wire50 = ( n_n275  &  _35036 ) | ( n_n275  &  _35037 ) ;
 assign wire645 = ( n_n100  &  _39746 ) | ( wire901  &  n_n100  &  _35946 ) ;
 assign wire2596 = ( wire63  &  n_n100 ) | ( n_n258  &  wire903  &  n_n100 ) ;
 assign wire2597 = ( n_n275  &  _35036  &  _39749 ) | ( n_n275  &  _35037  &  _39749 ) ;
 assign wire22203 = ( n_n94  &  _39750 ) | ( wire914  &  n_n94  &  _37163 ) ;
 assign n_n1286 = ( wire645 ) | ( wire2596 ) | ( wire2597 ) | ( wire22203 ) ;
 assign wire2593 = ( wire73  &  n_n100 ) | ( n_n100  &  wire220 ) | ( n_n100  &  wire22206 ) ;
 assign wire2594 = ( n_n94  &  wire22210 ) | ( n_n94  &  wire22211 ) ;
 assign wire2516 = ( n_n53  &  n_n82 ) | ( n_n53  &  wire144 ) | ( n_n53  &  wire47 ) ;
 assign wire22280 = ( n_n53  &  _39502 ) | ( wire907  &  n_n53  &  _36212 ) ;
 assign n_n1255 = ( wire461 ) | ( wire2516 ) | ( wire22280 ) ;
 assign n_n6848 = ( wire902  &  n_n258  &  n_n53 ) ;
 assign wire479 = ( n_n220  &  wire908  &  n_n53 ) | ( wire908  &  n_n256  &  n_n53 ) ;
 assign wire656 = ( wire902  &  n_n222  &  n_n53 ) | ( n_n222  &  wire908  &  n_n53 ) ;
 assign wire22286 = ( wire479 ) | ( wire656 ) | ( wire2507 ) ;
 assign wire22287 = ( wire629 ) | ( wire462 ) | ( wire2508 ) | ( wire22282 ) ;
 assign n_n1137 = ( n_n1255 ) | ( wire22286 ) | ( wire22287 ) ;
 assign wire2879 = ( wire95  &  n_n3 ) | ( n_n3  &  wire21913 ) ;
 assign wire21914 = ( n_n4  &  n_n8 ) | ( n_n4  &  n_n61 ) | ( n_n4  &  n_n62 ) ;
 assign n_n1157 = ( wire2879 ) | ( wire21914 ) | ( wire169  &  n_n10 ) ;
 assign wire1112 = ( wire75 ) | ( wire63 ) | ( n_n58 ) | ( wire223 ) ;
 assign n_n1295 = ( wire747 ) | ( wire22187 ) | ( wire22188 ) ;
 assign n_n1641 = ( n_n100  &  wire69 ) | ( n_n94  &  n_n103 ) ;
 assign wire22190 = ( n_n94  &  n_n38 ) | ( n_n94  &  n_n86 ) | ( n_n94  &  wire1334 ) ;
 assign wire22193 = ( n_n1645 ) | ( wire773 ) | ( wire49  &  n_n100 ) ;
 assign n_n1151 = ( n_n1295 ) | ( n_n1641 ) | ( wire22190 ) | ( wire22193 ) ;
 assign wire1113 = ( (~ i_14_)  &  i_13_  &  i_12_  &  wire902 ) | ( i_14_  &  (~ i_13_)  &  i_12_  &  wire902 ) | ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire902 ) | ( i_14_  &  i_13_  &  (~ i_12_)  &  wire902 ) | ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  wire902 ) ;
 assign wire22185 = ( n_n1624 ) | ( wire22181 ) | ( n_n100  &  wire1044 ) ;
 assign n_n1102 = ( n_n1151 ) | ( wire2602 ) | ( _39743 ) | ( _39744 ) ;
 assign n_n1284 = ( n_n4687 ) | ( wire22213 ) | ( wire22214 ) ;
 assign wire22219 = ( wire484 ) | ( wire2581 ) | ( wire22217 ) ;
 assign wire22220 = ( wire2583 ) | ( _1394 ) ;
 assign wire807 = ( (~ i_14_)  &  i_13_  &  i_12_  &  wire898 ) | ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire898 ) ;
 assign n_n4675 = ( n_n56  &  wire807 ) | ( n_n279  &  n_n56  &  wire904 ) ;
 assign n_n4681 = ( n_n56  &  n_n42 ) | ( n_n57  &  wire81 ) ;
 assign n_n1604 = ( n_n54  &  n_n56 ) | ( n_n57  &  wire51 ) ;
 assign wire497 = ( n_n220  &  n_n56  &  wire904 ) | ( n_n56  &  n_n256  &  wire904 ) ;
 assign wire22227 = ( n_n4960 ) | ( n_n4675 ) | ( n_n4681 ) | ( n_n1604 ) ;
 assign wire22228 = ( n_n4961 ) | ( wire497 ) | ( wire2571 ) | ( wire2572 ) ;
 assign n_n1101 = ( _39785 ) | ( _39786 ) ;
 assign n_n1298 = ( wire2566 ) | ( wire22231 ) | ( wire22232 ) ;
 assign wire22236 = ( n_n100  &  _39793 ) | ( wire907  &  n_n100  &  _36783 ) ;
 assign n_n1152 = ( n_n1298 ) | ( wire2560 ) | ( wire2561 ) | ( _39796 ) ;
 assign wire874 = ( wire22240 ) | ( wire22241 ) | ( wire22242 ) ;
 assign n_n1154 = ( wire874 ) | ( wire20755 ) | ( _1372 ) | ( _39805 ) ;
 assign n_n3881 = ( wire51  &  n_n100 ) | ( n_n54  &  n_n94 ) ;
 assign wire784 = ( wire166  &  n_n100 ) | ( wire180  &  n_n100 ) ;
 assign n_n1103 = ( n_n1152 ) | ( n_n1154 ) | ( wire2545 ) | ( _39811 ) ;
 assign wire647 = ( n_n6  &  n_n216 ) | ( n_n6  &  n_n203 ) | ( n_n6  &  wire20149 ) ;
 assign wire22785 = ( n_n228  &  wire902  &  n_n53 ) | ( n_n228  &  wire899  &  n_n53 ) ;
 assign wire356 = ( (~ i_14_)  &  i_15_  &  n_n253  &  n_n254 ) | ( i_14_  &  (~ i_15_)  &  n_n253  &  n_n254 ) | ( (~ i_14_)  &  (~ i_15_)  &  n_n253  &  n_n254 ) ;
 assign wire22613 = ( n_n206  &  n_n100 ) | ( n_n206  &  n_n94 ) | ( n_n226  &  n_n94 ) ;
 assign n_n850 = ( n_n4970 ) | ( wire22613 ) | ( n_n57  &  wire356 ) ;
 assign wire335 = ( (~ i_14_)  &  i_15_  &  n_n254  &  n_n267 ) | ( i_14_  &  (~ i_15_)  &  n_n254  &  n_n267 ) | ( (~ i_14_)  &  (~ i_15_)  &  n_n254  &  n_n267 ) ;
 assign wire1121 = ( n_n228  &  wire912 ) | ( n_n228  &  wire902 ) | ( n_n228  &  wire897 ) ;
 assign wire1120 = ( n_n228  &  wire912 ) | ( n_n228  &  wire902 ) | ( n_n228  &  wire897 ) ;
 assign wire2138 = ( n_n285  &  n_n271  &  n_n230  &  wire335 ) ;
 assign wire22616 = ( n_n226  &  n_n100 ) | ( n_n100  &  n_n63 ) | ( n_n94  &  n_n63 ) ;
 assign n_n4628 = ( n_n6  &  wire19457 ) | ( n_n6  &  n_n222  &  wire897 ) ;
 assign wire727 = ( n_n5  &  wire88 ) | ( n_n5  &  n_n31 ) | ( n_n5  &  n_n80 ) ;
 assign n_n431 = ( wire22403 ) | ( wire22404 ) | ( _40169 ) ;
 assign wire22409 = ( n_n53  &  n_n10 ) | ( n_n48  &  n_n13 ) | ( n_n53  &  n_n13 ) ;
 assign wire22412 = ( n_n4153 ) | ( n_n618 ) | ( wire2378 ) ;
 assign wire2374 = ( n_n48  &  wire57 ) | ( wire914  &  n_n279  &  n_n48 ) ;
 assign wire22414 = ( wire914  &  n_n256  &  n_n48 ) | ( wire912  &  n_n256  &  n_n48 ) ;
 assign wire22415 = ( n_n6  &  n_n54 ) | ( n_n53  &  n_n10 ) ;
 assign wire22416 = ( n_n246  &  n_n48 ) | ( n_n6  &  n_n98 ) ;
 assign n_n429 = ( wire2374 ) | ( wire22414 ) | ( wire22415 ) | ( wire22416 ) ;
 assign wire22400 = ( wire2392 ) | ( wire22399 ) ;
 assign wire22401 = ( wire624 ) | ( wire2393 ) | ( wire2398 ) | ( wire22395 ) ;
 assign n_n343 = ( _40200 ) | ( _40201 ) ;
 assign wire2361 = ( n_n5  &  wire320 ) | ( wire914  &  n_n5  &  n_n256 ) ;
 assign wire2356 = ( _830 ) | ( n_n6  &  n_n109 ) | ( n_n6  &  wire143 ) ;
 assign wire2353 = ( n_n5  &  wire245 ) | ( n_n5  &  n_n40 ) | ( n_n5  &  wire351 ) ;
 assign wire2354 = ( n_n6  &  n_n34 ) | ( n_n6  &  n_n81 ) | ( n_n6  &  wire47 ) ;
 assign n_n363 = ( wire2354 ) | ( _817 ) | ( _40252 ) | ( _40262 ) ;
 assign n_n438 = ( n_n6848 ) | ( wire2374 ) | ( wire22414 ) | ( n_n618 ) ;
 assign wire22446 = ( n_n48  &  n_n103 ) | ( n_n53  &  n_n103 ) | ( n_n53  &  wire140 ) ;
 assign n_n443 = ( n_n4183 ) | ( wire22451 ) | ( wire41  &  n_n53 ) ;
 assign wire22454 = ( n_n105  &  n_n48 ) | ( n_n105  &  n_n53 ) | ( n_n53  &  wire175 ) ;
 assign wire22457 = ( wire22456 ) | ( n_n57  &  wire1678 ) ;
 assign wire809 = ( n_n258  &  wire898  &  n_n48 ) ;
 assign wire22459 = ( i_15_  &  n_n256  &  n_n247 ) | ( (~ i_15_)  &  n_n256  &  n_n247 ) | ( i_15_  &  n_n256  &  n_n267 ) | ( (~ i_15_)  &  n_n256  &  n_n267 ) ;
 assign wire1128 = ( wire166 ) | ( wire57 ) | ( n_n113 ) | ( wire22459 ) ;
 assign wire22463 = ( wire2311 ) | ( wire22461 ) | ( n_n54  &  n_n48 ) ;
 assign wire22464 = ( wire2333 ) | ( wire22449 ) | ( n_n53  &  wire1128 ) ;
 assign n_n143 = ( i_9_  &  i_10_  &  i_12_  &  (~ i_11_) ) ;
 assign n_n39 = ( (~ i_14_)  &  i_13_  &  i_12_  &  wire912 ) ;
 assign n_n77 = ( (~ i_14_)  &  i_13_  &  i_12_  &  wire908 ) ;
 assign n_n67 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire913 ) ;
 assign wire1131 = ( (~ i_13_) ) | ( (~ i_12_) ) | ( (~ i_14_)  &  i_13_  &  i_12_ ) ;
 assign wire19213 = ( wire19212 ) | ( n_n228  &  wire903 ) ;
 assign wire1130 = ( wire19213 ) | ( n_n275  &  wire1131 ) ;
 assign wire5893 = ( (~ i_14_)  &  i_13_  &  i_12_  &  _34780 ) | ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  _34780 ) | ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  _34780 ) ;
 assign wire19215 = ( i_9_  &  i_10_  &  i_11_ ) | ( i_9_  &  (~ i_10_)  &  i_11_  &  n_n256 ) ;
 assign wire19216 = ( i_14_  &  i_13_  &  (~ i_12_)  &  wire899 ) | ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire899 ) ;
 assign wire19217 = ( n_n258  &  wire908 ) | ( n_n228  &  wire899 ) ;
 assign wire1132 = ( wire5893 ) | ( wire19215 ) | ( wire19216 ) | ( wire19217 ) ;
 assign wire190 = ( i_14_  &  (~ i_13_)  &  i_12_  &  wire897 ) | ( i_14_  &  i_13_  &  (~ i_12_)  &  wire897 ) | ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire897 ) ;
 assign n_n4941 = ( n_n56  &  wire57 ) | ( wire914  &  n_n279  &  n_n56 ) ;
 assign n_n4942 = ( n_n56  &  wire55 ) | ( n_n279  &  wire912  &  n_n56 ) ;
 assign wire157 = ( (~ i_14_)  &  i_13_  &  i_12_  &  wire914 ) | ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire914 ) | ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  wire914 ) ;
 assign wire728 = ( wire273  &  n_n56 ) | ( n_n56  &  wire157 ) ;
 assign wire729 = ( wire112  &  n_n57 ) | ( n_n57  &  wire277 ) ;
 assign n_n5685 = ( (~ i_7_)  &  i_6_  &  n_n260  &  n_n116 ) ;
 assign wire4889 = ( wire48  &  n_n128 ) | ( wire913  &  n_n220  &  n_n128 ) ;
 assign wire20020 = ( wire4892 ) | ( wire913  &  n_n220  &  n_n130 ) ;
 assign wire20021 = ( n_n5693 ) | ( wire452 ) | ( wire758 ) | ( wire4890 ) ;
 assign wire4882 = ( n_n264  &  n_n118  &  n_n231 ) | ( n_n118  &  n_n231  &  n_n230 ) ;
 assign wire20023 = ( n_n264  &  n_n118  &  n_n155 ) | ( n_n284  &  n_n118  &  n_n155 ) ;
 assign wire20027 = ( n_n5659 ) | ( n_n5673 ) | ( n_n5664 ) | ( wire587 ) ;
 assign wire794 = ( (~ i_7_)  &  i_6_  &  n_n116  &  n_n230 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n116  &  n_n230 ) ;
 assign n_n4394 = ( n_n285  &  n_n266  &  n_n230  &  wire247 ) ;
 assign n_n4381 = ( n_n57  &  wire63 ) | ( n_n281  &  n_n57  &  wire908 ) ;
 assign n_n3850 = ( n_n9  &  n_n56 ) | ( n_n57  &  wire132 ) ;
 assign wire5587 = ( n_n56  &  n_n7 ) | ( n_n56  &  wire50 ) | ( n_n56  &  n_n59 ) ;
 assign wire473 = ( wire5587 ) | ( n_n57  &  wire137 ) ;
 assign wire124 = ( i_14_  &  i_13_  &  i_12_  &  wire903 ) | ( i_14_  &  i_13_  &  (~ i_12_)  &  wire903 ) | ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire903 ) ;
 assign n_n4929 = ( n_n285  &  n_n266  &  n_n230  &  wire124 ) ;
 assign wire212 = ( (~ i_14_)  &  i_13_  &  i_12_  &  wire897 ) | ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire897 ) | ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  wire897 ) ;
 assign wire250 = ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  wire905 ) | ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire905 ) ;
 assign wire1141 = ( n_n229  &  n_n165  &  n_n284 ) | ( n_n165  &  n_n284  &  n_n283 ) ;
 assign wire4166 = ( n_n152  &  wire103 ) | ( n_n152  &  n_n220  &  wire905 ) ;
 assign wire20712 = ( n_n5796 ) | ( n_n139  &  n_n281  &  wire899 ) ;
 assign n_n4279 = ( n_n4970 ) | ( wire4166 ) | ( wire20712 ) ;
 assign wire4569 = ( n_n48  &  n_n7 ) | ( n_n48  &  wire50 ) | ( n_n48  &  n_n59 ) ;
 assign wire4570 = ( n_n53  &  wire50 ) | ( n_n228  &  n_n53  &  wire897 ) ;
 assign wire20273 = ( n_n53  &  _37155 ) | ( wire902  &  n_n53  &  _35049 ) ;
 assign n_n3978 = ( wire4569 ) | ( wire4570 ) | ( wire20273 ) ;
 assign n_n1346 = ( n_n3  &  n_n41 ) | ( n_n4  &  wire78 ) ;
 assign n_n884 = ( n_n4  &  wire88 ) | ( n_n4  &  wire902  &  n_n222 ) ;
 assign wire21228 = ( n_n1341 ) | ( n_n1346 ) | ( wire21225 ) ;
 assign n_n3908 = ( wire21228 ) | ( _3235 ) | ( _3236 ) | ( _38254 ) ;
 assign n_n3778 = ( n_n2  &  wire68 ) | ( n_n1  &  n_n42 ) ;
 assign n_n3229 = ( n_n3  &  n_n108 ) | ( n_n4  &  wire70 ) ;
 assign wire740 = ( wire44  &  n_n100 ) | ( n_n258  &  wire904  &  n_n100 ) ;
 assign n_n1555 = ( n_n95  &  n_n48 ) | ( n_n53  &  wire55 ) ;
 assign wire626 = ( n_n53  &  _37263 ) | ( wire908  &  n_n53  &  _35046 ) ;
 assign n_n3791 = ( n_n60  &  n_n53 ) | ( n_n8  &  n_n53 ) | ( n_n61  &  n_n53 ) ;
 assign wire478 = ( n_n53  &  _35118 ) | ( wire908  &  n_n53  &  _35120 ) ;
 assign wire20387 = ( n_n53  &  _37469 ) | ( wire902  &  n_n53  &  _35622 ) ;
 assign wire736 = ( n_n4073 ) | ( wire479 ) | ( wire478 ) | ( wire20387 ) ;
 assign wire20392 = ( n_n4068 ) | ( n_n4069 ) | ( wire20390 ) ;
 assign n_n2815 = ( n_n3964 ) | ( wire736 ) | ( wire20392 ) ;
 assign n_n2982 = ( n_n60  &  n_n4 ) | ( n_n4  &  n_n8 ) | ( n_n4  &  n_n226 ) ;
 assign wire349 = ( n_n228  &  n_n3  &  wire898 ) ;
 assign wire483 = ( wire88  &  n_n53 ) | ( n_n53  &  n_n31 ) | ( n_n53  &  n_n80 ) ;
 assign wire876 = ( n_n4076 ) | ( wire483 ) | ( n_n4  &  n_n257 ) ;
 assign wire20996 = ( wire876 ) | ( wire20993 ) | ( wire20994 ) ;
 assign n_n3097 = ( n_n3116 ) | ( n_n2815 ) | ( wire20996 ) ;
 assign n_n3099 = ( n_n3122 ) | ( wire21019 ) | ( _37976 ) | ( _37989 ) ;
 assign n_n3101 = ( n_n3128 ) | ( wire21054 ) | ( _37993 ) | ( _37994 ) ;
 assign wire21063 = ( n_n3124 ) | ( n_n3123 ) | ( wire21061 ) ;
 assign n_n3103 = ( n_n3132 ) | ( n_n3133 ) | ( wire21093 ) | ( _38057 ) ;
 assign wire21122 = ( wire21070 ) | ( n_n3130 ) | ( wire21120 ) | ( _38087 ) ;
 assign wire4694 = ( n_n5  &  wire79 ) | ( n_n5  &  n_n20 ) | ( n_n5  &  wire83 ) ;
 assign wire4695 = ( n_n6  &  wire44 ) | ( n_n6  &  n_n252 ) | ( n_n6  &  n_n15 ) ;
 assign n_n3864 = ( wire63  &  n_n100 ) | ( n_n228  &  wire902  &  n_n100 ) ;
 assign wire780 = ( n_n281  &  wire908  &  n_n100 ) ;
 assign n_n2702 = ( n_n106  &  n_n100 ) | ( wire160  &  n_n94 ) ;
 assign wire654 = ( n_n94  &  _36825 ) | ( wire914  &  n_n94  &  _34565 ) ;
 assign wire1372 = ( (~ i_14_)  &  i_13_  &  i_12_  &  wire913 ) | ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire913 ) ;
 assign n_n2398 = ( n_n94  &  wire1372 ) | ( wire913  &  n_n220  &  n_n94 ) ;
 assign wire1150 = ( wire60 ) | ( n_n204 ) | ( wire247 ) | ( wire210 ) ;
 assign n_n2724 = ( wire160  &  n_n100 ) | ( n_n66  &  n_n94 ) ;
 assign wire1156 = ( n_n270  &  _38788 ) | ( n_n270  &  _38789 ) ;
 assign wire3340 = ( n_n207  &  wire21536 ) | ( n_n225  &  wire903  &  n_n207 ) ;
 assign wire21537 = ( n_n5  &  n_n145 ) | ( n_n207  &  n_n67 ) ;
 assign wire21538 = ( n_n151  &  wire164 ) | ( n_n227  &  wire1156 ) ;
 assign n_n2133 = ( wire3340 ) | ( wire21537 ) | ( wire21538 ) ;
 assign wire388 = ( n_n94  &  _37878 ) | ( wire913  &  n_n94  &  _36810 ) ;
 assign wire747 = ( wire40  &  n_n94 ) | ( n_n281  &  n_n94  &  wire897 ) ;
 assign wire21540 = ( n_n70  &  n_n227 ) | ( n_n94  &  n_n200 ) ;
 assign wire21541 = ( n_n204  &  n_n94 ) | ( n_n227  &  n_n109 ) ;
 assign n_n2132 = ( wire388 ) | ( wire747 ) | ( wire21540 ) | ( wire21541 ) ;
 assign wire391 = ( wire907  &  n_n225  &  n_n100 ) | ( wire907  &  n_n256  &  n_n100 ) ;
 assign wire21549 = ( wire3324 ) | ( wire21544 ) | ( wire21545 ) | ( wire21546 ) ;
 assign wire330 = ( i_15_  &  n_n281  &  n_n247 ) | ( i_15_  &  n_n279  &  n_n247 ) | ( (~ i_15_)  &  n_n279  &  n_n247 ) ;
 assign wire241 = ( i_15_  &  n_n281  &  n_n267 ) | ( i_15_  &  n_n279  &  n_n267 ) | ( (~ i_15_)  &  n_n279  &  n_n267 ) ;
 assign wire1159 = ( wire153 ) | ( wire157 ) | ( wire330 ) | ( wire241 ) ;
 assign wire21425 = ( n_n4  &  n_n108 ) | ( n_n4  &  n_n70 ) | ( n_n4  &  n_n93 ) ;
 assign n_n2129 = ( wire3518 ) | ( wire21425 ) | ( n_n3  &  n_n186 ) ;
 assign wire21431 = ( wire476 ) | ( wire21426 ) | ( wire21428 ) ;
 assign wire21432 = ( wire3480 ) | ( wire21427 ) | ( _2633 ) ;
 assign n_n2274 = ( n_n53  &  n_n76 ) | ( n_n53  &  n_n26 ) | ( n_n53  &  n_n77 ) ;
 assign wire1163 = ( i_15_  &  n_n279  &  n_n270 ) | ( (~ i_15_)  &  n_n279  &  n_n270 ) | ( i_15_  &  n_n279  &  n_n259 ) | ( (~ i_15_)  &  n_n279  &  n_n259 ) ;
 assign wire2780 = ( n_n5  &  wire223 ) | ( n_n220  &  wire911  &  n_n5 ) ;
 assign wire2781 = ( n_n207  &  wire425 ) | ( n_n228  &  wire903  &  n_n207 ) ;
 assign wire22022 = ( n_n6  &  wire75 ) | ( n_n103  &  n_n207 ) ;
 assign n_n1217 = ( wire2780 ) | ( wire2781 ) | ( wire22022 ) ;
 assign n_n4687 = ( n_n57  &  wire807 ) | ( n_n279  &  n_n57  &  wire904 ) ;
 assign wire22213 = ( n_n258  &  n_n57  &  wire898 ) | ( n_n57  &  wire898  &  n_n222 ) ;
 assign wire22214 = ( n_n94  &  wire223 ) | ( n_n57  &  wire486 ) ;
 assign wire2503 = ( _1686 ) | ( n_n48  &  wire433 ) | ( n_n48  &  wire22290 ) ;
 assign wire750 = ( n_n2  &  wire200 ) | ( n_n2  &  wire112 ) ;
 assign n_n1433 = ( wire66  &  n_n53 ) | ( wire899  &  n_n256  &  n_n53 ) ;
 assign wire1171 = ( i_14_  &  (~ i_13_)  &  i_12_  &  wire907 ) | ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire907 ) | ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  wire907 ) ;
 assign wire22034 = ( n_n257  &  n_n53 ) | ( n_n2  &  wire85 ) ;
 assign wire22040 = ( wire456 ) | ( wire626 ) | ( _39817 ) ;
 assign wire22041 = ( n_n1433 ) | ( wire22035 ) | ( wire22039 ) ;
 assign n_n1120 = ( wire750 ) | ( wire22034 ) | ( wire22040 ) | ( wire22041 ) ;
 assign n_n1476 = ( n_n5  &  n_n197 ) | ( n_n6  &  wire62 ) ;
 assign wire2777 = ( _1248 ) | ( n_n6  &  wire247 ) | ( n_n6  &  wire220 ) ;
 assign wire589 = ( n_n56  &  n_n197 ) | ( n_n57  &  wire62 ) ;
 assign wire2525 = ( n_n57  &  n_n107 ) | ( n_n57  &  n_n112 ) | ( n_n57  &  wire52 ) ;
 assign wire22270 = ( n_n4921 ) | ( n_n4394 ) | ( wire481 ) | ( n_n4915 ) ;
 assign wire2521 = ( n_n56  &  wire22275 ) | ( n_n56  &  wire22276 ) ;
 assign wire22277 = ( wire2520 ) | ( wire2532 ) | ( wire2533 ) ;
 assign n_n3843 = ( n_n95  &  n_n53 ) | ( n_n48  &  wire81 ) ;
 assign wire19385 = ( n_n267  &  _35164 ) | ( n_n267  &  _35165 ) ;
 assign wire662 = ( n_n53  &  wire19385 ) | ( n_n256  &  wire900  &  n_n53 ) ;
 assign n_n1584 = ( n_n57  &  n_n197 ) | ( n_n56  &  wire69 ) ;
 assign wire706 = ( n_n285  &  n_n271  &  n_n230  &  wire165 ) ;
 assign wire406 = ( n_n258  &  wire899  &  n_n53 ) | ( n_n222  &  wire899  &  n_n53 ) ;
 assign n_n952 = ( n_n53  &  n_n197 ) | ( n_n53  &  n_n223 ) | ( n_n53  &  n_n221 ) ;
 assign wire1984 = ( n_n6  &  n_n37 ) | ( n_n6  &  wire126 ) | ( n_n6  &  wire89 ) ;
 assign wire22736 = ( n_n6  &  n_n104 ) | ( n_n5  &  n_n41 ) ;
 assign n_n819 = ( wire1984 ) | ( wire22736 ) | ( n_n5  &  wire126 ) ;
 assign wire930 = ( (~ i_1_)  &  (~ i_2_)  &  i_0_  &  _37619 ) ;
 assign n_n5673 = ( (~ i_7_)  &  i_6_  &  n_n264  &  n_n116 ) ;
 assign n_n59 = ( i_14_  &  i_13_  &  i_12_  &  wire897 ) ;
 assign n_n90 = ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  wire900 ) ;
 assign wire6020 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  _34919 ) | ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  _34919 ) ;
 assign wire19269 = ( n_n267 ) | ( n_n258  &  wire903 ) ;
 assign wire19270 = ( i_14_  &  i_13_  &  (~ i_12_)  &  wire903 ) | ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire903 ) ;
 assign wire19271 = ( n_n242  &  wire1182 ) | ( i_15_  &  n_n242  &  n_n222 ) ;
 assign wire1181 = ( wire6020 ) | ( wire19269 ) | ( wire19270 ) | ( wire19271 ) ;
 assign wire1187 = ( i_9_ ) | ( (~ i_9_)  &  i_10_ ) | ( (~ i_9_)  &  (~ i_10_)  &  i_11_ ) ;
 assign wire1186 = ( i_9_  &  i_10_ ) | ( (~ i_9_)  &  i_10_  &  i_11_ ) | ( i_9_  &  (~ i_10_)  &  i_11_ ) | ( (~ i_9_)  &  (~ i_10_)  &  (~ i_11_) ) ;
 assign wire5885 = ( n_n227  &  wire65 ) | ( n_n227  &  wire19220 ) | ( n_n227  &  wire19221 ) ;
 assign wire19223 = ( wire5900 ) | ( n_n227  &  wire1130 ) | ( n_n227  &  wire1132 ) ;
 assign wire19230 = ( n_n5063 ) | ( wire19228 ) | ( _6708 ) ;
 assign n_n5007 = ( n_n5020 ) | ( wire5885 ) | ( wire19223 ) | ( wire19230 ) ;
 assign wire936 = ( (~ i_1_)  &  (~ i_2_)  &  i_0_  &  _36585 ) ;
 assign wire198 = ( i_14_  &  (~ i_13_)  &  i_12_  &  wire902 ) | ( i_14_  &  i_13_  &  (~ i_12_)  &  wire902 ) | ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire902 ) ;
 assign wire760 = ( n_n57  &  wire167 ) | ( n_n56  &  wire190 ) ;
 assign wire119 = ( (~ i_14_)  &  i_13_  &  i_12_  &  wire903 ) | ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire903 ) | ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  wire903 ) ;
 assign wire761 = ( n_n57  &  wire190 ) | ( n_n56  &  wire119 ) ;
 assign wire762 = ( n_n57  &  wire140 ) | ( n_n57  &  wire165 ) ;
 assign wire5076 = ( n_n6  &  wire95 ) | ( n_n281  &  wire914  &  n_n6 ) ;
 assign wire19878 = ( n_n4826 ) | ( n_n4823 ) | ( wire584 ) | ( n_n4821 ) ;
 assign wire763 = ( n_n285  &  n_n266  &  n_n230  &  wire119 ) ;
 assign n_n4183 = ( wire579 ) | ( wire764 ) | ( n_n54  &  n_n53 ) ;
 assign n_n4770 = ( n_n5  &  wire99 ) | ( n_n5  &  wire41 ) | ( n_n5  &  wire254 ) ;
 assign n_n4160 = ( wire95  &  n_n53 ) | ( n_n228  &  wire912  &  n_n53 ) ;
 assign wire1279 = ( n_n247  &  _38062 ) | ( n_n247  &  _38063 ) ;
 assign n_n1645 = ( n_n94  &  wire1279 ) | ( wire912  &  n_n225  &  n_n94 ) ;
 assign wire767 = ( n_n100  &  n_n41 ) | ( n_n100  &  wire368 ) | ( n_n100  &  n_n88 ) ;
 assign wire21098 = ( n_n94  &  n_n41 ) | ( n_n94  &  wire77 ) | ( n_n94  &  n_n86 ) ;
 assign wire21101 = ( n_n1066 ) | ( n_n1645 ) | ( wire3778 ) ;
 assign n_n3309 = ( n_n108  &  n_n48 ) | ( wire70  &  n_n53 ) ;
 assign wire463 = ( n_n48  &  _37977 ) | ( wire914  &  n_n48  &  _37163 ) ;
 assign wire20999 = ( n_n108  &  n_n53 ) | ( n_n48  &  wire82 ) ;
 assign wire21003 = ( wire463 ) | ( _3503 ) | ( wire44  &  _38018 ) ;
 assign wire21004 = ( n_n4160 ) | ( wire20998 ) | ( _3498 ) ;
 assign n_n3124 = ( n_n3309 ) | ( wire20999 ) | ( wire21003 ) | ( wire21004 ) ;
 assign wire3852 = ( n_n48  &  n_n179 ) | ( n_n48  &  wire57 ) | ( n_n48  &  wire21009 ) ;
 assign wire681 = ( wire3852 ) | ( wire912  &  n_n256  &  n_n48 ) ;
 assign wire21013 = ( n_n3791 ) | ( n_n48  &  n_n147 ) | ( n_n48  &  n_n148 ) ;
 assign wire21014 = ( wire461 ) | ( wire3843 ) | ( wire21010 ) ;
 assign n_n3123 = ( n_n3184 ) | ( wire681 ) | ( wire21013 ) | ( wire21014 ) ;
 assign n_n3122 = ( wire21027 ) | ( wire21028 ) | ( _4342 ) | ( _37285 ) ;
 assign wire21035 = ( wire727 ) | ( n_n4632 ) | ( wire487 ) | ( wire21030 ) ;
 assign n_n3128 = ( n_n3324 ) | ( n_n4381 ) | ( wire21046 ) | ( wire21047 ) ;
 assign wire21054 = ( wire3852 ) | ( wire21051 ) | ( _3512 ) | ( _38014 ) ;
 assign n_n3587 = ( n_n53  &  wire42 ) | ( n_n279  &  wire899  &  n_n53 ) ;
 assign wire770 = ( n_n48  &  n_n76 ) | ( n_n48  &  n_n26 ) | ( n_n48  &  wire80 ) ;
 assign wire771 = ( wire88  &  n_n48 ) | ( n_n48  &  n_n29 ) | ( n_n48  &  wire49 ) ;
 assign n_n3132 = ( wire370 ) | ( wire788 ) | ( wire21077 ) | ( wire21081 ) ;
 assign n_n3133 = ( n_n3209 ) | ( wire21089 ) | ( wire21090 ) ;
 assign wire21116 = ( n_n3221 ) | ( wire21114 ) | ( _5922 ) | ( _35714 ) ;
 assign wire653 = ( _4177 ) | ( n_n57  &  wire453 ) | ( n_n57  &  n_n38 ) ;
 assign wire548 = ( n_n94  &  _36682 ) | ( n_n247  &  n_n94  &  _36683 ) ;
 assign wire773 = ( n_n100  &  wire140 ) | ( n_n100  &  wire165 ) ;
 assign wire774 = ( n_n220  &  wire907  &  n_n100 ) ;
 assign wire20056 = ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire912 ) | ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  wire912 ) ;
 assign wire1194 = ( wire57 ) | ( n_n113 ) | ( wire157 ) | ( wire20056 ) ;
 assign wire20060 = ( wire686 ) | ( wire391 ) | ( wire548 ) | ( wire774 ) ;
 assign n_n2665 = ( wire773 ) | ( wire20060 ) | ( _4977 ) | ( _36687 ) ;
 assign wire1196 = ( i_8_  &  n_n260  &  n_n272  &  n_n285 ) | ( (~ i_8_)  &  n_n260  &  n_n272  &  n_n285 ) ;
 assign wire1195 = ( n_n220  &  wire911 ) | ( n_n220  &  wire897 ) ;
 assign wire1198 = ( n_n220  &  wire912 ) | ( n_n220  &  wire898 ) | ( n_n220  &  wire900 ) ;
 assign wire3005 = ( n_n6  &  wire230 ) | ( n_n6  &  n_n222  &  wire897 ) ;
 assign wire3198 = ( n_n268  &  n_n58 ) | ( n_n268  &  wire429 ) | ( n_n268  &  wire21658 ) ;
 assign wire21660 = ( n_n268  &  wire273 ) | ( n_n265  &  n_n32 ) ;
 assign wire21665 = ( wire21662 ) | ( wire21663 ) | ( n_n268  &  wire247 ) ;
 assign n_n1697 = ( wire21665 ) | ( wire3190 ) | ( _2412 ) | ( _38945 ) ;
 assign wire690 = ( n_n3  &  _38969 ) | ( n_n3  &  wire898  &  _38971 ) ;
 assign wire270 = ( n_n267  &  _38965 ) | ( n_n267  &  _38966 ) ;
 assign wire3186 = ( n_n3  &  n_n99 ) | ( n_n3  &  n_n52 ) | ( n_n3  &  wire807 ) ;
 assign wire21657 = ( wire3203 ) | ( wire3211 ) | ( wire21651 ) | ( wire21655 ) ;
 assign wire21673 = ( wire3186 ) | ( wire3187 ) | ( wire21670 ) | ( wire21671 ) ;
 assign n_n1753 = ( wire21675 ) | ( wire21676 ) | ( wire21677 ) | ( wire21678 ) ;
 assign wire3159 = ( wire143  &  _39051 ) | ( wire21668  &  _39051 ) | ( _39048  &  _39051 ) ;
 assign wire21683 = ( wire690 ) | ( wire622 ) | ( wire21681 ) ;
 assign n_n1703 = ( n_n1753 ) | ( wire21683 ) | ( _39055 ) ;
 assign wire21697 = ( wire657 ) | ( wire21694 ) | ( wire21695 ) ;
 assign n_n1704 = ( n_n1757 ) | ( n_n1756 ) | ( wire21697 ) ;
 assign wire21699 = ( n_n281  &  wire899  &  n_n53 ) | ( wire899  &  n_n256  &  n_n53 ) ;
 assign wire21700 = ( n_n53  &  _39081 ) | ( wire902  &  n_n53  &  _35049 ) ;
 assign wire21701 = ( n_n220  &  wire905  &  n_n53 ) | ( n_n220  &  wire899  &  n_n53 ) ;
 assign wire21702 = ( n_n2  &  n_n37 ) | ( n_n53  &  wire1849 ) ;
 assign n_n1752 = ( wire21699 ) | ( wire21700 ) | ( wire21701 ) | ( wire21702 ) ;
 assign wire21648 = ( _39009 ) | ( n_n1  &  wire21647 ) ;
 assign wire21649 = ( wire3219 ) | ( wire3220 ) | ( wire3221 ) | ( wire3222 ) ;
 assign n_n1356 = ( n_n229  &  n_n284  &  n_n285  &  wire99 ) ;
 assign wire22043 = ( n_n4  &  n_n258  &  wire906 ) | ( n_n4  &  n_n258  &  wire908 ) ;
 assign wire22044 = ( n_n220  &  n_n4  &  wire902 ) | ( n_n220  &  n_n4  &  wire899 ) ;
 assign n_n1208 = ( wire476 ) | ( n_n1356 ) | ( wire22043 ) | ( wire22044 ) ;
 assign n_n639 = ( n_n264  &  n_n273  &  n_n285  &  wire140 ) ;
 assign wire694 = ( n_n53  &  wire61 ) | ( n_n281  &  wire902  &  n_n53 ) ;
 assign wire869 = ( wire902  &  n_n258  &  n_n53 ) | ( wire902  &  n_n222  &  n_n53 ) ;
 assign wire22053 = ( wire409 ) | ( wire479 ) | ( wire22050 ) ;
 assign wire22054 = ( wire22047 ) | ( wire22048 ) | ( wire22052 ) ;
 assign n_n1121 = ( n_n1208 ) | ( wire22053 ) | ( wire22054 ) ;
 assign n_n876 = ( n_n4  &  wire469 ) | ( n_n4  &  n_n222  &  wire899 ) ;
 assign wire850 = ( n_n268  &  wire20362 ) | ( n_n279  &  n_n268  &  wire897 ) ;
 assign wire22775 = ( n_n228  &  n_n1  &  wire899 ) | ( n_n228  &  n_n2  &  wire899 ) ;
 assign wire22776 = ( n_n268  &  wire56 ) | ( n_n206  &  wire135 ) ;
 assign n_n790 = ( wire850 ) | ( wire22775 ) | ( wire22776 ) ;
 assign wire743 = ( n_n4  &  _40205 ) | ( wire905  &  n_n4  &  _39673 ) ;
 assign wire232 = ( (~ i_15_)  &  n_n228  &  n_n242 ) | ( i_15_  &  n_n242  &  n_n258 ) ;
 assign wire22336 = ( wire913  &  n_n256 ) | ( wire908  &  n_n256 ) ;
 assign wire1213 = ( n_n17 ) | ( wire514 ) | ( wire232 ) | ( wire22336 ) ;
 assign wire22338 = ( wire2472 ) | ( wire2473 ) | ( wire22337 ) ;
 assign wire2463 = ( n_n3  &  n_n52 ) | ( n_n3  &  wire357 ) | ( n_n3  &  wire22340 ) ;
 assign wire22348 = ( wire2463 ) | ( wire22346 ) | ( _40414 ) ;
 assign wire22351 = ( n_n4  &  wire320 ) | ( n_n4  &  wire908  &  n_n256 ) ;
 assign wire642 = ( n_n4  &  _40208 ) | ( n_n4  &  wire908  &  _39470 ) ;
 assign wire351 = ( n_n247  &  _40253 ) | ( n_n247  &  _40254 ) ;
 assign wire22352 = ( wire914  &  n_n256 ) | ( wire907  &  n_n256 ) ;
 assign wire1217 = ( wire245 ) | ( n_n40 ) | ( wire351 ) | ( wire22352 ) ;
 assign wire19341 = ( wire5861 ) | ( wire19331 ) | ( wire19339 ) ;
 assign wire19284 = ( i_11_  &  n_n281  &  n_n163 ) | ( (~ i_11_)  &  n_n281  &  n_n163 ) | ( i_11_  &  n_n163  &  n_n278 ) | ( (~ i_11_)  &  n_n163  &  n_n278 ) ;
 assign wire19285 = ( wire5999 ) | ( n_n279  &  wire901 ) | ( n_n279  &  wire897 ) ;
 assign n_n5051 = ( n_n177  &  wire19284 ) | ( n_n177  &  wire19285 ) ;
 assign wire1223 = ( (~ i_9_) ) | ( i_9_  &  (~ i_10_)  &  i_12_  &  (~ i_11_) ) ;
 assign wire19288 = ( wire5990 ) | ( n_n177  &  wire19286 ) | ( n_n177  &  wire19287 ) ;
 assign n_n5017 = ( n_n5053 ) | ( n_n5051 ) | ( wire19288 ) ;
 assign wire1226 = ( i_7_  &  i_8_  &  i_6_ ) | ( (~ i_7_)  &  i_8_  &  i_6_ ) ;
 assign wire5874 = ( n_n264  &  n_n165  &  wire1226 ) ;
 assign wire5875 = ( _6995 ) | ( _6996 ) | ( _6997 ) ;
 assign wire19882 = ( n_n4834 ) | ( _5173 ) | ( _5174 ) ;
 assign n_n4633 = ( n_n6  &  wire65 ) | ( n_n6  &  wire902  &  n_n225 ) ;
 assign wire705 = ( n_n57  &  n_n108 ) | ( n_n56  &  wire60 ) ;
 assign wire1231 = ( n_n264  &  n_n229  &  n_n165 ) | ( n_n229  &  n_n165  &  n_n230 ) ;
 assign wire20719 = ( wire200  &  n_n56 ) | ( n_n56  &  wire277 ) ;
 assign wire20720 = ( wire268  &  n_n57 ) | ( wire200  &  n_n57 ) ;
 assign wire20721 = ( wire268  &  n_n56 ) | ( n_n57  &  wire277 ) ;
 assign wire20722 = ( wire112  &  n_n57 ) | ( wire112  &  n_n56 ) | ( n_n57  &  wire157 ) ;
 assign n_n4218 = ( wire20719 ) | ( wire20720 ) | ( wire20721 ) | ( wire20722 ) ;
 assign n_n4214 = ( n_n4259 ) | ( wire721 ) | ( _3878 ) | ( _37661 ) ;
 assign n_n4255 = ( wire5011 ) | ( _36959 ) ;
 assign wire20729 = ( n_n4920 ) | ( n_n4907 ) | ( n_n4922 ) | ( n_n4921 ) ;
 assign wire20733 = ( n_n4256 ) | ( wire20728 ) | ( _37666 ) ;
 assign n_n1370 = ( n_n268  &  wire55 ) | ( n_n265  &  n_n32 ) ;
 assign wire5591 = ( n_n264  &  n_n285  &  n_n263  &  n_n253 ) ;
 assign wire5592 = ( n_n264  &  n_n285  &  n_n261  &  n_n267 ) ;
 assign wire309 = ( wire5591 ) | ( wire5592 ) ;
 assign wire571 = ( n_n264  &  n_n285  &  n_n261  &  n_n275 ) ;
 assign wire737 = ( n_n264  &  n_n285  &  n_n263  &  n_n270 ) ;
 assign wire20300 = ( wire5591 ) | ( wire5592 ) | ( wire737 ) ;
 assign wire20301 = ( wire407 ) | ( wire457 ) | ( n_n53  &  wire77 ) ;
 assign wire20304 = ( n_n4183 ) | ( wire20299 ) | ( _4390 ) ;
 assign wire5510 = ( _6034 ) | ( wire137  &  n_n94 ) | ( wire132  &  n_n94 ) ;
 assign wire5514 = ( n_n100  &  wire246 ) | ( n_n100  &  wire256 ) ;
 assign wire5515 = ( wire73  &  n_n94 ) | ( n_n65  &  n_n94 ) | ( n_n94  &  wire19556 ) ;
 assign wire20155 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire911 ) | ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  wire911 ) ;
 assign n_n3598 = ( wire118  &  n_n94 ) | ( n_n220  &  wire899  &  n_n94 ) ;
 assign wire3800 = ( wire72  &  n_n100 ) | ( wire905  &  n_n258  &  n_n100 ) ;
 assign wire21083 = ( n_n226  &  n_n100 ) | ( wire208  &  n_n94 ) ;
 assign n_n3209 = ( n_n3598 ) | ( wire3800 ) | ( wire21083 ) ;
 assign wire628 = ( wire80  &  n_n100 ) | ( n_n100  &  wire69 ) | ( n_n100  &  n_n78 ) ;
 assign wire21105 = ( _3443 ) | ( _3444 ) | ( n_n31  &  n_n100 ) ;
 assign n_n4644 = ( n_n6  &  wire368 ) | ( n_n6  &  n_n247  &  _36683 ) ;
 assign n_n4636 = ( n_n5  &  wire368 ) | ( n_n5  &  n_n247  &  _36683 ) ;
 assign wire4745 = ( n_n5  &  wire71 ) | ( n_n5  &  n_n97 ) | ( n_n5  &  wire77 ) ;
 assign wire20131 = ( n_n6  &  n_n41 ) | ( n_n6  &  wire368 ) | ( n_n6  &  n_n88 ) ;
 assign wire21019 = ( n_n4636 ) | ( wire3837 ) | ( wire21017 ) ;
 assign wire21027 = ( wire389 ) | ( wire464 ) | ( wire463 ) | ( wire21021 ) ;
 assign wire21028 = ( wire21022 ) | ( wire21023 ) | ( _3550 ) ;
 assign n_n4632 = ( n_n6  &  wire80 ) | ( n_n6  &  wire902  &  n_n256 ) ;
 assign wire487 = ( n_n6  &  wire88 ) | ( n_n6  &  n_n31 ) | ( n_n6  &  n_n80 ) ;
 assign wire742 = ( n_n253  &  _35042  &  _38171 ) | ( n_n253  &  _35043  &  _38171 ) ;
 assign wire931 = ( n_n208  &  n_n285  &  n_n230  &  wire232 ) ;
 assign wire20362 = ( n_n275  &  _37442 ) | ( n_n275  &  _37444 ) ;
 assign wire20364 = ( n_n151  &  n_n6 ) | ( n_n207  &  wire232 ) ;
 assign n_n2876 = ( wire20364 ) | ( _4139 ) ;
 assign n_n3731 = ( n_n4  &  wire19407 ) | ( n_n4  &  n_n256  &  wire897 ) ;
 assign n_n1597 = ( n_n57  &  n_n104 ) | ( n_n56  &  wire78 ) ;
 assign wire3595 = ( _3041 ) | ( _3042 ) ;
 assign wire3588 = ( _3035 ) | ( _3036 ) | ( _3037 ) ;
 assign wire21318 = ( n_n1604 ) | ( _3027 ) | ( _3028 ) ;
 assign wire271 = ( i_15_  &  n_n242  &  n_n222 ) | ( (~ i_15_)  &  n_n242  &  n_n222 ) ;
 assign wire472 = ( i_15_  &  n_n222  &  n_n259 ) | ( (~ i_15_)  &  n_n222  &  n_n259 ) ;
 assign wire21723 = ( n_n57  &  wire271 ) | ( n_n56  &  wire472 ) ;
 assign wire21724 = ( n_n110  &  n_n57 ) | ( n_n110  &  n_n56 ) | ( n_n57  &  wire247 ) ;
 assign n_n1788 = ( wire21723 ) | ( wire21724 ) ;
 assign wire21713 = ( n_n56  &  n_n22 ) | ( n_n57  &  wire426 ) ;
 assign wire21714 = ( n_n57  &  wire212 ) | ( n_n56  &  wire212 ) ;
 assign wire21718 = ( wire21716 ) | ( n_n56  &  n_n76 ) | ( n_n56  &  wire165 ) ;
 assign wire21719 = ( wire3109 ) | ( n_n56  &  wire247 ) | ( n_n56  &  wire21715 ) ;
 assign n_n1715 = ( wire21713 ) | ( wire21714 ) | ( wire21718 ) | ( wire21719 ) ;
 assign wire1250 = ( n_n220  &  wire911 ) | ( n_n220  &  wire912 ) | ( n_n220  &  wire902 ) ;
 assign wire1249 = ( n_n220  &  wire902 ) | ( n_n220  &  wire899 ) ;
 assign wire1248 = ( n_n220  &  wire901 ) | ( n_n220  &  wire897 ) ;
 assign wire21729 = ( n_n111  &  n_n56 ) | ( n_n57  &  n_n76 ) ;
 assign wire21730 = ( n_n56  &  wire426 ) | ( n_n57  &  wire379 ) ;
 assign n_n1792 = ( wire21729 ) | ( wire21730 ) | ( n_n57  &  wire165 ) ;
 assign wire158 = ( i_15_  &  n_n282  &  n_n222 ) | ( (~ i_15_)  &  n_n282  &  n_n222 ) ;
 assign wire1251 = ( i_15_  &  n_n282  &  n_n222 ) | ( (~ i_15_)  &  n_n282  &  n_n222 ) | ( i_15_  &  n_n222  &  n_n247 ) | ( (~ i_15_)  &  n_n222  &  n_n247 ) ;
 assign wire21728 = ( wire3098 ) | ( wire3106 ) | ( wire21721 ) | ( wire21726 ) ;
 assign wire21739 = ( n_n1792 ) | ( wire3080 ) | ( wire21733 ) | ( wire21737 ) ;
 assign n_n1690 = ( n_n1788 ) | ( n_n1715 ) | ( wire21728 ) | ( wire21739 ) ;
 assign n_n1440 = ( n_n3  &  wire68 ) | ( n_n4  &  n_n42 ) ;
 assign wire300 = ( i_15_  &  n_n281  &  n_n267 ) | ( i_15_  &  n_n256  &  n_n267 ) | ( (~ i_15_)  &  n_n256  &  n_n267 ) ;
 assign n_n1173 = ( n_n1440 ) | ( _1801 ) | ( wire41  &  _39406 ) ;
 assign wire2740 = ( n_n4  &  wire66 ) | ( n_n4  &  wire42 ) | ( n_n4  &  n_n20 ) ;
 assign wire22064 = ( n_n4  &  n_n258  &  wire899 ) | ( n_n4  &  n_n222  &  wire899 ) ;
 assign n_n1210 = ( wire466 ) | ( wire2740 ) | ( wire22064 ) ;
 assign n_n6820 = ( wire911  &  n_n225  &  n_n94 ) ;
 assign wire1253 = ( n_n228  &  wire902 ) | ( n_n228  &  wire899 ) ;
 assign wire22765 = ( wire911  &  n_n279 ) | ( n_n225  &  wire903 ) ;
 assign wire22766 = ( i_14_  &  i_13_  &  i_12_  &  wire913 ) | ( (~ i_14_)  &  i_13_  &  i_12_  &  wire913 ) ;
 assign wire1254 = ( wire60 ) | ( n_n68 ) | ( wire22765 ) | ( wire22766 ) ;
 assign wire320 = ( n_n275  &  _40264 ) | ( n_n275  &  _40265 ) ;
 assign wire22335 = ( n_n275  &  _40268 ) | ( n_n275  &  _40269 ) ;
 assign n_n370 = ( _719 ) | ( _720 ) | ( _721 ) | ( _40313 ) ;
 assign wire276 = ( n_n270  &  _40217 ) | ( n_n270  &  _40218 ) ;
 assign wire182 = ( i_15_  &  n_n256  &  n_n270 ) | ( (~ i_15_)  &  n_n256  &  n_n270 ) ;
 assign wire405 = ( (~ i_15_)  &  n_n279  &  n_n275 ) | ( i_15_  &  n_n256  &  n_n275 ) | ( (~ i_15_)  &  n_n256  &  n_n275 ) ;
 assign wire22477 = ( i_14_  &  i_13_  &  (~ i_12_)  &  wire908 ) | ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire908 ) ;
 assign wire1259 = ( wire276 ) | ( wire182 ) | ( wire405 ) | ( wire22477 ) ;
 assign wire2304 = ( _705 ) | ( _706 ) | ( n_n56  &  wire22475 ) ;
 assign wire2305 = ( _702 ) | ( _703 ) ;
 assign wire2296 = ( wire166  &  n_n94 ) | ( n_n94  &  wire229 ) ;
 assign wire22483 = ( wire166  &  n_n100 ) | ( n_n258  &  wire900  &  n_n100 ) ;
 assign wire22487 = ( wire2291 ) | ( _675 ) ;
 assign wire877 = ( n_n83  &  n_n100 ) | ( n_n100  &  n_n36 ) | ( n_n100  &  n_n35 ) ;
 assign wire2277 = ( n_n256  &  n_n94  &  _40373 ) | ( n_n256  &  n_n94  &  _40375 ) ;
 assign wire22495 = ( n_n94  &  n_n41 ) | ( n_n100  &  n_n81 ) ;
 assign wire22496 = ( n_n258  &  wire901  &  n_n100 ) | ( wire901  &  n_n256  &  n_n100 ) ;
 assign n_n464 = ( wire877 ) | ( wire2277 ) | ( wire22495 ) | ( wire22496 ) ;
 assign wire688 = ( wire914  &  n_n256  &  n_n94 ) | ( wire912  &  n_n256  &  n_n94 ) ;
 assign wire358 = ( i_15_  &  n_n256  &  n_n247 ) | ( (~ i_15_)  &  n_n256  &  n_n247 ) ;
 assign wire1261 = ( wire57 ) | ( wire140 ) | ( n_n113 ) | ( wire358 ) ;
 assign wire22493 = ( wire22240 ) | ( wire22241 ) | ( wire22242 ) | ( wire22491 ) ;
 assign wire22494 = ( wire22492 ) | ( _654 ) | ( _655 ) ;
 assign wire22504 = ( n_n464 ) | ( wire22502 ) | ( n_n100  &  wire1261 ) ;
 assign wire5988 = ( i_5_  &  i_3_  &  n_n165  &  wire19291 ) ;
 assign n_n5048 = ( _6700 ) | ( _34842 ) ;
 assign wire315 = ( i_9_ ) | ( (~ i_9_)  &  i_10_ ) ;
 assign wire1265 = ( n_n165  &  n_n283  &  wire19294 ) | ( n_n165  &  n_n283  &  wire19296 ) ;
 assign wire1264 = ( n_n165  &  n_n273  &  wire19294 ) | ( n_n165  &  n_n273  &  wire19296 ) ;
 assign wire326 = ( (~ i_15_)  &  n_n281  &  n_n242 ) | ( i_15_  &  n_n242  &  n_n279 ) ;
 assign wire19260 = ( _6865 ) | ( _6866 ) | ( n_n130  &  _34687 ) ;
 assign wire19261 = ( wire5953 ) | ( _6848 ) | ( _6849 ) ;
 assign wire19263 = ( wire19243 ) | ( wire19250 ) | ( _34724 ) ;
 assign n_n4911 = ( n_n110  &  n_n57 ) | ( n_n56  &  wire82 ) ;
 assign n_n3736 = ( n_n4  &  wire80 ) | ( n_n4  &  wire908  &  n_n256 ) ;
 assign n_n1339 = ( n_n4  &  n_n76 ) | ( n_n3  &  wire56 ) ;
 assign n_n3579 = ( n_n65  &  n_n48 ) | ( wire44  &  n_n53 ) ;
 assign n_n4674 = ( n_n56  &  wire71 ) | ( n_n56  &  n_n256  &  wire904 ) ;
 assign wire3830 = ( n_n49  &  n_n48 ) | ( n_n48  &  wire71 ) | ( n_n48  &  wire68 ) ;
 assign wire3831 = ( n_n95  &  n_n53 ) | ( n_n53  &  n_n179 ) | ( n_n53  &  wire57 ) ;
 assign wire4492 = ( n_n207  &  n_n17 ) | ( n_n207  &  wire514 ) | ( n_n207  &  wire20365 ) ;
 assign wire20366 = ( n_n207  &  _37448 ) | ( wire913  &  n_n207  &  _36156 ) ;
 assign wire20367 = ( n_n104  &  n_n100 ) | ( n_n9  &  n_n207 ) ;
 assign n_n2875 = ( wire4492 ) | ( wire20366 ) | ( wire20367 ) ;
 assign wire3316 = ( n_n5  &  n_n93 ) | ( n_n5  &  n_n90 ) | ( n_n5  &  wire21389 ) ;
 assign wire3317 = ( n_n6  &  wire71 ) | ( n_n6  &  n_n279  &  wire904 ) ;
 assign n_n2145 = ( wire389 ) | ( wire3316 ) | ( wire3317 ) ;
 assign wire226 = ( n_n253  &  _38941 ) | ( n_n253  &  _38942 ) ;
 assign wire21832 = ( n_n48  &  n_n47 ) | ( n_n57  &  n_n150 ) ;
 assign n_n1785 = ( wire21832 ) | ( _2230 ) | ( n_n56  &  _39096 ) ;
 assign wire1291 = ( n_n220  &  wire912 ) | ( n_n220  &  wire898 ) | ( n_n220  &  wire897 ) ;
 assign wire1290 = ( n_n220  &  wire912 ) | ( n_n220  &  wire902 ) ;
 assign wire1289 = ( n_n220  &  wire901 ) | ( n_n220  &  wire900 ) ;
 assign wire2566 = ( wire154  &  n_n100 ) | ( wire64  &  n_n100 ) ;
 assign wire22231 = ( wire907  &  n_n279  &  n_n100 ) | ( wire907  &  n_n256  &  n_n100 ) ;
 assign wire22232 = ( n_n94  &  n_n41 ) | ( n_n94  &  n_n88 ) | ( n_n94  &  n_n87 ) ;
 assign wire687 = ( n_n94  &  wire50 ) | ( wire912  &  n_n256  &  n_n94 ) ;
 assign wire22066 = ( n_n10  &  n_n100 ) | ( n_n94  &  n_n39 ) ;
 assign wire22067 = ( n_n94  &  _39853 ) | ( wire911  &  n_n94  &  _34546 ) ;
 assign n_n1212 = ( wire825 ) | ( wire687 ) | ( wire22066 ) | ( wire22067 ) ;
 assign wire374 = ( n_n4  &  wire902  &  n_n258 ) | ( n_n4  &  wire902  &  n_n222 ) ;
 assign wire434 = ( wire907  &  n_n228  &  n_n100 ) | ( wire907  &  n_n279  &  n_n100 ) ;
 assign wire799 = ( n_n4  &  wire140 ) | ( n_n4  &  wire165 ) ;
 assign wire22075 = ( wire696 ) | ( wire548 ) | ( wire374 ) | ( wire434 ) ;
 assign wire22076 = ( wire799 ) | ( wire22070 ) | ( wire22071 ) ;
 assign n_n1123 = ( n_n1212 ) | ( wire22075 ) | ( wire22076 ) ;
 assign wire20755 = ( n_n177  &  n_n112 ) | ( n_n189  &  n_n109 ) ;
 assign wire229 = ( i_15_  &  n_n256  &  n_n267 ) | ( (~ i_15_)  &  n_n256  &  n_n267 ) ;
 assign n_n5664 = ( (~ i_7_)  &  (~ i_6_)  &  n_n118  &  n_n230 ) ;
 assign wire793 = ( i_7_  &  i_6_  &  n_n116  &  n_n230 ) | ( i_7_  &  (~ i_6_)  &  n_n116  &  n_n230 ) ;
 assign wire22240 = ( n_n255  &  n_n197 ) | ( n_n241  &  n_n104 ) ;
 assign wire22241 = ( n_n189  &  n_n113 ) | ( n_n177  &  n_n35 ) ;
 assign wire22242 = ( n_n241  &  n_n216 ) | ( n_n255  &  n_n41 ) ;
 assign wire1307 = ( wire913  &  n_n281 ) | ( n_n281  &  wire914 ) ;
 assign wire22512 = ( wire912  &  n_n258 ) | ( wire902  &  n_n258 ) ;
 assign wire22513 = ( i_15_  &  n_n256  &  n_n247 ) | ( (~ i_15_)  &  n_n256  &  n_n247 ) | ( i_15_  &  n_n256  &  n_n275 ) | ( (~ i_15_)  &  n_n256  &  n_n275 ) ;
 assign wire1311 = ( wire57 ) | ( n_n113 ) | ( wire22512 ) | ( wire22513 ) ;
 assign wire2258 = ( n_n2  &  n_n34 ) | ( n_n2  &  wire47 ) | ( n_n2  &  wire22519 ) ;
 assign wire624 = ( wire905  &  n_n256  &  n_n53 ) | ( wire899  &  n_n256  &  n_n53 ) ;
 assign wire233 = ( n_n282  &  _40015 ) | ( n_n282  &  _40016 ) ;
 assign wire22522 = ( n_n61  &  n_n53 ) | ( n_n257  &  n_n53 ) | ( n_n53  &  wire123 ) ;
 assign n_n408 = ( wire624 ) | ( wire22522 ) | ( n_n2  &  wire233 ) ;
 assign wire22524 = ( wire2246 ) | ( n_n2  &  wire166 ) | ( n_n2  &  wire22523 ) ;
 assign wire22527 = ( wire22511 ) | ( wire22518 ) | ( _40056 ) ;
 assign wire19909 = ( n_n4287 ) | ( n_n4892 ) | ( wire5023 ) ;
 assign n_n4736 = ( wire5033 ) | ( wire19909 ) | ( _5135 ) | ( _36515 ) ;
 assign wire481 = ( n_n220  &  wire905  &  n_n57 ) | ( wire905  &  n_n57  &  n_n256 ) ;
 assign n_n4913 = ( n_n57  &  wire84 ) | ( wire913  &  n_n279  &  n_n57 ) ;
 assign n_n4259 = ( n_n4912 ) | ( n_n4911 ) | ( n_n4913 ) ;
 assign n_n4915 = ( n_n110  &  n_n56 ) | ( n_n57  &  wire60 ) ;
 assign n_n4914 = ( n_n57  &  wire52 ) | ( wire911  &  n_n279  &  n_n57 ) ;
 assign wire721 = ( n_n4916 ) | ( n_n4915 ) | ( n_n4914 ) ;
 assign wire5589 = ( n_n56  &  wire70 ) | ( n_n56  &  wire44 ) ;
 assign wire20121 = ( n_n57  &  wire73 ) | ( n_n57  &  n_n65 ) | ( n_n57  &  n_n11 ) ;
 assign n_n4256 = ( wire5589 ) | ( wire20121 ) | ( n_n57  &  n_n12 ) ;
 assign wire101 = ( n_n282  &  _35947 ) | ( n_n282  &  _35948 ) ;
 assign wire5011 = ( n_n106  &  n_n56 ) | ( n_n56  &  n_n62 ) | ( n_n56  &  wire101 ) ;
 assign wire5552 = ( n_n56  &  wire73 ) | ( n_n56  &  n_n65 ) | ( n_n56  &  n_n12 ) ;
 assign wire465 = ( wire5552 ) | ( n_n57  &  wire44 ) ;
 assign wire5613 = ( n_n6  &  wire41 ) | ( n_n6  &  n_n279  &  wire898 ) ;
 assign n_n3786 = ( n_n1  &  n_n95 ) | ( n_n2  &  wire81 ) ;
 assign n_n3782 = ( n_n2  &  n_n42 ) | ( n_n1  &  wire81 ) ;
 assign wire723 = ( n_n2  &  wire19385 ) | ( n_n2  &  n_n256  &  wire900 ) ;
 assign wire19384 = ( (~ i_14_)  &  i_13_  &  i_12_  &  wire906 ) | ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire906 ) ;
 assign wire19440 = ( n_n3781 ) | ( n_n3786 ) | ( _6280 ) ;
 assign n_n4676 = ( n_n56  &  wire96 ) | ( n_n56  &  n_n222  &  wire904 ) ;
 assign n_n4686 = ( n_n57  &  wire71 ) | ( n_n57  &  n_n256  &  wire904 ) ;
 assign wire1322 = ( wire912  &  n_n258 ) | ( wire902  &  n_n258 ) | ( n_n258  &  wire898 ) ;
 assign wire3764 = ( n_n260  &  n_n285  &  n_n271  &  wire1322 ) ;
 assign wire21108 = ( n_n255  &  n_n197 ) | ( n_n189  &  n_n109 ) ;
 assign wire21109 = ( wire914  &  n_n279  &  n_n189 ) | ( n_n279  &  n_n189  &  wire904 ) ;
 assign wire21110 = ( n_n54  &  n_n100 ) | ( n_n189  &  n_n101 ) ;
 assign n_n3221 = ( wire3764 ) | ( wire21108 ) | ( wire21109 ) | ( wire21110 ) ;
 assign wire1323 = ( i_9_  &  i_10_  &  i_11_ ) | ( i_9_  &  (~ i_10_)  &  i_11_ ) | ( i_9_  &  (~ i_10_)  &  (~ i_11_) ) ;
 assign wire21046 = ( wire5031 ) | ( wire21043 ) | ( n_n60  &  n_n56 ) ;
 assign wire21047 = ( n_n4892 ) | ( wire4056 ) | ( wire20826 ) | ( wire21042 ) ;
 assign wire298 = ( _4514 ) | ( n_n53  &  n_n31 ) | ( n_n53  &  n_n80 ) ;
 assign n_n5675 = ( i_7_  &  i_6_  &  n_n116  &  n_n284 ) ;
 assign wire1327 = ( i_15_  &  n_n279  &  n_n247 ) | ( (~ i_15_)  &  n_n279  &  n_n247 ) | ( (~ i_15_)  &  n_n225  &  n_n247 ) ;
 assign wire3303 = ( n_n264  &  n_n285  &  n_n283  &  wire1327 ) ;
 assign wire21565 = ( n_n106  &  n_n53 ) | ( n_n48  &  n_n148 ) ;
 assign wire21566 = ( n_n6  &  n_n186 ) | ( n_n48  &  n_n135 ) ;
 assign n_n2146 = ( wire462 ) | ( wire3303 ) | ( wire21565 ) | ( wire21566 ) ;
 assign wire429 = ( i_15_  &  n_n222  &  n_n247 ) | ( (~ i_15_)  &  n_n222  &  n_n247 ) ;
 assign wire263 = ( n_n247  &  _38978 ) | ( n_n247  &  _38979 ) ;
 assign wire1329 = ( wire102 ) | ( wire263 ) | ( wire912  &  n_n256 ) ;
 assign wire1330 = ( n_n220  &  wire898 ) | ( n_n220  &  wire897 ) ;
 assign wire21770 = ( n_n8  &  n_n53 ) | ( n_n48  &  n_n147 ) ;
 assign wire21771 = ( n_n53  &  n_n147 ) | ( n_n48  &  n_n62 ) | ( n_n53  &  n_n62 ) ;
 assign wire21772 = ( n_n48  &  n_n64 ) | ( n_n53  &  n_n64 ) | ( n_n48  &  wire1330 ) ;
 assign n_n1774 = ( wire21770 ) | ( wire21771 ) | ( wire21772 ) ;
 assign wire3032 = ( _39274 ) | ( n_n53  &  wire195 ) | ( n_n53  &  _39273 ) ;
 assign wire3033 = ( _1997 ) | ( _1998 ) ;
 assign wire1333 = ( n_n275  &  _39703 ) | ( n_n275  &  _39704 ) ;
 assign wire22187 = ( n_n94  &  _39702 ) | ( wire903  &  n_n94  &  _36705 ) ;
 assign wire22188 = ( n_n94  &  n_n200 ) | ( n_n94  &  n_n24 ) | ( n_n94  &  wire1333 ) ;
 assign wire1334 = ( n_n247  &  _39707 ) | ( n_n247  &  _39708 ) ;
 assign n_n3884 = ( n_n100  &  wire19577 ) | ( n_n228  &  wire906  &  n_n100 ) ;
 assign wire580 = ( n_n227  &  wire22795 ) | ( n_n228  &  wire897  &  n_n227 ) ;
 assign wire22796 = ( n_n9  &  n_n207 ) | ( n_n94  &  n_n203 ) ;
 assign wire22797 = ( n_n9  &  n_n227 ) | ( n_n207  &  n_n59 ) ;
 assign n_n809 = ( wire931 ) | ( wire580 ) | ( wire22796 ) | ( wire22797 ) ;
 assign wire1340 = ( i_15_  &  n_n282  &  n_n225 ) | ( (~ i_15_)  &  n_n282  &  n_n225 ) | ( i_15_  &  n_n225  &  n_n247 ) | ( (~ i_15_)  &  n_n225  &  n_n247 ) ;
 assign wire1343 = ( i_15_  &  n_n282  &  n_n225 ) | ( (~ i_15_)  &  n_n282  &  n_n225 ) | ( i_15_  &  n_n225  &  n_n247 ) | ( (~ i_15_)  &  n_n225  &  n_n247 ) ;
 assign wire1344 = ( wire907  &  n_n258 ) | ( n_n258  &  wire903 ) ;
 assign wire22363 = ( n_n258  &  wire906 ) | ( wire905  &  n_n256 ) ;
 assign wire408 = ( n_n267  &  _40066 ) | ( n_n267  &  _40067 ) ;
 assign wire933 = ( wire913  &  n_n268  &  n_n258 ) ;
 assign wire414 = ( (~ i_15_)  &  n_n279  &  n_n282 ) | ( i_15_  &  n_n282  &  n_n256 ) | ( (~ i_15_)  &  n_n282  &  n_n256 ) ;
 assign wire357 = ( n_n253  &  _40068 ) | ( n_n253  &  _40069 ) ;
 assign wire22340 = ( n_n253  &  _40070 ) | ( n_n253  &  _40071 ) ;
 assign wire22533 = ( wire22532 ) | ( _1054 ) ;
 assign wire1354 = ( i_8_  &  n_n260  &  n_n285  &  n_n155 ) | ( (~ i_8_)  &  n_n260  &  n_n285  &  n_n155 ) ;
 assign wire1357 = ( wire914  &  n_n258 ) | ( n_n258  &  wire904 ) ;
 assign wire1355 = ( wire907  &  n_n258 ) | ( n_n258  &  wire906 ) ;
 assign wire22537 = ( wire2237 ) | ( wire2239 ) | ( wire2240 ) ;
 assign wire419 = ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  wire914 ) | ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire914 ) ;
 assign wire19604 = ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  wire913 ) | ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire913 ) ;
 assign wire20344 = ( n_n220  &  wire908  &  n_n53 ) | ( wire908  &  n_n256  &  n_n53 ) ;
 assign n_n4146 = ( wire478 ) | ( wire406 ) | ( n_n3587 ) | ( wire20344 ) ;
 assign wire20253 = ( wire376 ) | ( wire462 ) | ( wire464 ) | ( wire20248 ) ;
 assign wire20254 = ( n_n4094 ) | ( n_n4124 ) | ( n_n4090 ) | ( wire483 ) ;
 assign n_n3925 = ( wire470 ) | ( wire4602 ) | ( wire20253 ) | ( wire20254 ) ;
 assign wire21250 = ( n_n4068 ) | ( n_n4069 ) | ( wire21248 ) ;
 assign wire3707 = ( n_n3  &  n_n7 ) | ( n_n3  &  wire50 ) | ( n_n3  &  n_n59 ) ;
 assign wire3708 = ( n_n4  &  wire50 ) | ( n_n228  &  n_n4  &  wire897 ) ;
 assign wire21188 = ( n_n4  &  _38311 ) | ( n_n4  &  wire902  &  _35049 ) ;
 assign n_n3930 = ( wire3707 ) | ( wire3708 ) | ( wire21188 ) ;
 assign wire3702 = ( n_n3  &  wire208 ) | ( n_n3  &  wire199 ) ;
 assign wire21190 = ( n_n4  &  _38296 ) | ( n_n4  &  wire899  &  _37091 ) ;
 assign wire21191 = ( n_n4  &  n_n145 ) | ( n_n4  &  n_n7 ) | ( n_n4  &  n_n144 ) ;
 assign n_n3929 = ( wire3702 ) | ( wire21190 ) | ( wire21191 ) ;
 assign wire4587 = ( n_n53  &  wire74 ) | ( n_n225  &  n_n53  &  wire903 ) ;
 assign wire20259 = ( n_n53  &  n_n197 ) | ( n_n48  &  wire69 ) ;
 assign wire20262 = ( n_n4168 ) | ( wire4593 ) | ( wire20257 ) | ( n_n4073 ) ;
 assign wire20271 = ( wire20268 ) | ( wire20269 ) | ( _4469 ) | ( _37143 ) ;
 assign n_n3980 = ( n_n4160 ) | ( wire4565 ) | ( wire20275 ) ;
 assign wire20282 = ( wire882 ) | ( wire20277 ) | ( wire20278 ) | ( wire20279 ) ;
 assign n_n3920 = ( n_n3978 ) | ( n_n3980 ) | ( wire20282 ) ;
 assign wire4558 = ( _4426 ) | ( n_n48  &  n_n16 ) | ( n_n48  &  wire20155 ) ;
 assign wire20287 = ( wire456 ) | ( n_n4165 ) | ( wire20285 ) ;
 assign n_n3922 = ( wire4558 ) | ( wire20287 ) | ( _4429 ) | ( _37170 ) ;
 assign wire4552 = ( _4412 ) | ( _4413 ) | ( _4414 ) ;
 assign wire20293 = ( wire675 ) | ( wire4551 ) | ( wire4573 ) | ( wire4574 ) ;
 assign wire4530 = ( _4376 ) | ( _4377 ) ;
 assign wire20310 = ( wire912  &  n_n258  &  n_n53 ) | ( n_n258  &  wire901  &  n_n53 ) ;
 assign wire20319 = ( _4365 ) | ( _4366 ) | ( _37230 ) ;
 assign wire59 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire900 ) | ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  wire900 ) ;
 assign wire19582 = ( n_n3881 ) | ( _5925 ) | ( n_n105  &  n_n100 ) ;
 assign wire4131 = ( wire66  &  n_n100 ) | ( wire905  &  n_n222  &  n_n100 ) ;
 assign wire20756 = ( n_n197  &  n_n100 ) | ( n_n94  &  wire77 ) ;
 assign n_n3486 = ( n_n3610 ) | ( wire4131 ) | ( wire20756 ) ;
 assign wire20764 = ( wire20758 ) | ( wire20760 ) | ( n_n100  &  wire83 ) ;
 assign wire20765 = ( n_n1628 ) | ( n_n1058 ) | ( wire4120 ) | ( wire20759 ) ;
 assign n_n3403 = ( n_n3486 ) | ( wire20764 ) | ( wire20765 ) ;
 assign n_n3372 = ( n_n3403 ) | ( _35721 ) | ( _35722 ) | ( _37751 ) ;
 assign wire225 = ( i_15_  &  n_n228  &  n_n242 ) | ( (~ i_15_)  &  n_n242  &  n_n258 ) ;
 assign n_n2713 = ( n_n145  &  n_n100 ) | ( n_n94  &  wire225 ) ;
 assign wire5506 = ( n_n57  &  wire96 ) | ( n_n57  &  n_n222  &  wire904 ) ;
 assign wire370 = ( wire863 ) | ( n_n4687 ) | ( wire5506 ) ;
 assign wire130 = ( n_n242  &  _34536 ) | ( n_n242  &  _34537 ) ;
 assign wire4789 = ( n_n151  &  n_n100 ) | ( wire75  &  n_n100 ) | ( n_n206  &  n_n100 ) ;
 assign wire20775 = ( n_n1624 ) | ( n_n3604 ) | ( wire4117 ) | ( wire20772 ) ;
 assign wire20782 = ( wire370 ) | ( wire4789 ) | ( wire4790 ) | ( wire20779 ) ;
 assign n_n3371 = ( wire20782 ) | ( wire19565 ) | ( _37764 ) | ( _37772 ) ;
 assign wire19936 = ( n_n4920 ) | ( n_n4921 ) | ( n_n4916 ) | ( wire705 ) ;
 assign wire19914 = ( n_n4907 ) | ( _5118 ) | ( _5119 ) ;
 assign n_n3397 = ( n_n4781 ) | ( n_n4912 ) | ( n_n4911 ) | ( wire19914 ) ;
 assign wire788 = ( n_n56  &  n_n95 ) | ( n_n56  &  n_n49 ) | ( n_n56  &  wire71 ) ;
 assign wire21077 = ( n_n56  &  wire68 ) | ( n_n57  &  wire55 ) ;
 assign wire21081 = ( n_n4675 ) | ( n_n4676 ) | ( n_n4686 ) | ( wire21076 ) ;
 assign wire20374 = ( wire434 ) | ( wire20369 ) | ( wire20370 ) | ( wire20371 ) ;
 assign wire20376 = ( n_n281  &  wire906 ) | ( n_n228  &  wire901 ) ;
 assign wire1371 = ( wire132 ) | ( wire160 ) | ( wire184 ) | ( wire20376 ) ;
 assign wire20381 = ( wire20379 ) | ( n_n6  &  wire1371 ) ;
 assign wire20382 = ( n_n4823 ) | ( n_n4605 ) | ( wire4506 ) | ( wire20356 ) ;
 assign wire21389 = ( (~ i_14_)  &  i_13_  &  i_12_  &  wire906 ) | ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire906 ) ;
 assign n_n2158 = ( _2854 ) | ( n_n48  &  wire51 ) | ( n_n48  &  _38545 ) ;
 assign wire1378 = ( wire913  &  n_n281 ) | ( n_n281  &  wire905 ) | ( n_n281  &  wire908 ) ;
 assign wire1377 = ( i_8_  &  n_n153  &  n_n285  &  n_n230 ) | ( (~ i_8_)  &  n_n153  &  n_n285  &  n_n230 ) ;
 assign n_n4682 = ( n_n56  &  wire19384 ) | ( n_n281  &  n_n56  &  wire900 ) ;
 assign wire21445 = ( n_n281  &  wire905  &  n_n100 ) | ( n_n281  &  wire905  &  n_n94 ) ;
 assign wire21446 = ( n_n151  &  wire168 ) | ( n_n57  &  wire482 ) ;
 assign n_n2172 = ( n_n4686 ) | ( wire21445 ) | ( wire21446 ) ;
 assign wire482 = ( i_15_  &  n_n279  &  n_n253 ) | ( (~ i_15_)  &  n_n279  &  n_n253 ) ;
 assign wire1379 = ( i_15_  &  n_n279  &  n_n267 ) | ( (~ i_15_)  &  n_n279  &  n_n267 ) ;
 assign wire3452 = ( n_n57  &  wire19384 ) | ( n_n281  &  n_n57  &  wire900 ) ;
 assign wire21449 = ( n_n57  &  n_n42 ) | ( n_n57  &  wire1379 ) | ( n_n56  &  wire1379 ) ;
 assign wire21453 = ( n_n4674 ) | ( n_n4682 ) | ( wire3451 ) | ( wire21448 ) ;
 assign n_n2093 = ( n_n2172 ) | ( wire3452 ) | ( wire21449 ) | ( wire21453 ) ;
 assign wire86 = ( i_15_  &  n_n281  &  n_n282 ) | ( (~ i_15_)  &  n_n282  &  n_n225 ) ;
 assign n_n4666 = ( n_n57  &  wire86 ) | ( wire907  &  n_n57  &  n_n256 ) ;
 assign wire1383 = ( i_15_  &  n_n279  &  n_n282 ) | ( (~ i_15_)  &  n_n279  &  n_n282 ) | ( i_15_  &  n_n279  &  n_n270 ) | ( (~ i_15_)  &  n_n279  &  n_n270 ) ;
 assign wire21462 = ( n_n2398 ) | ( wire3441 ) | ( wire3442 ) | ( wire21459 ) ;
 assign wire21463 = ( wire3440 ) | ( wire3447 ) | ( wire21455 ) ;
 assign wire21470 = ( n_n2169 ) | ( _2888 ) | ( _38513 ) | ( _38522 ) ;
 assign wire425 = ( (~ i_14_)  &  i_13_  &  i_12_  &  wire897 ) | ( i_14_  &  i_13_  &  (~ i_12_)  &  wire897 ) ;
 assign wire657 = ( n_n94  &  wire228 ) | ( n_n256  &  n_n94  &  wire897 ) ;
 assign wire2939 = ( n_n100  &  wire230 ) | ( wire902  &  n_n256  &  n_n100 ) ;
 assign wire21857 = ( n_n94  &  wire425 ) | ( n_n222  &  wire903  &  n_n94 ) ;
 assign n_n1804 = ( wire657 ) | ( wire2939 ) | ( wire21857 ) ;
 assign wire448 = ( (~ i_15_)  &  n_n228  &  n_n267 ) | ( i_15_  &  n_n222  &  n_n267 ) | ( (~ i_15_)  &  n_n222  &  n_n267 ) ;
 assign wire2745 = ( n_n1  &  wire22058 ) | ( n_n1  &  wire22059 ) ;
 assign wire22061 = ( n_n3778 ) | ( _1305 ) | ( _1306 ) ;
 assign n_n1092 = ( n_n1120 ) | ( n_n1121 ) | ( wire2745 ) | ( wire22061 ) ;
 assign wire1491 = ( wire200 ) | ( wire112 ) | ( n_n79 ) | ( wire21930 ) ;
 assign wire21935 = ( n_n1341 ) | ( n_n1346 ) | ( wire21933 ) ;
 assign n_n1108 = ( wire21935 ) | ( _1737 ) | ( _1743 ) | ( _1744 ) ;
 assign wire1492 = ( wire67 ) | ( wire85 ) | ( n_n135 ) | ( wire347 ) ;
 assign wire21941 = ( n_n3242 ) | ( wire476 ) | ( n_n1356 ) | ( wire3662 ) ;
 assign wire519 = ( n_n3  &  wire40 ) | ( n_n4  &  n_n103 ) ;
 assign wire22625 = ( n_n4954 ) | ( wire2128 ) | ( n_n56  &  wire254 ) ;
 assign wire22626 = ( wire2129 ) | ( n_n57  &  wire277 ) | ( n_n56  &  wire277 ) ;
 assign wire22646 = ( wire2103 ) | ( wire2104 ) | ( wire22642 ) | ( wire22643 ) ;
 assign n_n742 = ( wire22646 ) | ( wire22639 ) | ( wire22640 ) | ( _40728 ) ;
 assign wire139 = ( i_15_  &  n_n225  &  n_n267 ) | ( (~ i_15_)  &  n_n225  &  n_n267 ) ;
 assign wire776 = ( n_n105  &  n_n94 ) | ( n_n46  &  n_n94 ) | ( n_n94  &  wire19577 ) ;
 assign wire22662 = ( n_n1066 ) | ( wire2082 ) | ( wire22658 ) ;
 assign wire22663 = ( wire767 ) | ( wire2081 ) | ( wire2089 ) | ( wire22659 ) ;
 assign wire22670 = ( wire19380 ) | ( wire19379 ) | ( wire22667 ) | ( wire22668 ) ;
 assign n_n744 = ( n_n772 ) | ( wire22662 ) | ( wire22663 ) | ( wire22670 ) ;
 assign n_n5679 = ( i_7_  &  i_6_  &  n_n116  &  n_n230 ) ;
 assign wire321 = ( n_n279  &  n_n247 ) | ( n_n247  &  _34594 ) ;
 assign wire331 = ( wire196 ) | ( i_13_  &  (~ i_12_)  &  n_n247 ) ;
 assign wire19319 = ( wire287 ) | ( n_n281  &  wire911 ) ;
 assign wire19320 = ( wire19318 ) | ( n_n242  &  wire152 ) ;
 assign wire1400 = ( wire321 ) | ( wire331 ) | ( wire19319 ) | ( wire19320 ) ;
 assign wire546 = ( n_n4  &  _35392 ) | ( n_n4  &  wire906  &  _35394 ) ;
 assign wire634 = ( n_n3  &  n_n66 ) | ( n_n4  &  n_n64 ) ;
 assign wire21257 = ( wire349 ) | ( wire546 ) | ( wire634 ) | ( wire19400 ) ;
 assign wire21258 = ( n_n4076 ) | ( wire483 ) | ( wire21252 ) | ( wire21253 ) ;
 assign wire4089 = ( n_n151  &  n_n3 ) | ( wire75  &  n_n3 ) | ( n_n206  &  n_n3 ) ;
 assign wire4090 = ( n_n4  &  wire225 ) | ( n_n4  &  wire130 ) ;
 assign n_n3406 = ( wire4089 ) | ( wire4090 ) | ( n_n3  &  n_n226 ) ;
 assign wire3698 = ( n_n3  &  wire113 ) | ( n_n3  &  wire101 ) ;
 assign wire21193 = ( n_n4  &  _38299 ) | ( wire914  &  n_n4  &  _34565 ) ;
 assign n_n3932 = ( n_n4015 ) | ( wire3698 ) | ( wire21193 ) ;
 assign wire21200 = ( wire546 ) | ( wire3688 ) | ( wire21195 ) ;
 assign wire21201 = ( wire3689 ) | ( wire21196 ) | ( wire21197 ) ;
 assign n_n3904 = ( n_n3932 ) | ( wire21200 ) | ( wire21201 ) ;
 assign n_n3806 = ( n_n6  &  wire208 ) | ( n_n5  &  n_n59 ) ;
 assign wire5780 = ( n_n3  &  wire73 ) | ( n_n3  &  n_n65 ) | ( n_n3  &  n_n12 ) ;
 assign wire19381 = ( n_n4  &  wire44 ) | ( n_n220  &  n_n4  &  wire900 ) ;
 assign n_n3408 = ( wire546 ) | ( wire5780 ) | ( wire19381 ) ;
 assign wire20793 = ( n_n1320 ) | ( n_n3229 ) | ( wire4081 ) ;
 assign n_n3374 = ( n_n3408 ) | ( wire20793 ) | ( _3636 ) | ( _37901 ) ;
 assign wire20798 = ( wire4302 ) | ( n_n4  &  n_n108 ) | ( n_n4  &  n_n70 ) ;
 assign wire19400 = ( n_n4  &  n_n12 ) | ( n_n3  &  n_n252 ) ;
 assign wire19401 = ( n_n3  &  _35478 ) | ( n_n3  &  wire898  &  _35480 ) ;
 assign wire633 = ( wire19400 ) | ( wire19401 ) | ( n_n3  &  n_n15 ) ;
 assign wire20804 = ( n_n3406 ) | ( wire633 ) | ( wire20802 ) ;
 assign n_n3362 = ( n_n3374 ) | ( wire20798 ) | ( wire20804 ) | ( _37910 ) ;
 assign wire4391 = ( n_n57  &  wire85 ) | ( n_n220  &  wire914  &  n_n57 ) ;
 assign wire20403 = ( n_n896 ) | ( n_n2986 ) | ( wire20401 ) ;
 assign n_n2817 = ( wire4472 ) | ( wire20397 ) | ( wire20400 ) | ( wire20403 ) ;
 assign wire4470 = ( n_n4  &  wire51 ) | ( n_n4  &  n_n43 ) | ( n_n4  &  wire59 ) ;
 assign wire533 = ( wire4470 ) | ( n_n4  &  wire19578 ) | ( n_n4  &  n_n92 ) ;
 assign wire20412 = ( wire876 ) | ( wire533 ) | ( wire20408 ) | ( wire20409 ) ;
 assign wire20484 = ( _37350 ) | ( _37351 ) ;
 assign n_n2804 = ( wire20542 ) | ( wire20540 ) | ( _37406 ) | ( _37407 ) ;
 assign wire20553 = ( wire20495 ) | ( _37422 ) | ( _37429 ) ;
 assign wire4319 = ( _4044 ) | ( _4045 ) | ( _4046 ) ;
 assign wire3292 = ( n_n6  &  wire80 ) | ( n_n6  &  n_n30 ) | ( n_n6  &  n_n101 ) ;
 assign wire21574 = ( n_n5  &  n_n171 ) | ( n_n6  &  wire69 ) ;
 assign n_n2140 = ( wire3292 ) | ( wire21574 ) | ( n_n5  &  wire67 ) ;
 assign wire3370 = ( n_n3  &  wire79 ) | ( n_n279  &  wire905  &  n_n3 ) ;
 assign wire21516 = ( n_n281  &  n_n4  &  wire904 ) | ( n_n281  &  n_n3  &  wire904 ) ;
 assign wire21517 = ( n_n4  &  n_n12 ) | ( n_n3  &  n_n12 ) | ( n_n3  &  wire83 ) ;
 assign n_n2099 = ( wire3370 ) | ( wire21516 ) | ( wire21517 ) ;
 assign wire281 = ( (~ i_14_)  &  i_13_  &  i_12_  &  wire905 ) | ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire905 ) | ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  wire905 ) ;
 assign wire338 = ( i_15_  &  n_n281  &  n_n259 ) | ( i_15_  &  n_n279  &  n_n259 ) | ( (~ i_15_)  &  n_n279  &  n_n259 ) ;
 assign wire858 = ( i_15_  &  n_n281  &  n_n275 ) | ( i_15_  &  n_n279  &  n_n275 ) | ( (~ i_15_)  &  n_n279  &  n_n275 ) ;
 assign wire1413 = ( wire119 ) | ( wire281 ) | ( wire338 ) | ( wire858 ) ;
 assign wire242 = ( i_15_  &  n_n281  &  n_n253 ) | ( i_15_  &  n_n279  &  n_n253 ) | ( (~ i_15_)  &  n_n279  &  n_n253 ) ;
 assign wire1416 = ( wire153 ) | ( wire255 ) | ( wire241 ) | ( wire242 ) ;
 assign n_n2097 = ( n_n100  &  wire330 ) | ( n_n100  &  wire1416 ) | ( n_n94  &  wire1416 ) ;
 assign wire3419 = ( n_n260  &  n_n285  &  n_n263  &  wire330 ) ;
 assign wire21482 = ( wire907  &  n_n279  &  n_n100 ) | ( n_n279  &  wire901  &  n_n100 ) ;
 assign wire21483 = ( n_n100  &  _38625 ) | ( wire907  &  n_n100  &  _36212 ) ;
 assign n_n2180 = ( wire391 ) | ( wire3419 ) | ( wire21482 ) | ( wire21483 ) ;
 assign wire1423 = ( i_8_  &  n_n260  &  n_n285  &  n_n155 ) | ( (~ i_8_)  &  n_n260  &  n_n285  &  n_n155 ) ;
 assign n_n3770 = ( n_n1  &  n_n76 ) | ( n_n2  &  wire56 ) ;
 assign wire21963 = ( i_14_  &  i_13_  &  i_12_  &  wire903 ) | ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire903 ) | ( i_14_  &  i_13_  &  (~ i_12_)  &  wire903 ) | ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  wire903 ) | ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire903 ) ;
 assign wire1424 = ( wire49 ) | ( n_n79 ) | ( wire212 ) | ( wire21963 ) ;
 assign wire22000 = ( n_n4  &  wire68 ) | ( n_n265  &  n_n62 ) ;
 assign wire22007 = ( n_n1370 ) | ( wire22005 ) | ( n_n268  &  wire273 ) ;
 assign wire587 = ( (~ i_7_)  &  i_6_  &  n_n260  &  n_n118 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n260  &  n_n118 ) ;
 assign wire4565 = ( wire113  &  n_n48 ) | ( n_n48  &  wire101 ) ;
 assign wire20275 = ( n_n53  &  _37158 ) | ( wire914  &  n_n53  &  _34565 ) ;
 assign wire3660 = ( _3222 ) | ( _3223 ) | ( n_n3  &  wire78 ) ;
 assign wire3661 = ( _3216 ) | ( _3217 ) | ( _3218 ) ;
 assign wire21236 = ( wire3653 ) | ( wire21233 ) | ( _3206 ) | ( _38268 ) ;
 assign n_n3709 = ( _6069 ) | ( _6070 ) | ( n_n56  &  _35566 ) ;
 assign wire882 = ( n_n53  &  _37160 ) | ( wire901  &  n_n53  &  _35946 ) ;
 assign wire4453 = ( _37323 ) | ( wire75  &  n_n53 ) | ( n_n53  &  _37322 ) ;
 assign wire20429 = ( wire516 ) | ( wire676 ) | ( wire882 ) | ( wire20424 ) ;
 assign wire20430 = ( n_n3791 ) | ( wire20425 ) | ( _4277 ) ;
 assign wire20452 = ( wire20449 ) | ( wire20450 ) | ( _4342 ) | ( _37285 ) ;
 assign wire20469 = ( n_n4381 ) | ( wire4417 ) | ( wire20460 ) | ( wire20461 ) ;
 assign wire20495 = ( n_n4920 ) | ( n_n4912 ) | ( wire20492 ) ;
 assign wire4360 = ( n_n100  &  wire20512 ) | ( n_n100  &  wire20513 ) | ( n_n100  &  wire20514 ) ;
 assign wire20516 = ( n_n3864 ) | ( wire4380 ) | ( _37376 ) ;
 assign wire20541 = ( _4209 ) | ( _4210 ) | ( _5967 ) | ( _5968 ) ;
 assign wire20542 = ( wire20520 ) | ( wire20525 ) | ( _37396 ) | ( _37398 ) ;
 assign wire19408 = ( n_n275  &  _35110 ) | ( n_n275  &  _35111 ) ;
 assign wire693 = ( n_n57  &  wire19408 ) | ( n_n57  &  n_n256  &  wire903 ) ;
 assign wire3277 = ( n_n53  &  n_n270  &  _38883 ) | ( n_n53  &  n_n270  &  _38885 ) ;
 assign wire21590 = ( n_n111  &  n_n48 ) | ( n_n48  &  n_n171 ) | ( n_n48  &  n_n38 ) ;
 assign n_n2154 = ( wire479 ) | ( wire478 ) | ( wire3277 ) | ( wire21590 ) ;
 assign wire3368 = ( n_n3  &  wire62 ) | ( n_n279  &  n_n3  &  wire899 ) ;
 assign wire1450 = ( n_n281  &  wire914 ) | ( n_n281  &  wire908 ) | ( n_n281  &  wire903 ) ;
 assign wire1451 = ( n_n220  &  wire912 ) | ( n_n220  &  wire898 ) ;
 assign wire823 = ( n_n268  &  wire124 ) | ( n_n268  &  wire212 ) ;
 assign wire22087 = ( wire22081 ) | ( wire22082 ) | ( wire22084 ) ;
 assign wire22088 = ( wire2725 ) | ( wire2726 ) | ( wire22083 ) ;
 assign n_n1124 = ( n_n1215 ) | ( wire22087 ) | ( wire22088 ) ;
 assign wire22095 = ( n_n1173 ) | ( n_n1210 ) | ( wire22093 ) ;
 assign n_n1093 = ( n_n1123 ) | ( n_n1124 ) | ( wire22095 ) ;
 assign wire381 = ( n_n94  &  _36808 ) | ( n_n222  &  n_n94  &  _36699 ) ;
 assign wire152 = ( i_13_  &  (~ i_12_) ) | ( i_14_  &  (~ i_13_)  &  (~ i_12_) ) ;
 assign wire21281 = ( wire913  &  n_n220  &  n_n268 ) | ( n_n220  &  n_n268  &  wire903 ) ;
 assign wire21089 = ( wire780 ) | ( wire654 ) | ( wire3791 ) | ( wire21085 ) ;
 assign wire21090 = ( n_n3864 ) | ( n_n2724 ) | ( wire3790 ) ;
 assign wire20573 = ( wire64 ) | ( wire453 ) | ( _37546 ) ;
 assign wire20574 = ( wire85 ) | ( wire19384 ) | ( _37548 ) ;
 assign wire20575 = ( wire89 ) | ( wire86 ) | ( _37550 ) ;
 assign wire20576 = ( wire55 ) | ( wire57 ) | ( _37552 ) ;
 assign wire1463 = ( wire20573 ) | ( wire20574 ) | ( wire20575 ) | ( wire20576 ) ;
 assign n_n2808 = ( n_n4  &  wire245 ) | ( n_n4  &  n_n39 ) | ( n_n4  &  wire1463 ) ;
 assign wire20435 = ( wire20434 ) | ( _4357 ) ;
 assign wire4435 = ( n_n6  &  wire40 ) | ( n_n6  &  n_n258  &  wire899 ) ;
 assign wire20437 = ( n_n6  &  wire69 ) | ( n_n6  &  n_n258  &  wire897 ) ;
 assign wire20442 = ( n_n4633 ) | ( n_n4632 ) | ( wire20438 ) ;
 assign wire20583 = ( wire20581 ) | ( _3979 ) | ( _3980 ) ;
 assign n_n2806 = ( wire20583 ) | ( _3988 ) | ( _37560 ) | ( _37565 ) ;
 assign wire792 = ( n_n4  &  n_n171 ) | ( n_n4  &  wire56 ) | ( n_n4  &  wire53 ) ;
 assign wire3272 = ( n_n48  &  n_n247  &  _38860 ) | ( n_n48  &  n_n247  &  _38862 ) ;
 assign wire21593 = ( n_n53  &  n_n280 ) | ( n_n53  &  n_n33 ) | ( n_n53  &  n_n35 ) ;
 assign n_n2155 = ( wire376 ) | ( wire464 ) | ( wire3272 ) | ( wire21593 ) ;
 assign wire21596 = ( n_n279  &  wire912 ) | ( n_n279  &  wire901 ) ;
 assign n_n3751 = ( n_n284  &  n_n285  &  n_n271  &  wire212 ) ;
 assign wire380 = ( n_n281  &  n_n94  &  wire897 ) | ( n_n256  &  n_n94  &  wire897 ) ;
 assign wire1474 = ( n_n260  &  n_n165  &  n_n208 ) | ( n_n260  &  n_n165  &  n_n273 ) ;
 assign wire20457 = ( n_n3019 ) | ( wire20455 ) | ( _4318 ) ;
 assign wire395 = ( n_n1  &  wire88 ) | ( n_n1  &  n_n29 ) | ( n_n1  &  wire49 ) ;
 assign wire20562 = ( n_n3259 ) | ( n_n3260 ) | ( wire4313 ) ;
 assign wire829 = ( n_n1  &  n_n171 ) | ( n_n1  &  wire56 ) | ( n_n1  &  wire53 ) ;
 assign wire21379 = ( wire913  &  n_n281 ) | ( n_n220  &  wire914 ) ;
 assign wire1485 = ( i_15_  &  n_n279  &  n_n282 ) | ( (~ i_15_)  &  n_n279  &  n_n282 ) | ( (~ i_15_)  &  n_n282  &  n_n225 ) ;
 assign wire21572 = ( wire376 ) | ( wire3296 ) | ( wire3297 ) | ( wire21569 ) ;
 assign wire21551 = ( n_n279  &  wire899 ) | ( n_n279  &  wire897 ) ;
 assign wire1486 = ( wire40 ) | ( n_n74 ) | ( wire21367 ) | ( wire21551 ) ;
 assign wire343 = ( (~ i_15_)  &  n_n228  &  n_n242 ) | ( i_15_  &  n_n242  &  n_n222 ) | ( (~ i_15_)  &  n_n242  &  n_n222 ) ;
 assign wire21930 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire902 ) | ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  wire902 ) ;
 assign wire2019 = ( n_n53  &  wire368 ) | ( n_n53  &  n_n88 ) | ( n_n53  &  wire145 ) ;
 assign wire22710 = ( n_n37  &  n_n48 ) | ( n_n48  &  wire89 ) | ( n_n48  &  n_n104 ) ;
 assign n_n834 = ( wire2019 ) | ( wire22710 ) ;
 assign n_n560 = ( n_n264  &  n_n273  &  n_n285  &  wire123 ) ;
 assign wire5834 = ( n_n223  &  n_n122 ) | ( n_n122  &  wire214 ) | ( n_n122  &  wire19344 ) ;
 assign wire5835 = ( n_n123  &  wire19347 ) | ( n_n123  &  wire19348 ) ;
 assign wire5843 = ( n_n124  &  n_n253 ) | ( n_n124  &  n_n143 ) | ( n_n124  &  wire214 ) ;
 assign wire5844 = ( n_n123  &  wire19342 ) | ( n_n123  &  n_n282  &  wire1074 ) ;
 assign n_n5009 = ( wire5834 ) | ( wire5835 ) | ( wire5843 ) | ( wire5844 ) ;
 assign wire4478 = ( n_n4  &  wire66 ) | ( wire905  &  n_n4  &  n_n222 ) ;
 assign wire716 = ( _38272 ) | ( n_n4  &  wire66 ) | ( n_n4  &  _37480 ) ;
 assign wire4344 = ( _4219 ) | ( _4220 ) | ( _4221 ) ;
 assign wire20532 = ( wire907  &  n_n228  &  n_n100 ) | ( wire907  &  n_n279  &  n_n100 ) ;
 assign wire20533 = ( n_n37  &  n_n100 ) | ( n_n104  &  n_n100 ) | ( n_n100  &  n_n84 ) ;
 assign wire3287 = ( n_n6  &  n_n84 ) | ( n_n6  &  n_n35 ) | ( n_n6  &  wire86 ) ;
 assign wire21579 = ( n_n111  &  n_n6 ) | ( n_n6  &  wire78 ) | ( n_n6  &  n_n38 ) ;
 assign n_n1598 = ( n_n111  &  n_n57 ) | ( n_n56  &  wire85 ) ;
 assign wire704 = ( wire200  &  n_n56 ) | ( wire112  &  n_n56 ) ;
 assign n_n3523 = ( n_n110  &  n_n1 ) | ( n_n2  &  wire82 ) ;
 assign wire21975 = ( i_14_  &  i_13_  &  i_12_  &  wire905 ) | ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire905 ) | ( i_14_  &  i_13_  &  (~ i_12_)  &  wire905 ) | ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  wire905 ) | ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire905 ) ;
 assign wire1514 = ( wire73 ) | ( n_n252 ) | ( wire100 ) | ( wire21975 ) ;
 assign n_n1591 = ( n_n57  &  wire69 ) | ( n_n56  &  n_n103 ) ;
 assign wire144 = ( i_15_  &  n_n282  &  n_n256 ) | ( (~ i_15_)  &  n_n282  &  n_n256 ) ;
 assign n_n618 = ( n_n48  &  n_n41 ) | ( n_n53  &  wire144 ) ;
 assign wire1517 = ( i_8_  &  n_n264  &  n_n285  &  n_n155 ) | ( (~ i_8_)  &  n_n264  &  n_n285  &  n_n155 ) ;
 assign wire5550 = ( n_n57  &  wire73 ) | ( n_n228  &  n_n57  &  wire900 ) ;
 assign wire5244 = ( n_n6  &  n_n83 ) | ( n_n6  &  wire89 ) | ( n_n6  &  wire85 ) ;
 assign wire5245 = ( n_n220  &  wire907  &  n_n5 ) ;
 assign wire19865 = ( n_n4864 ) | ( n_n4870 ) | ( wire5099 ) | ( wire19862 ) ;
 assign n_n4773 = ( wire389 ) | ( wire708 ) | ( n_n5  &  wire166 ) ;
 assign n_n4680 = ( n_n57  &  wire76 ) | ( n_n279  &  n_n57  &  wire900 ) ;
 assign wire468 = ( n_n1  &  wire60 ) | ( n_n1  &  n_n204 ) | ( n_n1  &  wire52 ) ;
 assign wire21609 = ( n_n279  &  wire899 ) | ( n_n279  &  wire897 ) ;
 assign wire1528 = ( wire40 ) | ( n_n74 ) | ( wire21367 ) | ( wire21609 ) ;
 assign wire369 = ( i_15_  &  n_n279  &  n_n270 ) | ( (~ i_15_)  &  n_n279  &  n_n270 ) ;
 assign wire1530 = ( i_15_  &  n_n279  &  n_n275 ) | ( (~ i_15_)  &  n_n279  &  n_n275 ) | ( i_15_  &  n_n279  &  n_n259 ) | ( (~ i_15_)  &  n_n279  &  n_n259 ) ;
 assign n_n4489 = ( n_n111  &  n_n130 ) | ( wire48  &  n_n128 ) ;
 assign n_n4677 = ( n_n56  &  wire68 ) | ( n_n57  &  n_n42 ) ;
 assign wire371 = ( wire913  &  n_n279 ) | ( wire914  &  n_n279 ) ;
 assign wire1545 = ( wire913  &  n_n279 ) | ( wire914  &  n_n279 ) | ( n_n279  &  wire905 ) ;
 assign wire20192 = ( n_n122  &  n_n109 ) | ( n_n121  &  wire371 ) | ( n_n122  &  wire371 ) ;
 assign wire20117 = ( n_n6  &  n_n54 ) | ( wire72  &  n_n56 ) ;
 assign wire4655 = ( _4811 ) | ( n_n57  &  n_n179 ) | ( n_n57  &  wire57 ) ;
 assign wire20199 = ( n_n4671 ) | ( wire4656 ) | ( n_n56  &  n_n95 ) ;
 assign wire20200 = ( n_n4675 ) | ( n_n4674 ) | ( n_n4676 ) | ( n_n1598 ) ;
 assign wire20209 = ( wire20206 ) | ( _36887 ) ;
 assign wire1552 = ( wire190 ) | ( wire124 ) | ( wire212 ) | ( wire119 ) ;
 assign wire19485 = ( n_n6  &  wire153 ) | ( n_n6  &  wire166 ) | ( n_n6  &  wire180 ) ;
 assign n_n3638 = ( n_n3417 ) | ( wire19387 ) | ( _6235 ) | ( _6236 ) ;
 assign wire19398 = ( n_n3751 ) | ( _6205 ) | ( _35468 ) | ( _35472 ) ;
 assign n_n3624 = ( n_n3638 ) | ( wire19398 ) | ( wire19393 ) | ( _35464 ) ;
 assign wire19405 = ( wire349 ) | ( wire19400 ) | ( wire19401 ) | ( wire5743 ) ;
 assign wire5734 = ( n_n4  &  wire61 ) | ( n_n279  &  n_n4  &  wire908 ) ;
 assign wire19413 = ( n_n3731 ) | ( n_n3736 ) | ( wire792 ) ;
 assign n_n3550 = ( n_n257  &  n_n227 ) | ( n_n240  &  n_n227 ) | ( n_n240  &  n_n207 ) ;
 assign wire20862 = ( n_n3525 ) | ( n_n3524 ) | ( _3692 ) ;
 assign n_n3380 = ( n_n3523 ) | ( wire20862 ) | ( _3695 ) | ( _37852 ) ;
 assign wire5569 = ( n_n53  &  n_n93 ) | ( n_n53  &  wire81 ) | ( n_n53  &  wire76 ) ;
 assign wire20836 = ( n_n2440 ) | ( wire20831 ) | ( wire20832 ) | ( wire20833 ) ;
 assign n_n3417 = ( wire455 ) | ( _6237 ) | ( _6238 ) ;
 assign wire4071 = ( n_n1  &  wire225 ) | ( n_n1  &  wire130 ) ;
 assign wire4073 = ( _3597 ) | ( _3598 ) ;
 assign wire20809 = ( n_n2  &  n_n226 ) | ( n_n268  &  wire247 ) ;
 assign wire5725 = ( n_n2  &  wire88 ) | ( n_n2  &  n_n29 ) | ( n_n2  &  wire49 ) ;
 assign wire5726 = ( n_n1  &  n_n22 ) | ( n_n1  &  n_n73 ) | ( n_n1  &  wire19408 ) ;
 assign n_n2598 = ( n_n3768 ) | ( wire829 ) | ( n_n2  &  n_n22 ) ;
 assign n_n2579 = ( n_n3768 ) | ( wire829 ) | ( _6301 ) | ( _36238 ) ;
 assign wire2975 = ( wire64  &  n_n53 ) | ( wire907  &  n_n222  &  n_n53 ) ;
 assign wire2976 = ( n_n282  &  _39005  &  _39122 ) | ( n_n282  &  _39006  &  _39122 ) ;
 assign wire21827 = ( n_n281  &  wire901  &  n_n53 ) | ( n_n222  &  wire901  &  n_n53 ) ;
 assign wire21828 = ( n_n53  &  n_n32 ) | ( n_n48  &  n_n88 ) ;
 assign n_n1781 = ( wire2975 ) | ( wire2976 ) | ( wire21827 ) | ( wire21828 ) ;
 assign n_n785 = ( n_n896 ) | ( wire712 ) | ( n_n4  &  wire139 ) ;
 assign wire22546 = ( n_n10  &  n_n100 ) | ( n_n94  &  n_n41 ) ;
 assign wire22547 = ( n_n100  &  n_n81 ) | ( n_n94  &  n_n86 ) ;
 assign wire22548 = ( wire57  &  n_n94 ) | ( n_n258  &  wire903  &  n_n94 ) ;
 assign n_n413 = ( wire434 ) | ( wire22546 ) | ( wire22547 ) | ( wire22548 ) ;
 assign wire471 = ( n_n279  &  wire903  &  n_n94 ) | ( n_n222  &  wire903  &  n_n94 ) ;
 assign wire22556 = ( wire22551 ) | ( wire22552 ) ;
 assign wire22557 = ( wire743 ) | ( wire2205 ) | ( n_n257  &  n_n227 ) ;
 assign wire22558 = ( wire658 ) | ( wire642 ) | ( wire471 ) | ( wire2206 ) ;
 assign n_n359 = ( n_n413 ) | ( wire22556 ) | ( wire22557 ) | ( wire22558 ) ;
 assign wire5238 = ( n_n6  &  n_n32 ) | ( n_n6  &  n_n81 ) | ( n_n6  &  wire86 ) ;
 assign wire5239 = ( n_n247  &  _36001  &  _36215 ) | ( n_n247  &  _36002  &  _36215 ) ;
 assign wire19900 = ( n_n4858 ) | ( wire5047 ) | ( _5153 ) ;
 assign wire1575 = ( wire913  &  n_n279 ) | ( wire914  &  n_n279 ) | ( n_n279  &  wire905 ) ;
 assign n_n4685 = ( n_n57  &  n_n95 ) | ( n_n56  &  wire81 ) ;
 assign wire19387 = ( wire5775 ) | ( wire19383 ) | ( n_n268  &  n_n59 ) ;
 assign wire19495 = ( n_n3791 ) | ( wire5606 ) | ( n_n9  &  n_n53 ) ;
 assign wire19489 = ( n_n3827 ) | ( wire771 ) | ( n_n3579 ) ;
 assign wire19490 = ( wire770 ) | ( wire5617 ) | ( wire5625 ) | ( wire5626 ) ;
 assign wire5720 = ( n_n2  &  wire73 ) | ( n_n2  &  n_n65 ) | ( n_n2  &  n_n12 ) ;
 assign wire20865 = ( wire4005 ) | ( wire5709 ) | ( n_n1  &  n_n12 ) ;
 assign wire20866 = ( n_n3519 ) | ( n_n3520 ) | ( wire4004 ) ;
 assign n_n3379 = ( wire5720 ) | ( wire20865 ) | ( wire20866 ) | ( _35346 ) ;
 assign wire4042 = ( n_n6  &  wire60 ) | ( n_n6  &  n_n204 ) | ( n_n6  &  wire1619 ) ;
 assign n_n3393 = ( n_n1536 ) | ( n_n3581 ) | ( wire20847 ) | ( _37833 ) ;
 assign wire20501 = ( _4260 ) | ( n_n57  &  n_n93 ) | ( n_n57  &  wire76 ) ;
 assign wire20502 = ( n_n4686 ) | ( wire4373 ) | ( wire20499 ) ;
 assign n_n2633 = ( n_n1  &  n_n108 ) | ( n_n2  &  wire60 ) ;
 assign wire5711 = ( n_n1  &  wire80 ) | ( n_n1  &  wire908  &  n_n256 ) ;
 assign wire812 = ( n_n3772 ) | ( n_n3770 ) | ( wire5711 ) ;
 assign wire19770 = ( wire395 ) | ( wire5215 ) | ( n_n111  &  n_n2 ) ;
 assign n_n2580 = ( wire812 ) | ( wire19770 ) | ( _6298 ) | ( _35368 ) ;
 assign wire1593 = ( wire913  &  n_n281 ) | ( n_n281  &  wire914 ) ;
 assign wire21668 = ( n_n267  &  _38972 ) | ( n_n267  &  _38973 ) ;
 assign wire21834 = ( i_15_  &  n_n222  &  n_n247 ) | ( i_15_  &  n_n222  &  n_n267 ) ;
 assign wire1594 = ( n_n44 ) | ( wire270 ) | ( wire21668 ) | ( wire21834 ) ;
 assign n_n1713 = ( n_n1785 ) | ( _2220 ) | ( _2223 ) | ( _2224 ) ;
 assign wire195 = ( n_n242  &  _39010 ) | ( n_n242  &  _39011 ) ;
 assign wire21748 = ( n_n220  &  wire912 ) | ( n_n220  &  wire898 ) ;
 assign wire21749 = ( n_n220  &  wire902 ) | ( n_n220  &  wire901 ) ;
 assign wire1597 = ( n_n17 ) | ( wire195 ) | ( wire21748 ) | ( wire21749 ) ;
 assign wire375 = ( n_n259  &  _38957 ) | ( n_n259  &  _38958 ) ;
 assign wire240 = ( i_15_  &  n_n225  &  n_n259 ) | ( i_15_  &  n_n222  &  n_n259 ) | ( (~ i_15_)  &  n_n222  &  n_n259 ) ;
 assign wire21746 = ( n_n220  &  wire898 ) | ( n_n220  &  wire901 ) ;
 assign wire1596 = ( n_n20 ) | ( wire375 ) | ( wire240 ) | ( wire21746 ) ;
 assign wire857 = ( i_15_  &  n_n242  &  n_n225 ) | ( i_15_  &  n_n242  &  n_n222 ) | ( (~ i_15_)  &  n_n242  &  n_n222 ) ;
 assign wire1599 = ( n_n20 ) | ( wire375 ) | ( wire240 ) | ( wire857 ) ;
 assign wire494 = ( i_15_  &  n_n222  &  n_n267 ) | ( (~ i_15_)  &  n_n222  &  n_n267 ) ;
 assign wire1600 = ( i_15_  &  n_n222  &  n_n253 ) | ( (~ i_15_)  &  n_n222  &  n_n253 ) | ( i_15_  &  n_n222  &  n_n267 ) | ( (~ i_15_)  &  n_n222  &  n_n267 ) ;
 assign wire21766 = ( wire21761 ) | ( wire21764 ) | ( n_n56  &  wire180 ) ;
 assign wire21767 = ( wire3045 ) | ( wire21741 ) | ( wire21742 ) | ( wire21762 ) ;
 assign wire21769 = ( wire21752 ) | ( wire21753 ) | ( wire21759 ) | ( wire21760 ) ;
 assign n_n1691 = ( wire21766 ) | ( wire21767 ) | ( wire21769 ) ;
 assign wire862 = ( n_n4  &  n_n54 ) | ( n_n4  &  n_n99 ) | ( n_n4  &  wire96 ) ;
 assign wire895 = ( n_n268  &  wire310 ) | ( n_n268  &  wire22769 ) ;
 assign wire855 = ( n_n268  &  wire55 ) | ( n_n268  &  wire368 ) | ( n_n268  &  n_n39 ) ;
 assign wire856 = ( n_n265  &  wire89 ) | ( n_n265  &  wire22772 ) ;
 assign wire1606 = ( n_n228  &  wire912 ) | ( n_n228  &  wire902 ) | ( n_n228  &  wire901 ) ;
 assign wire22778 = ( n_n1  &  n_n65 ) | ( n_n2  &  n_n65 ) | ( n_n1  &  n_n15 ) ;
 assign n_n750 = ( n_n790 ) | ( wire22780 ) | ( _40657 ) | ( _40658 ) ;
 assign wire22561 = ( n_n4  &  n_n257 ) | ( n_n53  &  n_n197 ) ;
 assign wire22562 = ( n_n3  &  n_n252 ) | ( n_n53  &  n_n26 ) ;
 assign wire22565 = ( n_n53  &  n_n31 ) | ( n_n53  &  wire140 ) | ( n_n53  &  n_n78 ) ;
 assign wire20134 = ( n_n1497 ) | ( _4681 ) ;
 assign wire20119 = ( n_n4892 ) | ( n_n4895 ) | ( wire5035 ) | ( wire5036 ) ;
 assign wire20122 = ( n_n4898 ) | ( wire5013 ) | ( wire5014 ) ;
 assign wire5439 = ( n_n165  &  n_n283  &  wire19294  &  wire923 ) ;
 assign wire609 = ( wire5439 ) | ( n_n220  &  wire914  &  n_n128 ) ;
 assign wire5721 = ( n_n253  &  _35042  &  _36253 ) | ( n_n253  &  _35043  &  _36253 ) ;
 assign wire19784 = ( n_n3525 ) | ( n_n3519 ) | ( n_n3520 ) | ( n_n3524 ) ;
 assign wire19778 = ( _5457 ) | ( _5458 ) | ( _36250 ) ;
 assign wire19787 = ( n_n2633 ) | ( _5425 ) | ( _5426 ) ;
 assign n_n2578 = ( wire19787 ) | ( _5435 ) | ( _36267 ) | ( _36273 ) ;
 assign wire19793 = ( wire19791 ) | ( _5422 ) | ( _36277 ) | ( _36282 ) ;
 assign n_n2572 = ( wire19784 ) | ( n_n2578 ) | ( wire19793 ) | ( _36264 ) ;
 assign wire19798 = ( n_n3781 ) | ( n_n3778 ) | ( _5405 ) ;
 assign wire19802 = ( n_n111  &  n_n1 ) | ( n_n1  &  wire453 ) | ( n_n1  &  n_n38 ) ;
 assign n_n2582 = ( wire806 ) | ( wire19802 ) | ( _36297 ) ;
 assign wire1627 = ( wire268 ) | ( n_n62 ) | ( wire277 ) | ( wire101 ) ;
 assign n_n1773 = ( wire679 ) | ( wire3018 ) | ( wire3019 ) | ( wire21786 ) ;
 assign wire21783 = ( wire21780 ) | ( n_n48  &  wire102 ) ;
 assign wire21784 = ( wire629 ) | ( wire21781 ) | ( n_n53  &  n_n34 ) ;
 assign wire21792 = ( wire631 ) | ( wire3012 ) | ( wire21790 ) ;
 assign n_n1709 = ( n_n1773 ) | ( wire21783 ) | ( wire21784 ) | ( wire21792 ) ;
 assign wire21794 = ( i_15_  &  n_n222  &  n_n247 ) | ( i_15_  &  n_n222  &  n_n267 ) ;
 assign wire1630 = ( n_n44 ) | ( wire270 ) | ( wire21668 ) | ( wire21794 ) ;
 assign wire21799 = ( wire3043 ) | ( n_n6  &  wire1329 ) | ( n_n6  &  wire1630 ) ;
 assign n_n1688 = ( n_n1709 ) | ( _1966 ) | ( _1967 ) | ( _39307 ) ;
 assign wire3000 = ( n_n6  &  n_n203 ) | ( n_n6  &  wire21805 ) | ( n_n6  &  wire21807 ) ;
 assign wire21808 = ( wire3003 ) | ( wire3004 ) | ( n_n6  &  n_n108 ) ;
 assign n_n1706 = ( wire3000 ) | ( wire21808 ) | ( _1952 ) | ( _39309 ) ;
 assign wire21813 = ( n_n5  &  n_n8 ) | ( n_n6  &  n_n58 ) ;
 assign wire21814 = ( n_n80  &  n_n227 ) | ( n_n144  &  wire1776 ) ;
 assign wire21817 = ( wire21811 ) | ( wire21815 ) | ( n_n5  &  wire1291 ) ;
 assign wire21825 = ( _1903 ) | ( _39337 ) | ( _39341 ) ;
 assign n_n1687 = ( n_n1706 ) | ( wire21817 ) | ( wire21825 ) | ( _39332 ) ;
 assign wire2960 = ( n_n48  &  n_n29 ) | ( n_n48  &  n_n80 ) | ( n_n48  &  wire61 ) ;
 assign wire2961 = ( n_n53  &  n_n24 ) | ( n_n53  &  wire104 ) | ( n_n53  &  wire228 ) ;
 assign wire21847 = ( wire2952 ) | ( wire21844 ) | ( wire21845 ) ;
 assign n_n1711 = ( wire21842 ) | ( wire21847 ) | ( _2215 ) | ( _39118 ) ;
 assign wire21855 = ( n_n1781 ) | ( wire2973 ) | ( wire2974 ) | ( wire21853 ) ;
 assign wire22675 = ( n_n228  &  wire898 ) | ( n_n258  &  wire899 ) ;
 assign wire22676 = ( i_15_  &  n_n242  &  n_n225 ) | ( (~ i_15_)  &  n_n242  &  n_n225 ) | ( i_15_  &  n_n225  &  n_n259 ) | ( (~ i_15_)  &  n_n225  &  n_n259 ) ;
 assign wire1637 = ( n_n221 ) | ( wire469 ) | ( wire22675 ) | ( wire22676 ) ;
 assign wire22678 = ( wire647 ) | ( wire2067 ) | ( n_n5  &  n_n197 ) ;
 assign wire275 = ( (~ i_14_)  &  i_15_  &  n_n270  &  n_n254 ) | ( i_14_  &  (~ i_15_)  &  n_n270  &  n_n254 ) | ( (~ i_14_)  &  (~ i_15_)  &  n_n270  &  n_n254 ) ;
 assign wire262 = ( (~ i_14_)  &  i_15_  &  n_n275  &  n_n254 ) | ( i_14_  &  (~ i_15_)  &  n_n275  &  n_n254 ) | ( (~ i_14_)  &  (~ i_15_)  &  n_n275  &  n_n254 ) ;
 assign wire887 = ( n_n227  &  wire198 ) | ( n_n207  &  wire262 ) ;
 assign wire1640 = ( n_n228  &  wire912 ) | ( n_n228  &  wire902 ) ;
 assign wire1639 = ( n_n228  &  wire912 ) | ( n_n228  &  wire898 ) | ( n_n228  &  wire897 ) ;
 assign wire1638 = ( n_n228  &  wire901 ) | ( n_n228  &  wire900 ) ;
 assign wire145 = ( i_15_  &  n_n225  &  n_n247 ) | ( (~ i_15_)  &  n_n225  &  n_n247 ) ;
 assign wire22687 = ( i_15_  &  n_n258  &  n_n275 ) | ( i_15_  &  n_n225  &  n_n275 ) | ( (~ i_15_)  &  n_n225  &  n_n275 ) ;
 assign wire1641 = ( wire19457 ) | ( n_n25 ) | ( wire145 ) | ( wire22687 ) ;
 assign wire22685 = ( wire887 ) | ( wire22683 ) ;
 assign wire22686 = ( wire2059 ) | ( wire22680 ) | ( wire22681 ) | ( wire22684 ) ;
 assign wire22693 = ( n_n4636 ) | ( wire487 ) | ( wire22689 ) | ( wire22692 ) ;
 assign wire1649 = ( n_n258  &  wire906 ) | ( n_n258  &  wire904 ) ;
 assign wire1647 = ( wire914  &  n_n258 ) | ( n_n258  &  wire906 ) | ( n_n258  &  wire904 ) ;
 assign wire19931 = ( wire760 ) | ( wire19928 ) | ( n_n57  &  wire198 ) ;
 assign wire19946 = ( wire763 ) | ( wire4974 ) | ( wire19943 ) | ( wire19944 ) ;
 assign wire19959 = ( wire19958 ) | ( _5230 ) | ( _5231 ) ;
 assign wire19953 = ( n_n4970 ) | ( n_n4967 ) | ( _36428 ) ;
 assign wire19967 = ( wire19965 ) | ( _36442 ) | ( _36443 ) | ( _36448 ) ;
 assign wire672 = ( wire273  &  n_n57 ) | ( n_n57  &  wire157 ) ;
 assign n_n3803 = ( n_n5  &  wire199 ) | ( n_n6  &  n_n7 ) ;
 assign wire20141 = ( n_n4635 ) | ( wire20137 ) | ( n_n6  &  wire78 ) ;
 assign wire20142 = ( n_n4633 ) | ( n_n4636 ) | ( n_n4632 ) | ( wire4727 ) ;
 assign wire20224 = ( n_n4920 ) | ( n_n4922 ) | ( n_n4921 ) ;
 assign n_n4551 = ( wire705 ) | ( wire721 ) | ( wire20224 ) | ( _4775 ) ;
 assign wire19537 = ( n_n56  &  wire49 ) | ( n_n57  &  n_n22 ) ;
 assign n_n3708 = ( n_n4926 ) | ( wire693 ) | ( wire19537 ) ;
 assign wire20228 = ( n_n4907 ) | ( wire636 ) | ( n_n4924 ) | ( wire5544 ) ;
 assign wire20232 = ( n_n4259 ) | ( wire465 ) | ( n_n3708 ) | ( wire20227 ) ;
 assign wire20872 = ( _3674 ) | ( _3675 ) | ( _37862 ) ;
 assign wire3989 = ( wire123  &  n_n227 ) | ( n_n227  &  wire20875 ) ;
 assign wire20881 = ( n_n4806 ) | ( n_n3550 ) | ( wire3988 ) | ( wire20876 ) ;
 assign wire3985 = ( n_n4  &  wire123 ) | ( n_n4  &  wire100 ) ;
 assign wire20882 = ( n_n4  &  n_n197 ) | ( n_n4  &  n_n223 ) | ( n_n4  &  n_n221 ) ;
 assign wire20888 = ( wire455 ) | ( wire388 ) | ( wire381 ) | ( wire20883 ) ;
 assign wire20889 = ( wire333 ) | ( n_n6820 ) | ( wire3975 ) | ( wire3976 ) ;
 assign n_n3385 = ( wire3985 ) | ( wire20882 ) | ( wire20888 ) | ( wire20889 ) ;
 assign wire20508 = ( n_n3604 ) | ( wire740 ) | ( wire20506 ) ;
 assign wire227 = ( i_14_  &  (~ i_13_)  &  i_12_  &  wire899 ) | ( i_14_  &  i_13_  &  (~ i_12_)  &  wire899 ) | ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire899 ) ;
 assign wire1662 = ( wire123 ) | ( wire100 ) | ( wire281 ) | ( wire227 ) ;
 assign wire1661 = ( n_n112 ) | ( wire165 ) | ( wire52 ) | ( wire167 ) ;
 assign wire1664 = ( wire190 ) | ( wire124 ) | ( wire212 ) | ( wire119 ) ;
 assign wire20068 = ( wire20066 ) | ( n_n94  &  wire140 ) | ( n_n94  &  wire1661 ) ;
 assign wire20073 = ( wire20072 ) | ( n_n100  &  wire1664 ) ;
 assign wire1668 = ( n_n220  &  wire912 ) | ( n_n220  &  wire900 ) | ( n_n220  &  wire897 ) ;
 assign wire21888 = ( n_n220  &  n_n4  &  wire902 ) | ( n_n220  &  n_n4  &  wire900 ) ;
 assign wire21889 = ( n_n4  &  n_n147 ) | ( n_n3  &  n_n14 ) ;
 assign wire426 = ( i_15_  &  n_n222  &  n_n275 ) | ( (~ i_15_)  &  n_n222  &  n_n275 ) ;
 assign wire134 = ( i_15_  &  n_n225  &  n_n253 ) | ( (~ i_15_)  &  n_n225  &  n_n253 ) ;
 assign wire544 = ( n_n53  &  n_n31 ) | ( n_n53  &  n_n80 ) | ( n_n53  &  n_n30 ) ;
 assign wire1669 = ( i_15_  &  n_n225  &  n_n270 ) | ( (~ i_15_)  &  n_n225  &  n_n270 ) | ( i_15_  &  n_n225  &  n_n259 ) | ( (~ i_15_)  &  n_n225  &  n_n259 ) ;
 assign wire22792 = ( wire608 ) | ( wire22786 ) | ( n_n4  &  wire1669 ) ;
 assign wire22793 = ( n_n876 ) | ( wire544 ) | ( wire22787 ) | ( wire22788 ) ;
 assign n_n755 = ( n_n785 ) | ( wire22792 ) | ( wire22793 ) ;
 assign wire22803 = ( _40568 ) | ( n_n94  &  n_n88 ) | ( n_n94  &  _36682 ) ;
 assign wire22804 = ( wire697 ) | ( wire22801 ) | ( n_n100  &  n_n33 ) ;
 assign wire22809 = ( n_n884 ) | ( wire564 ) | ( wire22805 ) | ( wire22806 ) ;
 assign n_n756 = ( n_n809 ) | ( wire22803 ) | ( wire22804 ) | ( wire22809 ) ;
 assign wire22814 = ( wire22785 ) | ( _399 ) | ( _40604 ) ;
 assign wire403 = ( wire914  &  n_n258 ) | ( n_n258  &  wire903 ) ;
 assign wire1673 = ( wire905  &  n_n258 ) | ( n_n258  &  wire908 ) ;
 assign wire22451 = ( wire407 ) | ( wire457 ) | ( n_n56  &  n_n257 ) ;
 assign wire1678 = ( wire907  &  n_n258 ) | ( wire905  &  n_n258 ) | ( n_n258  &  wire908 ) ;
 assign wire1677 = ( wire914  &  n_n258 ) | ( n_n258  &  wire908 ) ;
 assign wire1676 = ( wire913  &  n_n258 ) | ( n_n258  &  wire903 ) ;
 assign wire292 = ( (~ i_15_)  &  n_n242  &  n_n279 ) | ( i_15_  &  n_n242  &  n_n256 ) | ( (~ i_15_)  &  n_n242  &  n_n256 ) ;
 assign wire1682 = ( wire913  &  n_n258 ) | ( wire914  &  n_n258 ) | ( n_n258  &  wire908 ) ;
 assign wire1680 = ( wire905  &  n_n258 ) | ( n_n258  &  wire908 ) ;
 assign wire1679 = ( wire907  &  n_n258 ) | ( n_n258  &  wire903 ) ;
 assign wire1687 = ( n_n229  &  n_n165  &  n_n284 ) | ( n_n165  &  n_n284  &  n_n283 ) ;
 assign wire5758 = ( n_n4  &  wire19384 ) | ( n_n281  &  n_n4  &  wire900 ) ;
 assign wire19393 = ( wire557 ) | ( wire374 ) | ( wire5754 ) ;
 assign wire20897 = ( n_n257  &  n_n53 ) | ( n_n1  &  wire68 ) ;
 assign wire20904 = ( wire634 ) | ( wire20898 ) | ( wire20900 ) ;
 assign wire20905 = ( n_n2272 ) | ( n_n952 ) | ( n_n560 ) | ( wire20899 ) ;
 assign n_n3383 = ( wire20897 ) | ( wire20904 ) | ( wire20905 ) | ( _3589 ) ;
 assign wire1696 = ( i_15_  &  n_n242  &  n_n222 ) | ( (~ i_15_)  &  n_n242  &  n_n222 ) | ( i_15_  &  n_n222  &  n_n275 ) | ( (~ i_15_)  &  n_n222  &  n_n275 ) ;
 assign wire21652 = ( n_n268  &  n_n22 ) | ( n_n2  &  n_n144 ) ;
 assign wire379 = ( i_15_  &  n_n222  &  n_n270 ) | ( (~ i_15_)  &  n_n222  &  n_n270 ) ;
 assign wire2011 = ( _560 ) | ( _561 ) ;
 assign wire22714 = ( wire2012 ) | ( wire22712 ) | ( n_n54  &  n_n48 ) ;
 assign wire22717 = ( wire22700 ) | ( wire22701 ) | ( wire22708 ) | ( wire22709 ) ;
 assign wire22744 = ( n_n819 ) | ( wire22742 ) | ( _455 ) | ( _40538 ) ;
 assign wire22763 = ( _379 ) | ( _380 ) | ( _382 ) | ( _40607 ) ;
 assign wire22822 = ( n_n750 ) | ( wire22820 ) | ( _40648 ) | ( _40649 ) ;
 assign wire1703 = ( wire913  &  n_n220 ) | ( n_n220  &  wire914 ) | ( n_n220  &  wire905 ) ;
 assign wire1707 = ( n_n281  &  wire911 ) | ( n_n281  &  wire912 ) | ( n_n281  &  wire899 ) ;
 assign wire1706 = ( n_n281  &  wire911 ) | ( n_n281  &  wire912 ) | ( n_n281  &  wire899 ) ;
 assign wire5671 = ( wire120  &  n_n207 ) | ( wire19457  &  n_n207 ) | ( n_n207  &  n_n25 ) ;
 assign wire19458 = ( n_n31  &  n_n227 ) | ( n_n103  &  n_n207 ) ;
 assign n_n3686 = ( wire5671 ) | ( wire19458 ) | ( n_n5  &  wire208 ) ;
 assign wire1717 = ( wire911  &  n_n228 ) | ( n_n228  &  wire897 ) ;
 assign wire236 = ( i_15_  &  n_n225  &  n_n270 ) | ( i_15_  &  n_n222  &  n_n270 ) | ( (~ i_15_)  &  n_n222  &  n_n270 ) ;
 assign wire74 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire897 ) | ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  wire897 ) ;
 assign wire424 = ( i_15_  &  n_n225  &  n_n275 ) | ( i_15_  &  n_n222  &  n_n275 ) | ( (~ i_15_)  &  n_n222  &  n_n275 ) ;
 assign wire1730 = ( wire74 ) | ( wire424 ) | ( n_n220  &  wire903 ) ;
 assign wire1733 = ( wire124 ) | ( n_n258  &  wire897 ) ;
 assign wire1737 = ( wire905  &  n_n258 ) | ( n_n258  &  wire908 ) | ( n_n258  &  wire903 ) ;
 assign wire22403 = ( n_n246  &  n_n48 ) | ( n_n61  &  n_n53 ) ;
 assign wire22404 = ( wire905  &  n_n258  &  n_n53 ) | ( n_n258  &  n_n53  &  wire903 ) ;
 assign wire1740 = ( i_5_  &  (~ i_3_)  &  i_4_  &  n_n118 ) | ( (~ i_5_)  &  (~ i_3_)  &  i_4_  &  n_n118 ) | ( i_5_  &  (~ i_3_)  &  (~ i_4_)  &  n_n118 ) | ( (~ i_5_)  &  (~ i_3_)  &  (~ i_4_)  &  n_n118 ) ;
 assign wire19465 = ( wire455 ) | ( wire374 ) | ( wire19461 ) ;
 assign wire19466 = ( wire799 ) | ( wire471 ) | ( wire19460 ) ;
 assign wire19467 = ( wire747 ) | ( wire5660 ) | ( wire5661 ) ;
 assign wire19523 = ( wire473 ) | ( wire19519 ) | ( wire19520 ) | ( wire19522 ) ;
 assign wire1747 = ( wire140 ) | ( wire165 ) | ( wire167 ) | ( wire198 ) ;
 assign wire1753 = ( n_n228  &  wire902 ) | ( n_n228  &  wire898 ) | ( n_n228  &  wire901 ) ;
 assign wire1752 = ( n_n228  &  wire912 ) | ( n_n228  &  wire898 ) | ( n_n228  &  wire901 ) ;
 assign wire1755 = ( (~ i_15_)  &  n_n279  &  n_n253 ) | ( i_15_  &  n_n256  &  n_n253 ) | ( (~ i_15_)  &  n_n256  &  n_n253 ) ;
 assign wire20075 = ( n_n100  &  n_n81 ) | ( n_n94  &  n_n39 ) ;
 assign wire20076 = ( wire57  &  n_n94 ) | ( n_n100  &  n_n33 ) ;
 assign n_n2671 = ( wire548 ) | ( wire434 ) | ( wire20075 ) | ( wire20076 ) ;
 assign wire20094 = ( wire4800 ) | ( _4943 ) | ( _4944 ) ;
 assign n_n2673 = ( n_n3598 ) | ( wire380 ) | ( wire471 ) | ( wire20096 ) ;
 assign wire20104 = ( wire381 ) | ( wire20099 ) | ( wire20101 ) ;
 assign n_n2659 = ( n_n2673 ) | ( wire20104 ) | ( _36813 ) ;
 assign wire2994 = ( n_n6  &  wire195 ) | ( n_n220  &  n_n6  &  wire898 ) ;
 assign wire3018 = ( n_n53  &  wire21785 ) | ( wire907  &  n_n222  &  n_n53 ) ;
 assign wire3019 = ( n_n220  &  wire911  &  wire185 ) ;
 assign wire21786 = ( n_n37  &  n_n53 ) | ( n_n48  &  n_n144 ) ;
 assign wire1773 = ( n_n220  &  wire902 ) | ( n_n220  &  wire901 ) | ( n_n220  &  wire899 ) ;
 assign wire1772 = ( n_n220  &  wire912 ) | ( n_n220  &  wire902 ) ;
 assign wire1771 = ( n_n220  &  wire911 ) | ( n_n220  &  wire897 ) ;
 assign wire1776 = ( i_8_  &  n_n272  &  n_n285  &  n_n230 ) | ( (~ i_8_)  &  n_n272  &  n_n285  &  n_n230 ) ;
 assign wire1777 = ( n_n228  &  wire912 ) | ( n_n228  &  wire902 ) | ( n_n228  &  wire897 ) ;
 assign wire22829 = ( n_n228  &  n_n4  &  wire902 ) | ( n_n228  &  n_n4  &  wire899 ) ;
 assign wire22830 = ( n_n3  &  n_n226 ) | ( n_n4  &  n_n59 ) ;
 assign wire20153 = ( n_n4624 ) | ( wire411 ) | ( _4622 ) ;
 assign wire20157 = ( n_n1476 ) | ( _4605 ) ;
 assign wire1786 = ( i_14_  &  i_13_  &  i_12_  &  wire904 ) | ( (~ i_14_)  &  i_13_  &  i_12_  &  wire904 ) | ( i_14_  &  i_13_  &  (~ i_12_)  &  wire904 ) | ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire904 ) ;
 assign wire3578 = ( _2984 ) | ( _2985 ) | ( n_n56  &  wire62 ) ;
 assign wire21675 = ( n_n4  &  n_n64 ) | ( n_n53  &  n_n27 ) ;
 assign wire21676 = ( n_n53  &  n_n76 ) | ( n_n3  &  n_n14 ) ;
 assign wire21677 = ( n_n4  &  n_n144 ) | ( n_n53  &  n_n78 ) ;
 assign wire21678 = ( n_n53  &  n_n29 ) | ( n_n53  &  n_n80 ) | ( n_n53  &  n_n28 ) ;
 assign wire622 = ( n_n4  &  _39052 ) | ( n_n4  &  wire899  &  _35752 ) ;
 assign wire1794 = ( (~ i_15_)  &  n_n242  &  n_n222 ) | ( i_15_  &  n_n242  &  n_n256 ) ;
 assign wire22341 = ( i_14_  &  i_13_  &  (~ i_12_)  &  wire906 ) | ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire906 ) ;
 assign wire22572 = ( wire2196 ) | ( wire22570 ) ;
 assign wire22573 = ( wire2200 ) | ( wire22566 ) | ( wire22567 ) | ( wire22571 ) ;
 assign wire22581 = ( wire2463 ) | ( wire22578 ) | ( _848 ) | ( _40234 ) ;
 assign n_n341 = ( n_n359 ) | ( wire22572 ) | ( wire22573 ) | ( wire22581 ) ;
 assign wire1797 = ( wire913  &  n_n279 ) | ( wire914  &  n_n279 ) | ( n_n279  &  wire905 ) ;
 assign wire1796 = ( n_n260  &  n_n229  &  n_n165 ) | ( n_n260  &  n_n165  &  n_n283 ) ;
 assign wire19565 = ( n_n4681 ) | ( n_n4686 ) | ( _6010 ) ;
 assign wire19566 = ( wire863 ) | ( n_n4687 ) | ( wire5506 ) | ( wire5494 ) ;
 assign wire1803 = ( n_n259  &  _39114 ) | ( n_n259  &  _39115 ) ;
 assign wire21864 = ( wire893 ) | ( wire2929 ) ;
 assign wire21865 = ( n_n4477 ) | ( wire21861 ) | ( wire21862 ) ;
 assign wire21874 = ( wire667 ) | ( wire2919 ) | ( wire21872 ) ;
 assign wire21877 = ( n_n1804 ) | ( wire2920 ) | ( wire2927 ) | ( wire2928 ) ;
 assign wire20096 = ( n_n94  &  _36803 ) | ( wire903  &  n_n94  &  _35109 ) ;
 assign wire3576 = ( n_n56  &  n_n7 ) | ( n_n56  &  wire50 ) | ( n_n56  &  n_n59 ) ;
 assign wire3577 = ( n_n57  &  wire208 ) | ( n_n57  &  wire50 ) | ( n_n57  &  n_n59 ) ;
 assign n_n2431 = ( wire3576 ) | ( wire3577 ) | ( _38451 ) ;
 assign wire441 = ( (~ i_15_)  &  n_n279  &  n_n259 ) | ( i_15_  &  n_n256  &  n_n259 ) | ( (~ i_15_)  &  n_n256  &  n_n259 ) ;
 assign wire1814 = ( n_n197 ) | ( wire42 ) | ( wire275 ) | ( wire441 ) ;
 assign wire1813 = ( n_n216 ) | ( wire52 ) | ( wire190 ) | ( wire292 ) ;
 assign wire1825 = ( n_n281  &  wire914 ) | ( n_n281  &  wire907 ) ;
 assign wire20176 = ( n_n3806 ) | ( n_n3803 ) | ( wire20174 ) ;
 assign wire1829 = ( i_5_  &  (~ i_3_)  &  i_4_  &  n_n118 ) | ( (~ i_5_)  &  (~ i_3_)  &  i_4_  &  n_n118 ) | ( i_5_  &  (~ i_3_)  &  (~ i_4_)  &  n_n118 ) ;
 assign wire3720 = ( n_n139  &  n_n135 ) | ( n_n139  &  wire419 ) | ( n_n139  &  wire19604 ) ;
 assign wire21168 = ( wire21164 ) | ( wire21165 ) | ( _3263 ) ;
 assign wire3558 = ( _3021 ) | ( _3022 ) | ( _3023 ) ;
 assign wire21352 = ( wire3562 ) | ( wire3563 ) | ( wire3565 ) | ( wire21337 ) ;
 assign wire362 = ( i_15_  &  n_n282  &  n_n225 ) | ( i_15_  &  n_n282  &  n_n222 ) | ( (~ i_15_)  &  n_n282  &  n_n222 ) ;
 assign wire1835 = ( wire154 ) | ( n_n34 ) | ( wire236 ) | ( wire362 ) ;
 assign wire161 = ( i_15_  &  n_n242  &  n_n225 ) | ( (~ i_15_)  &  n_n242  &  n_n225 ) ;
 assign wire22835 = ( n_n228  &  wire912 ) | ( n_n228  &  wire898 ) ;
 assign wire22833 = ( n_n258  &  wire899 ) | ( n_n228  &  wire900 ) ;
 assign wire1836 = ( n_n221 ) | ( wire469 ) | ( wire128 ) | ( wire22833 ) ;
 assign wire1849 = ( n_n259  &  _39084 ) | ( n_n259  &  _39085 ) ;
 assign wire47 = ( i_14_  &  i_13_  &  (~ i_12_)  &  wire907 ) | ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire907 ) ;
 assign wire19575 = ( i_14_  &  i_13_  &  (~ i_12_)  &  wire904 ) | ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire904 ) ;
 assign wire87 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire912 ) | ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  wire912 ) ;
 assign wire110 = ( i_15_  &  n_n242  &  n_n256 ) | ( (~ i_15_)  &  n_n242  &  n_n256 ) ;
 assign wire288 = ( (~ i_12_) ) | ( i_13_  &  i_12_ ) ;
 assign wire148 = ( (~ i_12_) ) | ( i_13_  &  i_12_ ) | ( (~ i_14_)  &  (~ i_13_)  &  i_12_ ) ;
 assign wire187 = ( i_15_  &  n_n256  &  n_n259 ) | ( (~ i_15_)  &  n_n256  &  n_n259 ) ;
 assign wire196 = ( i_9_  &  (~ i_10_)  &  i_11_ ) | ( i_9_  &  (~ i_10_)  &  i_12_  &  (~ i_11_) ) ;
 assign wire197 = ( i_13_  &  (~ i_12_) ) | ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_) ) ;
 assign wire214 = ( n_n259  &  _34625 ) | ( n_n259  &  _34626 ) ;
 assign wire215 = ( (~ i_9_)  &  i_10_  &  i_11_ ) | ( (~ i_9_)  &  i_10_  &  i_12_  &  (~ i_11_) ) ;
 assign wire220 = ( n_n253  &  _39553 ) | ( n_n253  &  _39554 ) ;
 assign wire230 = ( n_n270  &  _39001 ) | ( n_n270  &  _39002 ) ;
 assign wire231 = ( i_15_  &  n_n256  &  n_n275 ) | ( (~ i_15_)  &  n_n256  &  n_n275 ) ;
 assign wire243 = ( i_15_  &  n_n225  &  n_n267 ) | ( i_15_  &  n_n222  &  n_n267 ) | ( (~ i_15_)  &  n_n222  &  n_n267 ) ;
 assign wire246 = ( n_n267  &  _35531 ) | ( n_n267  &  _35532 ) ;
 assign wire256 = ( n_n267  &  _35529 ) | ( n_n267  &  _35530 ) ;
 assign wire274 = ( (~ i_15_)  &  n_n228  &  n_n259 ) | ( i_15_  &  n_n222  &  n_n259 ) | ( (~ i_15_)  &  n_n222  &  n_n259 ) ;
 assign wire19238 = ( n_n267 ) | ( n_n279  &  wire912 ) ;
 assign wire19253 = ( n_n247  &  _34548 ) | ( n_n247  &  _34549 ) ;
 assign wire287 = ( (~ i_9_)  &  (~ i_10_)  &  i_11_ ) | ( (~ i_9_)  &  (~ i_10_)  &  i_12_  &  (~ i_11_) ) ;
 assign wire291 = ( n_n282  &  _39565 ) | ( n_n282  &  _39566 ) ;
 assign wire304 = ( (~ i_14_)  &  i_15_  &  n_n247  &  n_n254 ) | ( i_14_  &  (~ i_15_)  &  n_n247  &  n_n254 ) | ( (~ i_14_)  &  (~ i_15_)  &  n_n247  &  n_n254 ) ;
 assign wire305 = ( (~ i_14_)  &  i_15_  &  n_n254  &  n_n259 ) | ( i_14_  &  (~ i_15_)  &  n_n254  &  n_n259 ) | ( (~ i_14_)  &  (~ i_15_)  &  n_n254  &  n_n259 ) ;
 assign wire311 = ( (~ i_15_)  &  n_n228  &  n_n253 ) | ( i_15_  &  n_n222  &  n_n253 ) | ( (~ i_15_)  &  n_n222  &  n_n253 ) ;
 assign wire325 = ( i_15_  &  n_n281  &  n_n242 ) | ( i_15_  &  n_n242  &  n_n256 ) | ( (~ i_15_)  &  n_n242  &  n_n256 ) ;
 assign wire328 = ( i_9_  &  i_10_ ) | ( i_9_  &  (~ i_10_)  &  i_11_ ) ;
 assign wire342 = ( i_15_  &  n_n281  &  n_n247 ) | ( i_15_  &  n_n256  &  n_n247 ) | ( (~ i_15_)  &  n_n256  &  n_n247 ) ;
 assign wire345 = ( i_15_  &  n_n281  &  n_n275 ) | ( i_15_  &  n_n256  &  n_n275 ) | ( (~ i_15_)  &  n_n256  &  n_n275 ) ;
 assign wire348 = ( (~ i_14_)  &  i_15_  &  n_n242  &  n_n254 ) | ( i_14_  &  (~ i_15_)  &  n_n242  &  n_n254 ) | ( (~ i_14_)  &  (~ i_15_)  &  n_n242  &  n_n254 ) ;
 assign wire352 = ( i_9_  &  i_10_  &  i_11_ ) | ( i_9_  &  i_10_  &  i_12_  &  (~ i_11_) ) ;
 assign wire361 = ( i_15_  &  n_n225  &  n_n253 ) | ( i_15_  &  n_n222  &  n_n253 ) | ( (~ i_15_)  &  n_n222  &  n_n253 ) ;
 assign wire397 = ( wire215 ) | ( n_n242  &  n_n222 ) ;
 assign wire413 = ( i_15_  &  n_n279  &  n_n259 ) | ( (~ i_15_)  &  n_n279  &  n_n259 ) ;
 assign wire428 = ( i_15_  &  n_n225  &  n_n247 ) | ( i_15_  &  n_n222  &  n_n247 ) | ( (~ i_15_)  &  n_n222  &  n_n247 ) ;
 assign wire431 = ( i_15_  &  n_n281  &  n_n270 ) | ( i_15_  &  n_n256  &  n_n270 ) | ( (~ i_15_)  &  n_n256  &  n_n270 ) ;
 assign wire433 = ( (~ i_15_)  &  n_n228  &  n_n282 ) | ( i_15_  &  n_n282  &  n_n222 ) | ( (~ i_15_)  &  n_n282  &  n_n222 ) ;
 assign wire435 = ( n_n143 ) | ( n_n259  &  _34625 ) | ( n_n259  &  _34626 ) ;
 assign wire437 = ( i_15_  &  n_n281  &  n_n282 ) | ( i_15_  &  n_n282  &  n_n256 ) | ( (~ i_15_)  &  n_n282  &  n_n256 ) ;
 assign wire444 = ( (~ i_15_)  &  n_n279  &  n_n247 ) | ( i_15_  &  n_n256  &  n_n247 ) | ( (~ i_15_)  &  n_n256  &  n_n247 ) ;
 assign wire1874 = ( n_n281  &  wire907 ) | ( n_n228  &  wire912 ) ;
 assign wire1918 = ( _40796 ) | ( n_n270  &  _35064 ) | ( n_n270  &  _35065 ) ;
 assign wire962 = ( i_9_  &  (~ i_10_)  &  i_11_ ) | ( i_9_  &  (~ i_10_)  &  (~ i_11_) ) ;
 assign wire965 = ( (~ i_12_) ) | ( i_13_  &  i_12_ ) | ( (~ i_14_)  &  (~ i_13_)  &  i_12_ ) ;
 assign wire968 = ( (~ i_12_) ) | ( i_13_  &  i_12_ ) | ( (~ i_14_)  &  (~ i_13_)  &  i_12_ ) ;
 assign wire971 = ( (~ i_12_) ) | ( i_13_  &  i_12_ ) | ( (~ i_14_)  &  (~ i_13_)  &  i_12_ ) ;
 assign wire1074 = ( i_13_  &  (~ i_12_) ) | ( i_14_  &  (~ i_13_)  &  (~ i_12_) ) ;
 assign wire1101 = ( n_n281  &  wire914 ) | ( n_n281  &  wire907 ) | ( n_n281  &  wire904 ) ;
 assign wire1135 = ( (~ i_14_)  &  i_13_  &  (~ i_12_) ) | ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_) ) ;
 assign wire1182 = ( (~ i_14_)  &  i_13_  &  (~ i_12_) ) | ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_) ) ;
 assign wire1199 = ( n_n220  &  wire898 ) | ( n_n220  &  wire900 ) ;
 assign wire1225 = ( (~ i_9_)  &  i_10_  &  i_11_ ) | ( (~ i_9_)  &  i_10_  &  (~ i_11_) ) ;
 assign wire1317 = ( i_9_ ) | ( (~ i_9_)  &  i_10_ ) ;
 assign wire1501 = ( (~ i_9_)  &  i_10_  &  (~ i_11_) ) | ( i_9_  &  (~ i_10_)  &  (~ i_11_) ) ;
 assign wire1619 = ( n_n112 ) | ( wire52 ) | ( wire247 ) | ( wire210 ) ;
 assign wire1792 = ( n_n17 ) | ( wire195 ) | ( wire240 ) | ( wire857 ) ;
 assign wire22841 = ( i_15_  &  n_n258  &  n_n247 ) | ( i_15_  &  n_n225  &  n_n247 ) | ( (~ i_15_)  &  n_n225  &  n_n247 ) ;
 assign wire238 = ( n_n3  &  wire368 ) | ( n_n3  &  n_n88 ) | ( n_n3  &  wire22841 ) ;
 assign wire505 = ( n_n228  &  wire169  &  wire901 ) ;
 assign wire22816 = ( i_15_  &  n_n258  &  n_n267 ) | ( i_15_  &  n_n225  &  n_n267 ) | ( (~ i_15_)  &  n_n225  &  n_n267 ) ;
 assign wire529 = ( n_n3  &  n_n46 ) | ( n_n3  &  wire19577 ) | ( n_n3  &  wire22816 ) ;
 assign wire543 = ( n_n1  &  wire254 ) | ( n_n1  &  wire356 ) ;
 assign wire550 = ( n_n260  &  n_n285  &  n_n283  &  wire224 ) ;
 assign wire564 = ( wire914  &  n_n228  &  _40573 ) | ( wire911  &  n_n228  &  _40573 ) ;
 assign wire22795 = ( n_n259  &  _40564 ) | ( n_n259  &  _40565 ) ;
 assign wire608 = ( n_n3  &  n_n253  &  _40544 ) | ( n_n3  &  n_n253  &  _40546 ) ;
 assign wire22772 = ( i_15_  &  n_n282  &  n_n225 ) | ( (~ i_15_)  &  n_n282  &  n_n225 ) ;
 assign wire22769 = ( (~ i_14_)  &  wire914  &  n_n254 ) | ( i_14_  &  wire911  &  n_n254 ) ;
 assign wire1970 = ( _358 ) | ( n_n2  &  wire275 ) | ( n_n2  &  wire348 ) ;
 assign wire22752 = ( wire60 ) | ( n_n204 ) | ( wire227 ) | ( wire348 ) ;
 assign wire1971 = ( n_n1  &  wire262 ) | ( n_n1  &  wire305 ) | ( n_n1  &  wire22752 ) ;
 assign wire22746 = ( i_15_  &  n_n258  &  n_n247 ) | ( i_15_  &  n_n225  &  n_n247 ) | ( (~ i_15_)  &  n_n225  &  n_n247 ) ;
 assign wire1976 = ( n_n4  &  wire368 ) | ( n_n4  &  n_n88 ) | ( n_n4  &  wire22746 ) ;
 assign wire1977 = ( n_n6  &  n_n41 ) | ( n_n6  &  wire139 ) | ( n_n6  &  wire145 ) ;
 assign wire22730 = ( n_n228  &  wire912 ) | ( n_n228  &  wire898 ) ;
 assign wire22719 = ( i_15_  &  n_n258  &  n_n267 ) | ( i_15_  &  n_n225  &  n_n267 ) | ( (~ i_15_)  &  n_n225  &  n_n267 ) ;
 assign wire2012 = ( n_n53  &  n_n46 ) | ( n_n53  &  wire19577 ) | ( n_n53  &  wire139 ) ;
 assign wire2022 = ( n_n264  &  n_n285  &  n_n283  &  wire1343 ) ;
 assign wire2023 = ( n_n225  &  n_n53  &  _40472 ) | ( n_n225  &  n_n53  &  _40474 ) ;
 assign wire2030 = ( n_n48  &  wire120 ) | ( n_n48  &  wire19457 ) | ( n_n48  &  n_n25 ) ;
 assign wire2034 = ( n_n53  &  wire128 ) | ( n_n53  &  n_n203 ) | ( n_n53  &  wire20149 ) ;
 assign wire22696 = ( i_15_  &  n_n242  &  n_n225 ) | ( (~ i_15_)  &  n_n242  &  n_n225 ) | ( i_15_  &  n_n225  &  n_n270 ) | ( (~ i_15_)  &  n_n225  &  n_n270 ) ;
 assign wire2035 = ( n_n48  &  n_n203 ) | ( n_n48  &  wire20149 ) | ( n_n48  &  wire22696 ) ;
 assign wire2041 = ( n_n53  &  wire120 ) | ( n_n53  &  wire19457 ) | ( n_n53  &  n_n25 ) ;
 assign wire2059 = ( n_n208  &  n_n285  &  n_n230  &  wire190 ) ;
 assign wire2067 = ( n_n5  &  n_n203 ) | ( n_n5  &  wire20149 ) | ( n_n5  &  wire161 ) ;
 assign wire22664 = ( i_15_  &  n_n225  &  n_n253 ) | ( (~ i_15_)  &  n_n225  &  n_n253 ) | ( i_15_  &  n_n225  &  n_n267 ) | ( (~ i_15_)  &  n_n225  &  n_n267 ) ;
 assign wire2072 = ( n_n99  &  n_n100 ) | ( n_n100  &  wire96 ) | ( n_n100  &  wire22664 ) ;
 assign wire2081 = ( n_n260  &  n_n285  &  n_n261  &  wire1340 ) ;
 assign wire22657 = ( i_15_  &  n_n258  &  n_n282 ) | ( i_15_  &  n_n282  &  n_n225 ) | ( (~ i_15_)  &  n_n282  &  n_n225 ) ;
 assign wire2082 = ( n_n37  &  n_n94 ) | ( wire89  &  n_n94 ) | ( n_n94  &  wire22657 ) ;
 assign wire2089 = ( n_n99  &  n_n94 ) | ( n_n94  &  wire96 ) | ( n_n94  &  wire134 ) ;
 assign wire22650 = ( (~ i_15_)  &  n_n225  &  n_n247 ) | ( i_15_  &  n_n225  &  n_n275 ) | ( (~ i_15_)  &  n_n225  &  n_n275 ) ;
 assign wire2103 = ( n_n57  &  wire275 ) | ( n_n57  &  wire262 ) ;
 assign wire2104 = ( n_n56  &  wire198 ) | ( n_n56  &  wire262 ) | ( n_n56  &  wire304 ) ;
 assign wire22631 = ( i_15_  &  n_n258  &  n_n253 ) | ( i_15_  &  n_n225  &  n_n253 ) | ( (~ i_15_)  &  n_n225  &  n_n253 ) ;
 assign wire2122 = ( n_n99  &  n_n53 ) | ( n_n53  &  wire96 ) | ( n_n53  &  wire22631 ) ;
 assign wire2128 = ( n_n56  &  wire301 ) | ( n_n56  &  wire356 ) ;
 assign wire2129 = ( n_n57  &  wire301 ) | ( n_n57  &  wire335 ) | ( n_n57  &  wire304 ) ;
 assign wire2162 = ( n_n4  &  wire128 ) | ( wire911  &  n_n4  &  n_n258 ) ;
 assign wire22598 = ( i_15_  &  n_n242  &  n_n225 ) | ( (~ i_15_)  &  n_n242  &  n_n225 ) | ( i_15_  &  n_n225  &  n_n270 ) | ( (~ i_15_)  &  n_n225  &  n_n270 ) ;
 assign wire22597 = ( i_15_  &  n_n258  &  n_n275 ) | ( i_15_  &  n_n225  &  n_n275 ) | ( (~ i_15_)  &  n_n225  &  n_n275 ) ;
 assign wire2170 = ( n_n3  &  n_n103 ) | ( n_n3  &  wire19457 ) | ( n_n3  &  n_n25 ) ;
 assign wire2173 = ( n_n3  &  n_n37 ) | ( n_n3  &  wire126 ) | ( n_n3  &  wire89 ) ;
 assign wire2174 = ( n_n4  &  n_n37 ) | ( n_n4  &  wire89 ) | ( n_n4  &  n_n104 ) ;
 assign wire2176 = ( wire913  &  n_n258  &  wire169 ) ;
 assign wire2183 = ( wire143  &  _40229 ) | ( wire22341  &  _40229 ) | ( _40226  &  _40229 ) ;
 assign wire2196 = ( n_n197  &  n_n227 ) | ( wire42  &  n_n227 ) | ( n_n227  &  wire441 ) ;
 assign wire2200 = ( n_n216  &  n_n207 ) | ( n_n207  &  n_n212 ) | ( n_n207  &  wire52 ) ;
 assign wire2205 = ( n_n4  &  wire65 ) | ( n_n4  &  wire902  &  n_n256 ) ;
 assign wire2206 = ( wire913  &  n_n258  &  wire278 ) ;
 assign wire2225 = ( n_n2  &  wire187 ) | ( n_n2  &  n_n258  &  wire904 ) ;
 assign wire2235 = ( wire123  &  wire1354 ) | ( n_n258  &  wire899  &  wire1354 ) ;
 assign wire2237 = ( n_n1  &  n_n112 ) | ( n_n1  &  wire52 ) | ( n_n1  &  wire110 ) ;
 assign wire2239 = ( n_n1  &  wire187 ) | ( wire911  &  n_n1  &  n_n258 ) ;
 assign wire22535 = ( i_15_  &  n_n242  &  n_n258 ) | ( i_15_  &  n_n242  &  n_n256 ) | ( (~ i_15_)  &  n_n242  &  n_n256 ) ;
 assign wire2240 = ( n_n2  &  n_n112 ) | ( n_n2  &  wire52 ) | ( n_n2  &  wire22535 ) ;
 assign wire2246 = ( n_n1  &  wire175 ) | ( n_n1  &  n_n258  &  wire900 ) ;
 assign wire22519 = ( i_14_  &  (~ i_13_)  &  i_12_  &  wire907 ) | ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire907 ) ;
 assign wire22515 = ( wire902  &  n_n258 ) | ( n_n258  &  wire897 ) ;
 assign wire22516 = ( i_11_  &  i_15_  &  n_n163  &  n_n256 ) | ( (~ i_11_)  &  i_15_  &  n_n163  &  n_n256 ) | ( i_11_  &  (~ i_15_)  &  n_n163  &  n_n256 ) | ( (~ i_11_)  &  (~ i_15_)  &  n_n163  &  n_n256 ) ;
 assign wire2260 = ( n_n1  &  wire124 ) | ( n_n1  &  wire22515 ) | ( n_n1  &  wire22516 ) ;
 assign wire2263 = ( n_n1  &  wire140 ) | ( n_n1  &  wire182 ) ;
 assign wire22506 = ( n_n258  &  wire898 ) | ( n_n258  &  wire901 ) ;
 assign wire2264 = ( n_n2  &  wire41 ) | ( n_n2  &  wire175 ) | ( n_n2  &  wire22506 ) ;
 assign wire2267 = ( n_n2  &  wire112 ) | ( n_n2  &  wire144 ) ;
 assign wire2268 = ( n_n1  &  wire112 ) | ( n_n1  &  n_n258  &  wire901 ) ;
 assign wire2269 = ( n_n104  &  n_n94 ) | ( wire57  &  n_n94 ) | ( n_n94  &  n_n113 ) ;
 assign wire2291 = ( n_n105  &  n_n94 ) | ( wire41  &  n_n94 ) | ( n_n94  &  wire175 ) ;
 assign wire22475 = ( (~ i_15_)  &  n_n279  &  n_n253 ) | ( i_15_  &  n_n256  &  n_n253 ) | ( (~ i_15_)  &  n_n256  &  n_n253 ) ;
 assign wire22471 = ( i_14_  &  i_13_  &  (~ i_12_)  &  wire908 ) | ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire908 ) ;
 assign wire2306 = ( n_n57  &  wire276 ) | ( n_n57  &  wire182 ) | ( n_n57  &  wire22471 ) ;
 assign wire2311 = ( wire41  &  n_n48 ) | ( n_n48  &  wire175 ) ;
 assign wire2333 = ( wire112  &  n_n48 ) | ( n_n48  &  wire144 ) ;
 assign wire2336 = ( wire124  &  wire1517 ) | ( wire1517  &  wire231 ) ;
 assign wire2344 = ( _793 ) | ( n_n6  &  n_n73 ) | ( n_n6  &  wire320 ) ;
 assign wire22436 = ( wire908  &  n_n256 ) | ( n_n256  &  wire903 ) ;
 assign wire22429 = ( wire907  &  n_n256 ) | ( n_n256  &  wire904 ) ;
 assign wire2364 = ( _897 ) | ( n_n6  &  n_n52 ) | ( n_n6  &  wire22340 ) ;
 assign wire22407 = ( wire907  &  n_n258 ) | ( n_n258  &  wire904 ) ;
 assign wire22408 = ( wire914  &  n_n258 ) | ( n_n258  &  wire904 ) ;
 assign wire2378 = ( wire112  &  n_n53 ) | ( n_n53  &  wire22408 ) ;
 assign wire2392 = ( n_n53  &  n_n112 ) | ( n_n53  &  wire52 ) | ( n_n53  &  wire110 ) ;
 assign wire2393 = ( n_n48  &  wire123 ) | ( n_n48  &  wire140 ) | ( n_n48  &  wire182 ) ;
 assign wire2398 = ( n_n48  &  n_n112 ) | ( n_n48  &  wire52 ) | ( n_n48  &  wire110 ) ;
 assign wire22387 = ( i_15_  &  n_n256  &  n_n275 ) | ( (~ i_15_)  &  n_n256  &  n_n275 ) | ( i_15_  &  n_n256  &  n_n259 ) | ( (~ i_15_)  &  n_n256  &  n_n259 ) ;
 assign wire2403 = ( n_n100  &  wire123 ) | ( n_n100  &  wire124 ) | ( n_n100  &  wire22387 ) ;
 assign wire2425 = ( n_n56  &  wire357 ) | ( n_n56  &  n_n222  &  wire904 ) ;
 assign wire22376 = ( n_n267  &  _40124 ) | ( n_n267  &  _40125 ) ;
 assign wire2426 = ( n_n57  &  wire76 ) | ( n_n57  &  wire229 ) | ( n_n57  &  wire22376 ) ;
 assign wire2427 = ( n_n285  &  n_n266  &  n_n230  &  wire1755 ) ;
 assign wire22374 = ( n_n267  &  _40133 ) | ( n_n267  &  _40134 ) ;
 assign wire2428 = ( n_n56  &  wire76 ) | ( n_n56  &  wire229 ) | ( n_n56  &  wire22374 ) ;
 assign wire2472 = ( n_n3  &  n_n78 ) | ( n_n3  &  wire65 ) | ( n_n3  &  wire276 ) ;
 assign wire2473 = ( n_n4  &  n_n199 ) | ( n_n4  &  n_n73 ) | ( n_n4  &  wire22335 ) ;
 assign wire2478 = ( n_n56  &  wire40 ) | ( n_n56  &  n_n74 ) | ( n_n56  &  wire140 ) ;
 assign wire2486 = ( _1515 ) | ( _1516 ) | ( n_n56  &  wire346 ) ;
 assign wire2491 = ( _1509 ) | ( _1510 ) | ( n_n57  &  wire433 ) ;
 assign wire2495 = ( wire51  &  n_n53 ) | ( n_n53  &  n_n90 ) | ( n_n53  &  wire448 ) ;
 assign wire22290 = ( i_15_  &  n_n281  &  n_n253 ) | ( i_15_  &  n_n256  &  n_n253 ) | ( (~ i_15_)  &  n_n256  &  n_n253 ) ;
 assign wire2507 = ( n_n48  &  wire57 ) | ( n_n48  &  n_n113 ) | ( n_n48  &  n_n39 ) ;
 assign wire2508 = ( n_n53  &  wire61 ) | ( n_n53  &  n_n79 ) | ( n_n53  &  n_n101 ) ;
 assign wire2520 = ( n_n57  &  n_n246 ) | ( n_n57  &  wire73 ) | ( n_n57  &  wire220 ) ;
 assign wire22275 = ( wire66 ) | ( wire274 ) | ( wire899  &  n_n256 ) ;
 assign wire22276 = ( n_n107 ) | ( wire83 ) | ( wire220 ) | ( wire22273 ) ;
 assign wire2532 = ( n_n56  &  n_n246 ) | ( n_n56  &  n_n147 ) | ( n_n56  &  wire291 ) ;
 assign wire2533 = ( n_n57  &  wire63 ) | ( n_n57  &  n_n147 ) | ( n_n57  &  wire291 ) ;
 assign wire2534 = ( n_n56  &  wire223 ) | ( n_n220  &  wire911  &  n_n56 ) ;
 assign wire22259 = ( n_n275  &  _39536 ) | ( n_n275  &  _39537 ) ;
 assign wire2545 = ( _1338 ) | ( n_n94  &  wire807 ) | ( n_n94  &  _39809 ) ;
 assign wire2560 = ( n_n111  &  n_n100 ) | ( n_n100  &  wire158 ) | ( n_n100  &  wire342 ) ;
 assign wire2561 = ( wire200  &  n_n94 ) | ( n_n94  &  wire85 ) | ( n_n94  &  wire78 ) ;
 assign wire2571 = ( n_n56  &  n_n50 ) | ( n_n56  &  wire300 ) | ( n_n56  &  wire311 ) ;
 assign wire2572 = ( n_n57  &  wire55 ) | ( wire914  &  n_n228  &  n_n57 ) ;
 assign wire2581 = ( wire63  &  n_n94 ) | ( wire913  &  n_n258  &  n_n94 ) ;
 assign wire2583 = ( wire75  &  n_n100 ) | ( n_n100  &  n_n58 ) | ( n_n100  &  wire223 ) ;
 assign wire22206 = ( n_n247  &  _39753 ) | ( n_n247  &  _39754 ) ;
 assign wire22210 = ( wire66 ) | ( wire22208 ) | ( wire899  &  n_n256 ) ;
 assign wire22211 = ( n_n107 ) | ( wire83 ) | ( wire220 ) | ( wire291 ) ;
 assign wire2601 = ( n_n260  &  n_n285  &  n_n263  &  wire1113 ) ;
 assign wire2602 = ( _1427 ) | ( _1428 ) | ( _1429 ) ;
 assign wire2623 = ( n_n94  &  wire232 ) | ( n_n94  &  wire110 ) | ( n_n94  &  wire274 ) ;
 assign wire22170 = ( (~ i_15_)  &  n_n228  &  n_n270 ) | ( i_15_  &  n_n222  &  n_n270 ) | ( (~ i_15_)  &  n_n222  &  n_n270 ) ;
 assign wire2631 = ( _1473 ) | ( n_n48  &  wire345 ) | ( n_n48  &  wire22170 ) ;
 assign wire22162 = ( n_n267  &  _39683 ) | ( n_n267  &  _39684 ) ;
 assign wire2637 = ( wire95  &  n_n53 ) | ( n_n53  &  wire220 ) | ( n_n53  &  wire22162 ) ;
 assign wire22167 = ( wire66 ) | ( wire22164 ) | ( wire905  &  n_n222 ) ;
 assign wire22168 = ( wire73 ) | ( n_n107 ) | ( wire187 ) | ( wire220 ) ;
 assign wire2640 = ( n_n53  &  wire62 ) | ( n_n281  &  wire911  &  n_n53 ) ;
 assign wire2652 = ( n_n6  &  wire166 ) | ( n_n6  &  wire180 ) | ( n_n6  &  n_n50 ) ;
 assign wire22139 = ( n_n220  &  wire911 ) | ( wire907  &  n_n228 ) ;
 assign wire2659 = ( n_n53  &  wire22139 ) | ( wire907  &  n_n222  &  n_n53 ) ;
 assign wire2676 = ( n_n6  &  n_n102 ) | ( n_n6  &  wire807 ) | ( n_n6  &  wire311 ) ;
 assign wire2703 = ( n_n5  &  wire55 ) | ( n_n5  &  n_n87 ) | ( n_n5  &  wire342 ) ;
 assign wire2708 = ( n_n5  &  n_n246 ) | ( n_n5  &  n_n147 ) | ( n_n5  &  wire291 ) ;
 assign wire2709 = ( n_n6  &  wire63 ) | ( n_n6  &  n_n147 ) | ( n_n6  &  wire291 ) ;
 assign wire2725 = ( n_n240  &  n_n207 ) | ( n_n207  &  n_n17 ) | ( n_n207  &  wire514 ) ;
 assign wire2726 = ( wire49  &  n_n227 ) | ( n_n228  &  wire908  &  n_n227 ) ;
 assign wire22058 = ( wire19578 ) | ( wire300 ) | ( n_n222  &  wire906 ) ;
 assign wire22059 = ( wire99 ) | ( n_n46 ) | ( wire81 ) | ( wire77 ) ;
 assign wire2774 = ( n_n5  &  n_n240 ) | ( n_n5  &  wire63 ) | ( n_n5  &  wire50 ) ;
 assign wire22033 = ( n_n275  &  _39902 ) | ( n_n275  &  _39903 ) ;
 assign wire22024 = ( n_n267  &  _39890 ) | ( n_n267  &  _39891 ) ;
 assign wire2784 = ( n_n6  &  wire274 ) | ( n_n281  &  n_n6  &  wire899 ) ;
 assign wire22001 = ( n_n220  &  wire911 ) | ( n_n258  &  wire903 ) ;
 assign wire2813 = ( n_n2  &  wire95 ) | ( n_n220  &  n_n2  &  wire898 ) ;
 assign wire2814 = ( n_n1  &  wire95 ) | ( n_n220  &  n_n1  &  wire901 ) ;
 assign wire2822 = ( _1166 ) | ( _1167 ) | ( _1168 ) ;
 assign wire21979 = ( wire514 ) | ( wire325 ) | ( wire911  &  n_n225 ) ;
 assign wire21980 = ( wire73 ) | ( wire60 ) | ( n_n18 ) | ( wire21977 ) ;
 assign wire2825 = ( n_n1  &  wire21979 ) | ( n_n1  &  wire21980 ) ;
 assign wire2827 = ( wire75  &  wire1423 ) | ( n_n220  &  wire899  &  wire1423 ) ;
 assign wire21971 = ( n_n275  &  _39950 ) | ( n_n275  &  _39951 ) ;
 assign wire2830 = ( n_n2  &  wire63 ) | ( n_n2  &  wire21971 ) ;
 assign wire2831 = ( n_n1  &  n_n257 ) | ( n_n1  &  wire63 ) | ( n_n1  &  wire50 ) ;
 assign wire2839 = ( _1203 ) | ( _1204 ) | ( _1205 ) ;
 assign wire21953 = ( wire112 ) | ( wire65 ) | ( wire902  &  n_n225 ) ;
 assign wire21954 = ( wire200 ) | ( wire49 ) | ( wire78 ) | ( n_n79 ) ;
 assign wire2842 = ( n_n1  &  wire21953 ) | ( n_n1  &  wire21954 ) ;
 assign wire2845 = ( n_n4  &  wire40 ) | ( n_n4  &  n_n74 ) | ( n_n4  &  wire346 ) ;
 assign wire2864 = ( n_n4  &  wire95 ) | ( n_n220  &  n_n4  &  wire898 ) ;
 assign wire2874 = ( wire75  &  n_n4 ) | ( n_n4  &  wire50 ) ;
 assign wire21913 = ( n_n220  &  wire901 ) | ( n_n258  &  wire903 ) ;
 assign wire2883 = ( n_n4  &  wire514 ) | ( n_n4  &  n_n68 ) | ( n_n4  &  wire325 ) ;
 assign wire2885 = ( n_n3  &  wire123 ) | ( n_n3  &  wire100 ) ;
 assign wire2888 = ( n_n208  &  n_n284  &  n_n285  &  wire992 ) ;
 assign wire2889 = ( _1760 ) | ( n_n3  &  wire343 ) | ( n_n3  &  wire431 ) ;
 assign wire2893 = ( n_n3  &  wire154 ) | ( n_n3  &  n_n247  &  _36683 ) ;
 assign wire21892 = ( n_n220  &  wire898 ) | ( n_n220  &  wire897 ) ;
 assign wire2917 = ( n_n3  &  n_n29 ) | ( n_n3  &  n_n80 ) | ( n_n3  &  wire61 ) ;
 assign wire2918 = ( n_n4  &  n_n24 ) | ( n_n4  &  wire104 ) | ( n_n4  &  wire228 ) ;
 assign wire2919 = ( wire154  &  n_n94 ) | ( n_n94  &  n_n34 ) | ( n_n94  &  wire263 ) ;
 assign wire2920 = ( n_n260  &  n_n285  &  n_n261  &  wire1835 ) ;
 assign wire2927 = ( _2145 ) | ( _2146 ) ;
 assign wire2928 = ( _2137 ) | ( _2138 ) | ( _2139 ) ;
 assign wire2929 = ( n_n100  &  n_n97 ) | ( n_n100  &  wire226 ) | ( n_n100  &  wire361 ) ;
 assign wire2942 = ( n_n53  &  wire61 ) | ( n_n222  &  wire908  &  n_n53 ) ;
 assign wire2943 = ( n_n247  &  _36974  &  _39131 ) | ( n_n247  &  _36975  &  _39131 ) ;
 assign wire2952 = ( n_n48  &  wire230 ) | ( n_n222  &  n_n48  &  _36699 ) ;
 assign wire2973 = ( n_n37  &  n_n48 ) | ( n_n83  &  n_n48 ) | ( wire64  &  n_n48 ) ;
 assign wire2974 = ( n_n53  &  wire102 ) | ( n_n53  &  n_n86 ) | ( n_n53  &  wire263 ) ;
 assign wire21821 = ( wire902  &  n_n222 ) | ( n_n222  &  wire901 ) ;
 assign wire21805 = ( i_14_  &  i_13_  &  (~ i_12_)  &  wire899 ) | ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  wire899 ) ;
 assign wire21807 = ( wire84 ) | ( n_n71 ) | ( n_n69 ) | ( wire143 ) ;
 assign wire3003 = ( n_n5  &  n_n29 ) | ( n_n5  &  n_n80 ) | ( n_n5  &  wire61 ) ;
 assign wire3004 = ( n_n6  &  n_n24 ) | ( n_n6  &  wire104 ) | ( n_n6  &  wire228 ) ;
 assign wire21789 = ( i_14_  &  i_13_  &  (~ i_12_)  &  wire898 ) | ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  wire898 ) ;
 assign wire3012 = ( n_n6  &  n_n52 ) | ( n_n6  &  wire807 ) | ( n_n6  &  wire21789 ) ;
 assign wire21785 = ( n_n225  &  wire901 ) | ( n_n220  &  wire897 ) ;
 assign wire3043 = ( n_n5  &  n_n37 ) | ( n_n5  &  n_n83 ) | ( n_n5  &  wire64 ) ;
 assign wire3045 = ( n_n285  &  n_n271  &  n_n230  &  wire1600 ) ;
 assign wire3056 = ( n_n94  &  n_n78 ) | ( n_n94  &  n_n69 ) | ( n_n94  &  wire230 ) ;
 assign wire3065 = ( n_n260  &  n_n285  &  n_n263  &  wire236 ) ;
 assign wire3072 = ( n_n220  &  wire899  &  wire1196 ) ;
 assign wire3080 = ( n_n285  &  n_n271  &  n_n230  &  wire1251 ) ;
 assign wire3098 = ( n_n285  &  n_n271  &  n_n230  &  wire1250 ) ;
 assign wire3106 = ( n_n56  &  wire100 ) | ( n_n56  &  wire1199 ) ;
 assign wire3109 = ( n_n57  &  wire100 ) | ( n_n57  &  wire472 ) ;
 assign wire3120 = ( n_n1  &  n_n97 ) | ( n_n1  &  wire226 ) | ( n_n1  &  wire361 ) ;
 assign wire3178 = ( n_n3  &  n_n44 ) | ( n_n3  &  wire270 ) | ( n_n3  &  wire21668 ) ;
 assign wire3179 = ( n_n4  &  n_n88 ) | ( n_n4  &  n_n44 ) | ( n_n4  &  wire21668 ) ;
 assign wire3187 = ( n_n267  &  _38965  &  _38968 ) | ( n_n267  &  _38966  &  _38968 ) ;
 assign wire3190 = ( n_n265  &  wire200 ) | ( n_n265  &  wire158 ) ;
 assign wire21658 = ( n_n220  &  wire914 ) | ( n_n220  &  wire911 ) ;
 assign wire3203 = ( n_n260  &  n_n273  &  n_n285  &  wire1773 ) ;
 assign wire21650 = ( n_n220  &  wire898 ) | ( n_n220  &  wire901 ) ;
 assign wire3211 = ( n_n2  &  n_n20 ) | ( n_n2  &  wire375 ) | ( n_n2  &  wire21650 ) ;
 assign wire3213 = ( n_n3  &  n_n37 ) | ( n_n3  &  n_n83 ) | ( n_n3  &  wire64 ) ;
 assign wire3214 = ( n_n4  &  wire102 ) | ( n_n4  &  n_n86 ) | ( n_n4  &  wire263 ) ;
 assign wire3219 = ( n_n1  &  n_n20 ) | ( n_n1  &  wire375 ) | ( n_n1  &  wire1792 ) ;
 assign wire21642 = ( wire236 ) | ( wire230 ) | ( wire902  &  n_n256 ) ;
 assign wire3220 = ( n_n2  &  wire1792 ) | ( n_n2  &  wire21642 ) ;
 assign wire3221 = ( _2306 ) | ( _2307 ) ;
 assign wire21639 = ( wire362 ) | ( wire87 ) | ( n_n220  &  wire914 ) ;
 assign wire21640 = ( n_n42 ) | ( wire59 ) | ( wire243 ) | ( wire428 ) ;
 assign wire3222 = ( n_n1  &  wire21639 ) | ( n_n1  &  wire21640 ) ;
 assign wire3228 = ( n_n3  &  wire102 ) | ( n_n3  &  n_n86 ) | ( n_n3  &  wire263 ) ;
 assign wire3232 = ( wire48  &  n_n127 ) | ( wire913  &  n_n220  &  n_n127 ) ;
 assign wire21584 = ( n_n279  &  wire912 ) | ( n_n279  &  wire900 ) ;
 assign wire21576 = ( n_n279  &  wire912 ) | ( n_n279  &  wire901 ) ;
 assign wire3296 = ( n_n264  &  n_n273  &  n_n285  &  wire1485 ) ;
 assign wire3297 = ( wire913  &  n_n281  &  wire185 ) ;
 assign wire3324 = ( wire913  &  n_n281  &  _38794 ) | ( n_n281  &  wire903  &  _38794 ) ;
 assign wire21536 = ( wire913  &  n_n279 ) | ( n_n279  &  wire897 ) ;
 assign wire3375 = ( n_n100  &  wire167 ) | ( n_n100  &  wire235 ) | ( n_n100  &  wire157 ) ;
 assign wire3376 = ( wire268  &  n_n94 ) | ( n_n94  &  wire436 ) | ( n_n94  &  wire157 ) ;
 assign wire3382 = ( n_n285  &  n_n266  &  n_n230  &  wire1530 ) ;
 assign wire3393 = ( wire1378  &  wire1377 ) ;
 assign wire3400 = ( n_n48  &  n_n93 ) | ( n_n48  &  n_n90 ) | ( n_n48  &  wire21389 ) ;
 assign wire3401 = ( n_n53  &  wire71 ) | ( n_n53  &  n_n102 ) | ( n_n53  &  wire77 ) ;
 assign wire3402 = ( n_n285  &  n_n271  &  n_n230  &  wire1095 ) ;
 assign wire3409 = ( n_n279  &  wire1094  &  _38556 ) | ( n_n279  &  wire1094  &  _38558 ) ;
 assign wire3413 = ( n_n56  &  n_n70 ) | ( n_n56  &  wire79 ) | ( n_n56  &  wire413 ) ;
 assign wire3416 = ( n_n56  &  wire264 ) | ( n_n56  &  n_n73 ) | ( n_n56  &  wire19408 ) ;
 assign wire3440 = ( n_n100  &  n_n148 ) | ( n_n100  &  wire210 ) | ( n_n100  &  wire399 ) ;
 assign wire21457 = ( n_n281  &  wire907 ) | ( n_n281  &  wire904 ) ;
 assign wire21458 = ( n_n281  &  wire914 ) | ( n_n281  &  wire908 ) ;
 assign wire3441 = ( n_n94  &  wire21457 ) | ( n_n94  &  wire21458 ) ;
 assign wire3442 = ( n_n281  &  wire903  &  wire168 ) ;
 assign wire3447 = ( n_n94  &  wire281 ) | ( n_n94  &  wire338 ) ;
 assign wire3451 = ( n_n56  &  n_n253  &  _38483 ) | ( n_n56  &  n_n253  &  _38485 ) ;
 assign wire3469 = ( n_n1  &  wire255 ) | ( n_n1  &  wire242 ) ;
 assign wire3470 = ( n_n264  &  n_n273  &  n_n285  &  wire1163 ) ;
 assign wire3480 = ( n_n3  &  wire71 ) | ( n_n279  &  n_n3  &  wire904 ) ;
 assign wire3499 = ( n_n2  &  wire281 ) | ( n_n2  &  wire338 ) | ( n_n2  &  wire1101 ) ;
 assign wire3500 = ( n_n1  &  n_n60 ) | ( n_n1  &  wire210 ) | ( n_n1  &  wire1101 ) ;
 assign wire3520 = ( n_n265  &  wire252 ) | ( n_n265  &  n_n81 ) | ( n_n265  &  wire86 ) ;
 assign wire21383 = ( i_15_  &  n_n242  &  n_n279 ) | ( (~ i_15_)  &  n_n242  &  n_n279 ) | ( i_15_  &  n_n279  &  n_n247 ) | ( (~ i_15_)  &  n_n279  &  n_n247 ) ;
 assign wire3544 = ( wire72  &  n_n57 ) | ( n_n57  &  n_n257 ) | ( n_n57  &  n_n7 ) ;
 assign wire3550 = ( n_n57  &  wire44 ) | ( n_n57  &  n_n252 ) | ( n_n57  &  n_n15 ) ;
 assign wire3551 = ( _2959 ) | ( _2960 ) | ( _2961 ) ;
 assign wire3562 = ( _3011 ) | ( _3012 ) ;
 assign wire3563 = ( _3006 ) | ( _3007 ) | ( _3008 ) ;
 assign wire3565 = ( _3000 ) | ( _3001 ) | ( _3002 ) ;
 assign wire3584 = ( n_n57  &  wire246 ) | ( n_n57  &  wire256 ) ;
 assign wire3585 = ( n_n281  &  n_n56  &  wire906 ) ;
 assign wire3627 = ( n_n282  &  _35947  &  _38361 ) | ( n_n282  &  _35948  &  _38361 ) ;
 assign wire21266 = ( n_n220  &  wire912 ) | ( wire913  &  n_n258 ) ;
 assign wire3629 = ( n_n268  &  wire160 ) | ( n_n268  &  n_n59 ) | ( n_n268  &  wire21266 ) ;
 assign wire3642 = ( wire95  &  n_n3 ) | ( n_n3  &  n_n11 ) | ( n_n3  &  n_n148 ) ;
 assign wire3653 = ( n_n54  &  n_n3 ) | ( n_n3  &  n_n99 ) | ( n_n3  &  wire96 ) ;
 assign wire3662 = ( n_n4  &  wire912  &  n_n258 ) ;
 assign wire3674 = ( _3195 ) | ( _3196 ) | ( _3197 ) ;
 assign wire3680 = ( _3178 ) | ( _3179 ) ;
 assign wire3681 = ( _3173 ) | ( _3174 ) | ( _3175 ) ;
 assign wire3682 = ( _3187 ) | ( _3188 ) | ( _3189 ) ;
 assign wire3688 = ( n_n3  &  wire73 ) | ( n_n3  &  n_n65 ) | ( n_n3  &  n_n12 ) ;
 assign wire3689 = ( n_n4  &  wire44 ) | ( n_n4  &  n_n252 ) | ( n_n4  &  n_n15 ) ;
 assign wire3712 = ( n_n152  &  n_n220  &  wire914 ) ;
 assign wire3725 = ( wire54  &  n_n128 ) | ( n_n111  &  n_n128 ) | ( n_n110  &  n_n128 ) ;
 assign wire3726 = ( wire48  &  n_n130 ) | ( wire54  &  n_n130 ) | ( n_n110  &  n_n130 ) ;
 assign wire3733 = ( wire48  &  n_n121 ) | ( wire54  &  n_n121 ) | ( n_n110  &  n_n121 ) ;
 assign wire3736 = ( n_n9  &  n_n3 ) | ( n_n3  &  wire63 ) | ( n_n3  &  wire184 ) ;
 assign wire3778 = ( wire453  &  n_n94 ) | ( wire71  &  n_n94 ) | ( n_n94  &  n_n97 ) ;
 assign wire3790 = ( wire199  &  n_n94 ) | ( wire70  &  n_n94 ) | ( n_n94  &  n_n14 ) ;
 assign wire3791 = ( n_n247  &  _34581  &  _38049 ) | ( n_n247  &  _34582  &  _38049 ) ;
 assign wire3821 = ( n_n264  &  n_n285  &  n_n263  &  wire1323 ) ;
 assign wire3837 = ( n_n5  &  wire87 ) | ( wire914  &  n_n5  &  n_n225 ) ;
 assign wire3843 = ( wire63  &  n_n48 ) | ( n_n228  &  wire902  &  n_n48 ) ;
 assign wire21009 = ( n_n247  &  _38006 ) | ( n_n247  &  _38007 ) ;
 assign wire3896 = ( wire118  &  n_n5 ) | ( n_n5  &  wire199 ) | ( n_n5  &  n_n144 ) ;
 assign wire3924 = ( n_n268  &  wire95 ) | ( n_n268  &  n_n11 ) | ( n_n268  &  wire157 ) ;
 assign wire3931 = ( n_n1  &  wire72 ) | ( n_n228  &  n_n1  &  wire902 ) ;
 assign wire20917 = ( n_n229  &  n_n165  &  n_n284 ) | ( n_n165  &  n_n284  &  n_n283 ) ;
 assign wire3946 = ( n_n165  &  n_n283  &  wire19294  &  wire923 ) ;
 assign wire3967 = ( n_n5  &  wire100 ) | ( n_n5  &  wire281 ) ;
 assign wire3968 = ( n_n6  &  wire118 ) | ( n_n6  &  wire70 ) | ( n_n6  &  n_n14 ) ;
 assign wire3975 = ( n_n4  &  wire166 ) | ( wire905  &  n_n4  &  n_n225 ) ;
 assign wire3976 = ( n_n94  &  wire130 ) | ( wire911  &  n_n228  &  n_n94 ) ;
 assign wire20874 = ( i_15_  &  n_n242  &  n_n258 ) | ( i_15_  &  n_n242  &  n_n256 ) | ( (~ i_15_)  &  n_n242  &  n_n256 ) ;
 assign wire3988 = ( n_n207  &  n_n112 ) | ( n_n207  &  wire52 ) | ( n_n207  &  wire20874 ) ;
 assign wire20875 = ( i_15_  &  n_n258  &  n_n259 ) | ( i_15_  &  n_n256  &  n_n259 ) | ( (~ i_15_)  &  n_n256  &  n_n259 ) ;
 assign wire4004 = ( n_n1  &  wire72 ) | ( n_n1  &  n_n226 ) | ( n_n1  &  n_n257 ) ;
 assign wire4005 = ( n_n2  &  wire66 ) | ( n_n2  &  wire899  &  n_n256 ) ;
 assign wire4016 = ( wire75  &  n_n48 ) | ( n_n206  &  n_n48 ) | ( wire44  &  n_n48 ) ;
 assign wire20839 = ( i_14_  &  i_13_  &  i_12_  &  wire905 ) | ( (~ i_14_)  &  i_13_  &  i_12_  &  wire905 ) | ( i_14_  &  i_13_  &  (~ i_12_)  &  wire905 ) | ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire905 ) ;
 assign wire20840 = ( (~ i_14_)  &  i_13_  &  i_12_  &  wire899 ) | ( i_14_  &  (~ i_13_)  &  i_12_  &  wire899 ) | ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire899 ) | ( i_14_  &  i_13_  &  (~ i_12_)  &  wire899 ) | ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire899 ) | ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  wire899 ) ;
 assign wire4036 = ( n_n5  &  wire60 ) | ( wire911  &  n_n279  &  n_n5 ) ;
 assign wire4044 = ( wire72  &  n_n57 ) | ( wire905  &  n_n258  &  n_n57 ) ;
 assign wire4056 = ( wire72  &  n_n56 ) | ( wire905  &  n_n258  &  n_n56 ) ;
 assign wire4062 = ( wire79  &  n_n48 ) | ( wire905  &  n_n256  &  n_n48 ) ;
 assign wire4081 = ( n_n4  &  wire19738 ) | ( wire913  &  n_n4  &  n_n256 ) ;
 assign wire4100 = ( wire118  &  n_n100 ) | ( n_n220  &  wire899  &  n_n100 ) ;
 assign wire4117 = ( wire79  &  n_n94 ) | ( n_n94  &  n_n20 ) | ( n_n94  &  wire83 ) ;
 assign wire4120 = ( wire79  &  n_n100 ) | ( wire899  &  n_n256  &  n_n100 ) ;
 assign wire4159 = ( wire250  &  wire1231 ) | ( n_n281  &  wire899  &  wire1231 ) ;
 assign wire4170 = ( wire250  &  wire1141 ) | ( n_n281  &  wire899  &  wire1141 ) ;
 assign wire4183 = ( n_n6  &  wire57 ) | ( wire914  &  n_n6  &  n_n279 ) ;
 assign wire4202 = ( i_7_  &  i_6_  &  n_n165  &  wire19294 ) ;
 assign wire20637 = ( n_n260  &  n_n229  &  n_n165 ) | ( n_n229  &  n_n165  &  n_n284 ) ;
 assign wire20638 = ( n_n260  &  n_n165  &  n_n283 ) | ( n_n165  &  n_n284  &  n_n283 ) ;
 assign wire4248 = ( n_n4  &  wire101 ) | ( n_n281  &  wire914  &  n_n4 ) ;
 assign wire4267 = ( n_n106  &  n_n265 ) | ( n_n265  &  wire268 ) | ( n_n265  &  wire101 ) ;
 assign wire4276 = ( _4013 ) | ( _4014 ) | ( _4015 ) ;
 assign wire4281 = ( _4005 ) | ( _4006 ) | ( _4007 ) ;
 assign wire20585 = ( n_n220  &  wire907 ) | ( n_n220  &  wire903 ) ;
 assign wire4285 = ( n_n4  &  n_n73 ) | ( n_n4  &  wire19408 ) | ( n_n4  &  wire20585 ) ;
 assign wire4313 = ( n_n111  &  n_n1 ) | ( n_n1  &  n_n32 ) | ( n_n1  &  wire85 ) ;
 assign wire4330 = ( n_n100  &  wire19578 ) | ( n_n222  &  wire906  &  n_n100 ) ;
 assign wire20512 = ( wire20510 ) | ( n_n275  &  _35051 ) | ( n_n275  &  _35052 ) ;
 assign wire20513 = ( wire75 ) | ( wire72 ) | ( _37370 ) ;
 assign wire20514 = ( wire73 ) | ( n_n65 ) | ( wire160 ) | ( wire184 ) ;
 assign wire4373 = ( n_n57  &  wire55 ) | ( n_n57  &  n_n42 ) | ( n_n57  &  wire81 ) ;
 assign wire4380 = ( wire137  &  n_n100 ) | ( wire113  &  n_n100 ) ;
 assign wire4409 = ( _4295 ) | ( _4296 ) | ( _4297 ) ;
 assign wire4417 = ( wire75  &  n_n57 ) | ( wire913  &  n_n281  &  n_n57 ) ;
 assign wire4418 = ( n_n264  &  n_n285  &  n_n261  &  n_n267 ) ;
 assign wire4423 = ( n_n6  &  wire19578 ) | ( n_n6  &  n_n222  &  wire906 ) ;
 assign wire4463 = ( _4271 ) | ( _4272 ) | ( _4273 ) ;
 assign wire20365 = ( wire913  &  n_n258 ) | ( n_n228  &  wire897 ) ;
 assign wire4506 = ( n_n6  &  wire137 ) | ( n_n6  &  wire113 ) | ( n_n6  &  n_n10 ) ;
 assign wire4520 = ( n_n53  &  wire225 ) | ( n_n53  &  wire130 ) ;
 assign wire4551 = ( n_n53  &  wire246 ) | ( n_n53  &  wire256 ) ;
 assign wire4573 = ( wire73  &  n_n48 ) | ( n_n65  &  n_n48 ) | ( n_n48  &  wire83 ) ;
 assign wire4574 = ( wire44  &  n_n53 ) | ( n_n53  &  n_n252 ) | ( n_n53  &  n_n15 ) ;
 assign wire4617 = ( i_7_  &  i_6_  &  wire1829 ) | ( (~ i_7_)  &  i_6_  &  wire1829 ) ;
 assign wire4618 = ( i_7_  &  i_6_  &  n_n284  &  n_n118 ) ;
 assign wire20213 = ( n_n229  &  n_n165  &  n_n284 ) | ( n_n165  &  n_n284  &  n_n283 ) ;
 assign wire4636 = ( n_n132  &  wire1575 ) | ( wire1575  &  wire20213 ) ;
 assign wire4641 = ( wire1797  &  wire1796 ) ;
 assign wire4656 = ( n_n56  &  wire89 ) | ( wire907  &  n_n56  &  n_n222 ) ;
 assign wire20180 = ( n_n228  &  wire898 ) | ( n_n281  &  wire906 ) ;
 assign wire4690 = ( n_n151  &  n_n5 ) | ( wire75  &  n_n5 ) | ( n_n206  &  n_n5 ) ;
 assign wire4691 = ( n_n6  &  wire225 ) | ( n_n220  &  n_n6  &  wire911 ) ;
 assign wire4711 = ( n_n6  &  wire79 ) | ( n_n6  &  wire899  &  n_n256 ) ;
 assign wire4727 = ( n_n5  &  wire87 ) | ( wire914  &  n_n5  &  n_n225 ) ;
 assign wire4750 = ( n_n6  &  n_n105 ) | ( n_n6  &  wire71 ) | ( n_n6  &  n_n97 ) ;
 assign wire20107 = ( n_n220  &  wire911 ) | ( n_n281  &  wire903 ) ;
 assign wire4766 = ( n_n151  &  n_n94 ) | ( n_n206  &  n_n94 ) | ( n_n94  &  wire20107 ) ;
 assign wire4790 = ( n_n242  &  _34536  &  _37766 ) | ( n_n242  &  _34537  &  _37766 ) ;
 assign wire20089 = ( i_14_  &  i_13_  &  i_12_  &  wire906 ) | ( (~ i_14_)  &  i_13_  &  i_12_  &  wire906 ) | ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire906 ) | ( i_14_  &  i_13_  &  (~ i_12_)  &  wire906 ) | ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  wire906 ) | ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire906 ) ;
 assign wire20090 = ( (~ i_14_)  &  i_13_  &  i_12_  &  wire900 ) | ( i_14_  &  (~ i_13_)  &  i_12_  &  wire900 ) | ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire900 ) | ( i_14_  &  i_13_  &  (~ i_12_)  &  wire900 ) | ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire900 ) | ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  wire900 ) ;
 assign wire4800 = ( n_n94  &  wire20089 ) | ( n_n94  &  wire20090 ) ;
 assign wire20086 = ( (~ i_14_)  &  i_13_  &  i_12_  &  wire898 ) | ( i_14_  &  (~ i_13_)  &  i_12_  &  wire898 ) | ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire898 ) | ( i_14_  &  i_13_  &  (~ i_12_)  &  wire898 ) | ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire898 ) | ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  wire898 ) ;
 assign wire20087 = ( i_14_  &  i_13_  &  i_12_  &  wire904 ) | ( (~ i_14_)  &  i_13_  &  i_12_  &  wire904 ) | ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire904 ) | ( i_14_  &  i_13_  &  (~ i_12_)  &  wire904 ) | ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  wire904 ) | ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire904 ) ;
 assign wire4805 = ( n_n94  &  wire20086 ) | ( n_n94  &  wire20087 ) ;
 assign wire4807 = ( wire273  &  n_n100 ) | ( wire200  &  n_n100 ) | ( n_n100  &  wire157 ) ;
 assign wire4808 = ( wire268  &  n_n94 ) | ( wire200  &  n_n94 ) | ( n_n94  &  wire277 ) ;
 assign wire4817 = ( n_n94  &  wire190 ) | ( n_n94  &  wire198 ) | ( n_n94  &  wire119 ) ;
 assign wire4844 = ( wire73  &  n_n100 ) | ( n_n65  &  n_n100 ) | ( n_n12  &  n_n100 ) ;
 assign wire4845 = ( wire70  &  n_n94 ) | ( n_n94  &  n_n14 ) | ( n_n94  &  wire256 ) ;
 assign wire4849 = ( n_n94  &  wire123 ) | ( n_n94  &  wire100 ) | ( n_n94  &  wire227 ) ;
 assign wire4856 = ( n_n60  &  n_n94 ) | ( n_n9  &  n_n94 ) | ( wire63  &  n_n94 ) ;
 assign wire4869 = ( n_n60  &  n_n100 ) | ( wire63  &  n_n100 ) | ( wire137  &  n_n100 ) ;
 assign wire4870 = ( n_n94  &  n_n7 ) | ( n_n94  &  wire50 ) | ( n_n94  &  n_n59 ) ;
 assign wire4871 = ( (~ i_7_)  &  i_6_  &  n_n165  &  wire19294 ) | ( i_7_  &  (~ i_6_)  &  n_n165  &  wire19294 ) ;
 assign wire4890 = ( i_7_  &  i_6_  &  n_n165  &  wire19294 ) ;
 assign wire4892 = ( n_n165  &  n_n273  &  n_n163  &  wire19296 ) ;
 assign wire4896 = ( wire48  &  wire1079 ) | ( wire913  &  n_n220  &  wire1079 ) ;
 assign wire4899 = ( wire48  &  n_n152 ) | ( wire913  &  n_n152  &  n_n220 ) ;
 assign wire4900 = ( i_7_  &  i_6_  &  n_n165  &  wire19294 ) | ( (~ i_7_)  &  i_6_  &  n_n165  &  wire19294 ) | ( i_7_  &  (~ i_6_)  &  n_n165  &  wire19294 ) ;
 assign wire4902 = ( wire48  &  wire1076 ) | ( wire913  &  n_n220  &  wire1076 ) ;
 assign wire4905 = ( wire949  &  n_n128 ) | ( wire949  &  n_n122 ) ;
 assign wire4928 = ( i_7_  &  i_6_  &  n_n260  &  n_n118 ) | ( (~ i_7_)  &  i_6_  &  n_n260  &  n_n118 ) | ( i_7_  &  (~ i_6_)  &  n_n260  &  n_n118 ) ;
 assign wire4939 = ( n_n56  &  wire153 ) | ( n_n56  &  wire41 ) ;
 assign wire4947 = ( wire54  &  n_n128 ) | ( wire913  &  n_n220  &  n_n128 ) ;
 assign wire4974 = ( n_n56  &  wire61 ) | ( n_n279  &  n_n56  &  wire908 ) ;
 assign wire5002 = ( wire95  &  n_n57 ) | ( n_n281  &  wire914  &  n_n57 ) ;
 assign wire5012 = ( n_n282  &  _35947  &  _36525 ) | ( n_n282  &  _35948  &  _36525 ) ;
 assign wire5013 = ( wire95  &  n_n56 ) | ( n_n281  &  wire914  &  n_n56 ) ;
 assign wire5014 = ( n_n57  &  wire63 ) | ( n_n228  &  wire902  &  n_n57 ) ;
 assign wire5023 = ( wire75  &  n_n56 ) | ( wire913  &  n_n281  &  n_n56 ) ;
 assign wire5036 = ( n_n275  &  _35051  &  _36954 ) | ( n_n275  &  _35052  &  _36954 ) ;
 assign wire5047 = ( n_n6  &  wire80 ) | ( n_n6  &  wire908  &  n_n256 ) ;
 assign wire5048 = ( n_n5  &  wire57 ) | ( n_n279  &  n_n5  &  wire912 ) ;
 assign wire5054 = ( n_n6  &  wire42 ) | ( n_n6  &  n_n279  &  wire899 ) ;
 assign wire5059 = ( n_n6  &  wire50 ) | ( n_n281  &  n_n6  &  wire903 ) ;
 assign wire5091 = ( n_n6  &  wire55 ) | ( n_n6  &  n_n279  &  wire912 ) ;
 assign wire5099 = ( n_n6  &  wire273 ) | ( wire914  &  n_n6  &  n_n225 ) ;
 assign wire19848 = ( wire913  &  n_n258 ) | ( n_n228  &  wire897 ) ;
 assign wire5138 = ( wire48  &  n_n124 ) | ( n_n124  &  n_n110 ) | ( n_n124  &  n_n163 ) ;
 assign wire5144 = ( n_n264  &  n_n229  &  n_n165  &  n_n163 ) ;
 assign wire5160 = ( n_n2  &  wire137 ) | ( n_n2  &  wire132 ) ;
 assign wire19814 = ( n_n281  &  wire908 ) | ( n_n228  &  wire897 ) ;
 assign wire5161 = ( n_n1  &  n_n7 ) | ( n_n1  &  wire50 ) | ( n_n1  &  wire19814 ) ;
 assign wire5184 = ( n_n2  &  wire95 ) | ( n_n2  &  n_n11 ) | ( n_n2  &  n_n148 ) ;
 assign wire5205 = ( n_n1  &  wire95 ) | ( n_n1  &  n_n148 ) | ( n_n1  &  wire101 ) ;
 assign wire5215 = ( n_n2  &  wire453 ) | ( wire914  &  n_n2  &  n_n256 ) ;
 assign wire5219 = ( n_n220  &  wire914  &  n_n2 ) ;
 assign wire5228 = ( n_n6  &  wire80 ) | ( n_n6  &  wire908  &  n_n256 ) ;
 assign wire5240 = ( n_n5  &  n_n171 ) | ( n_n5  &  wire56 ) | ( n_n5  &  wire53 ) ;
 assign wire5241 = ( n_n220  &  n_n6  &  wire908 ) ;
 assign wire5242 = ( n_n5  &  n_n22 ) | ( n_n5  &  n_n73 ) | ( n_n5  &  wire19408 ) ;
 assign wire5243 = ( wire897  &  _35097  &  _36218 ) | ( wire897  &  _35099  &  _36218 ) ;
 assign wire5262 = ( n_n6  &  wire19738 ) | ( wire913  &  n_n6  &  n_n256 ) ;
 assign wire19713 = ( i_14_  &  i_13_  &  i_12_  &  wire905 ) | ( (~ i_14_)  &  i_13_  &  i_12_  &  wire905 ) | ( i_14_  &  i_13_  &  (~ i_12_)  &  wire905 ) | ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire905 ) ;
 assign wire19714 = ( (~ i_14_)  &  i_13_  &  i_12_  &  wire899 ) | ( i_14_  &  (~ i_13_)  &  i_12_  &  wire899 ) | ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire899 ) | ( i_14_  &  i_13_  &  (~ i_12_)  &  wire899 ) | ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire899 ) | ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  wire899 ) ;
 assign wire5299 = ( n_n57  &  wire19713 ) | ( n_n57  &  wire19714 ) ;
 assign wire5327 = ( n_n60  &  n_n56 ) | ( n_n56  &  wire63 ) | ( n_n56  &  wire160 ) ;
 assign wire5328 = ( _35954 ) | ( n_n57  &  wire101 ) | ( n_n57  &  _35949 ) ;
 assign wire19683 = ( n_n228  &  wire901 ) | ( n_n281  &  wire904 ) ;
 assign wire5357 = ( _5617 ) | ( _5618 ) | ( _5619 ) ;
 assign wire5362 = ( n_n56  &  wire225 ) | ( n_n56  &  wire130 ) ;
 assign wire19668 = ( wire911  &  n_n228 ) | ( n_n281  &  wire905 ) ;
 assign wire5371 = ( _36091 ) | ( n_n5  &  wire71 ) ;
 assign wire5372 = ( _5604 ) | ( n_n6  &  wire453 ) | ( n_n6  &  wire55 ) ;
 assign wire5390 = ( n_n6  &  wire95 ) | ( n_n281  &  wire914  &  n_n6 ) ;
 assign wire5400 = ( n_n6  &  wire113 ) | ( n_n6  &  wire101 ) ;
 assign wire5411 = ( i_7_  &  i_6_  &  wire943 ) | ( i_7_  &  (~ i_6_)  &  wire943 ) ;
 assign wire5412 = ( i_7_  &  (~ i_6_)  &  n_n284  &  n_n118 ) ;
 assign wire5413 = ( i_7_  &  i_6_  &  n_n284  &  n_n118 ) ;
 assign wire5426 = ( wire54  &  n_n130 ) | ( wire54  &  n_n121 ) | ( wire54  &  n_n122 ) ;
 assign wire5430 = ( wire54  &  wire1687 ) | ( n_n220  &  wire914  &  wire1687 ) ;
 assign wire5441 = ( n_n165  &  n_n283  &  wire19296  &  wire923 ) ;
 assign wire5442 = ( n_n165  &  n_n273  &  n_n163  &  wire19296 ) ;
 assign wire5445 = ( n_n111  &  n_n124 ) | ( wire103  &  n_n124 ) | ( wire266  &  n_n124 ) ;
 assign wire19605 = ( (~ i_9_)  &  (~ i_10_) ) | ( n_n281  &  wire911 ) ;
 assign wire5472 = ( wire19578  &  n_n94 ) | ( n_n222  &  wire906  &  n_n94 ) ;
 assign wire5494 = ( n_n281  &  wire908  &  n_n94 ) ;
 assign wire5509 = ( n_n100  &  n_n7 ) | ( n_n100  &  wire50 ) | ( n_n100  &  n_n59 ) ;
 assign wire19556 = ( n_n228  &  wire898 ) | ( n_n281  &  wire906 ) ;
 assign wire19548 = ( (~ i_14_)  &  i_13_  &  i_12_  &  wire903 ) | ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire903 ) | ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  wire903 ) ;
 assign wire5516 = ( n_n94  &  wire19457 ) | ( n_n94  &  n_n25 ) | ( n_n94  &  wire19548 ) ;
 assign wire5517 = ( wire80  &  n_n100 ) | ( wire902  &  n_n256  &  n_n100 ) ;
 assign wire5544 = ( n_n56  &  wire61 ) | ( n_n279  &  n_n56  &  wire908 ) ;
 assign wire5564 = ( n_n49  &  n_n48 ) | ( n_n48  &  wire71 ) | ( n_n48  &  wire68 ) ;
 assign wire5565 = ( n_n53  &  n_n42 ) | ( n_n53  &  n_n90 ) | ( n_n53  &  wire19384 ) ;
 assign wire5577 = ( n_n56  &  wire63 ) | ( n_n281  &  n_n56  &  wire908 ) ;
 assign wire5588 = ( n_n275  &  _35053  &  _35956 ) | ( n_n275  &  _35054  &  _35956 ) ;
 assign wire5590 = ( n_n281  &  n_n57  &  wire906 ) ;
 assign wire5596 = ( n_n53  &  wire53 ) | ( n_n279  &  n_n53  &  wire897 ) ;
 assign wire5606 = ( wire137  &  n_n53 ) | ( wire132  &  n_n53 ) ;
 assign wire19491 = ( n_n228  &  wire902 ) | ( n_n281  &  wire903 ) ;
 assign wire5617 = ( wire70  &  n_n53 ) | ( n_n220  &  n_n53  &  wire903 ) ;
 assign wire5625 = ( wire70  &  n_n48 ) | ( wire73  &  n_n48 ) | ( n_n12  &  n_n48 ) ;
 assign wire5626 = ( wire73  &  n_n53 ) | ( n_n65  &  n_n53 ) | ( n_n12  &  n_n53 ) ;
 assign wire5640 = ( wire88  &  n_n227 ) | ( n_n80  &  n_n227 ) | ( wire114  &  n_n227 ) ;
 assign wire5642 = ( n_n5  &  wire50 ) | ( n_n281  &  n_n5  &  wire903 ) ;
 assign wire5643 = ( n_n6  &  wire50 ) | ( n_n6  &  n_n228  &  wire897 ) ;
 assign wire5650 = ( n_n5  &  wire165 ) | ( n_n5  &  wire167 ) ;
 assign wire5651 = ( n_n6  &  wire199 ) | ( n_n6  &  wire70 ) | ( n_n6  &  n_n14 ) ;
 assign wire5656 = ( n_n5  &  wire246 ) | ( n_n5  &  wire256 ) ;
 assign wire19469 = ( n_n228  &  wire900 ) | ( n_n281  &  wire904 ) ;
 assign wire5657 = ( n_n6  &  wire73 ) | ( n_n6  &  n_n12 ) | ( n_n6  &  wire19469 ) ;
 assign wire5660 = ( n_n4  &  wire166 ) | ( n_n4  &  n_n225  &  wire908 ) ;
 assign wire5661 = ( n_n94  &  wire50 ) | ( n_n281  &  wire903  &  n_n94 ) ;
 assign wire5681 = ( n_n4  &  wire153 ) | ( n_n4  &  wire180 ) ;
 assign wire5699 = ( n_n1  &  wire70 ) | ( n_n228  &  n_n1  &  wire902 ) ;
 assign wire5709 = ( n_n2  &  wire70 ) | ( n_n2  &  wire44 ) ;
 assign wire5743 = ( n_n4  &  wire137 ) | ( n_n4  &  wire132 ) ;
 assign wire5749 = ( n_n1  &  wire137 ) | ( n_n1  &  wire132 ) ;
 assign wire5754 = ( n_n4  &  wire88 ) | ( n_n4  &  n_n222  &  wire908 ) ;
 assign wire5775 = ( n_n3  &  n_n93 ) | ( n_n3  &  wire81 ) | ( n_n3  &  wire76 ) ;
 assign wire5778 = ( n_n268  &  n_n7 ) | ( n_n268  &  wire50 ) | ( n_n268  &  wire119 ) ;
 assign wire5797 = ( n_n139  &  wire48 ) | ( n_n139  &  wire913  &  n_n220 ) ;
 assign wire5812 = ( i_7_  &  i_6_  &  n_n260  &  n_n118 ) | ( i_7_  &  (~ i_6_)  &  n_n260  &  n_n118 ) ;
 assign wire5813 = ( i_7_  &  i_6_  &  n_n118  &  n_n230 ) | ( (~ i_7_)  &  i_6_  &  n_n118  &  n_n230 ) | ( i_7_  &  (~ i_6_)  &  n_n118  &  n_n230 ) ;
 assign wire19350 = ( i_5_  &  (~ i_6_)  &  (~ i_3_)  &  (~ i_4_) ) ;
 assign wire5824 = ( i_1_  &  (~ i_2_)  &  (~ i_0_)  &  wire19350 ) ;
 assign wire19344 = ( wire352 ) | ( n_n281  &  wire914 ) | ( n_n281  &  wire905 ) ;
 assign wire19347 = ( wire215 ) | ( wire152  &  wire1501 ) ;
 assign wire19348 = ( wire19345 ) | ( n_n281  &  wire911 ) | ( n_n281  &  wire912 ) ;
 assign wire19342 = ( wire287 ) | ( n_n281  &  wire901 ) ;
 assign wire19237 = ( i_12_  &  n_n247 ) | ( i_14_  &  i_13_  &  (~ i_12_)  &  n_n247 ) ;
 assign wire5848 = ( n_n128  &  n_n147 ) | ( n_n128  &  wire328 ) | ( n_n128  &  wire19237 ) ;
 assign wire19334 = ( n_n222  &  n_n247 ) | ( n_n247  &  _34585 ) ;
 assign wire5850 = ( n_n165  &  n_n266  &  n_n230 ) ;
 assign wire19332 = ( n_n222  &  n_n259 ) | ( n_n259  &  _34637 ) ;
 assign wire5854 = ( wire72  &  n_n127 ) | ( n_n127  &  wire352 ) | ( n_n127  &  wire19332 ) ;
 assign wire19329 = ( wire214 ) | ( wire19311 ) | ( _34627 ) ;
 assign wire19330 = ( n_n179 ) | ( wire19253 ) | ( wire19326 ) | ( wire19327 ) ;
 assign wire5861 = ( n_n130  &  wire19329 ) | ( n_n130  &  wire19330 ) ;
 assign wire5862 = ( n_n165  &  n_n208  &  n_n230 ) ;
 assign wire19244 = ( i_12_  &  n_n242 ) | ( i_14_  &  i_13_  &  (~ i_12_)  &  n_n242 ) ;
 assign wire5863 = ( n_n124  &  n_n150 ) | ( n_n124  &  wire326 ) | ( n_n124  &  wire19244 ) ;
 assign wire19313 = ( _34558 ) | ( wire913  &  n_n281 ) ;
 assign wire5877 = ( n_n284  &  n_n285  &  n_n271  &  wire1186 ) ;
 assign wire5878 = ( n_n284  &  n_n285  &  n_n266  &  wire1187 ) ;
 assign wire5879 = ( n_n285  &  n_n263  &  _34819 ) ;
 assign wire5880 = ( n_n285  &  n_n261  &  _34822 ) ;
 assign wire19220 = ( n_n247 ) | ( wire911  &  n_n258 ) ;
 assign wire19221 = ( n_n242  &  wire148 ) | ( n_n270  &  wire1135 ) ;
 assign wire19211 = ( n_n242  &  n_n225 ) | ( i_15_  &  n_n242  &  n_n279 ) ;
 assign wire5900 = ( n_n207  &  wire19211 ) | ( wire911  &  n_n228  &  n_n207 ) ;
 assign wire19197 = ( i_9_ ) | ( wire907  &  n_n258 ) ;
 assign wire19198 = ( i_11_  &  n_n163  &  wire148 ) | ( (~ i_11_)  &  n_n163  &  wire971 ) ;
 assign wire19252 = ( _34692 ) | ( n_n281  &  wire905 ) ;
 assign wire5953 = ( n_n132  &  n_n223 ) | ( n_n132  &  wire214 ) | ( n_n132  &  wire19252 ) ;
 assign wire5955 = ( n_n139  &  n_n150 ) | ( n_n139  &  wire326 ) | ( n_n139  &  wire19244 ) ;
 assign wire5973 = ( i_6_  &  n_n165  &  wire19296 ) | ( i_7_  &  (~ i_6_)  &  n_n165  &  wire19296 ) ;
 assign wire5985 = ( n_n285  &  n_n230  &  _34843 ) ;
 assign wire19291 = ( i_7_  &  i_6_  &  (~ i_4_) ) ;
 assign wire5990 = ( n_n285  &  n_n283  &  n_n230  &  wire1223 ) ;
 assign wire5999 = ( (~ i_9_)  &  i_10_  &  i_12_  &  i_11_ ) | ( (~ i_9_)  &  (~ i_10_)  &  i_12_  &  i_11_ ) | ( (~ i_9_)  &  (~ i_10_)  &  i_12_  &  (~ i_11_) ) ;
 assign wire6008 = ( n_n207  &  _34910 ) | ( (~ n_n254)  &  n_n207  &  _34908 ) ;
 assign wire6014 = ( i_13_  &  (~ i_12_)  &  _34914 ) | ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  _34914 ) ;
 assign wire19274 = ( n_n143 ) | ( n_n281  &  n_n253 ) ;
 assign wire19275 = ( n_n279  &  wire898 ) | ( n_n279  &  wire899 ) ;
 assign wire6009 = ( n_n189  &  wire6014 ) | ( n_n189  &  wire19274 ) | ( n_n189  &  wire19275 ) ;
 assign wire19212 = ( (~ i_9_)  &  i_10_  &  i_11_ ) | ( (~ i_9_)  &  (~ i_10_)  &  (~ i_11_) ) ;
 assign wire19228 = ( wire5877 ) | ( wire5878 ) | ( wire5879 ) | ( wire5880 ) ;
 assign wire19233 = ( i_9_  &  i_10_ ) | ( (~ i_9_)  &  i_10_  &  (~ i_11_)  &  n_n279 ) ;
 assign wire19243 = ( _6821 ) | ( _6822 ) | ( wire326  &  _34713 ) ;
 assign wire19250 = ( wire5955 ) | ( _6812 ) | ( _6813 ) ;
 assign wire19254 = ( (~ i_9_)  &  (~ i_10_) ) | ( (~ i_9_)  &  i_10_  &  i_11_ ) ;
 assign wire19255 = ( wire19254 ) | ( n_n281  &  wire914 ) ;
 assign wire19264 = ( i_9_  &  i_10_  &  i_11_ ) | ( (~ i_9_)  &  (~ i_10_)  &  (~ i_11_) ) ;
 assign wire19278 = ( n_n207  &  wire1071 ) | ( n_n207  &  wire1181 ) ;
 assign wire19286 = ( n_n149 ) | ( wire911  &  n_n279 ) ;
 assign wire19287 = ( n_n279  &  wire900 ) | ( wire197  &  wire1225 ) ;
 assign wire19297 = ( wire5985 ) | ( i_9_  &  i_10_  &  wire1265 ) | ( (~ i_9_)  &  (~ i_10_)  &  wire1265 ) ;
 assign wire19299 = ( i_7_  &  i_8_  &  (~ i_6_) ) | ( i_7_  &  (~ i_8_)  &  (~ i_6_)  &  wire1317 ) ;
 assign wire19300 = ( (~ i_7_)  &  (~ i_6_) ) | ( (~ i_7_)  &  i_8_  &  i_6_ ) | ( (~ i_7_)  &  (~ i_8_)  &  i_6_  &  wire315 ) ;
 assign wire19301 = ( i_1_  &  (~ i_2_)  &  (~ i_0_)  &  _34860 ) ;
 assign wire19302 = ( wire5973 ) | ( wire19299  &  wire19301 ) | ( wire19300  &  wire19301 ) ;
 assign wire19303 = ( wire19297 ) | ( wire19302 ) | ( wire315  &  wire1264 ) ;
 assign wire19305 = ( n_n5017 ) | ( wire6008 ) | ( wire6009 ) | ( wire19278 ) ;
 assign wire19307 = ( (~ i_9_)  &  (~ i_10_) ) | ( n_n279  &  wire912 ) ;
 assign wire19311 = ( n_n242  &  n_n222 ) | ( i_15_  &  n_n242  &  n_n279 ) ;
 assign wire19318 = ( i_9_  &  i_10_ ) | ( (~ i_9_)  &  i_10_  &  i_11_ ) | ( (~ i_9_)  &  i_10_  &  i_12_  &  (~ i_11_) ) ;
 assign wire19323 = ( wire5863 ) | ( n_n126  &  wire1400 ) ;
 assign wire19326 = ( (~ i_9_)  &  i_10_  &  i_11_ ) | ( i_9_  &  (~ i_10_)  &  i_11_ ) | ( (~ i_9_)  &  i_10_  &  i_12_  &  (~ i_11_) ) | ( i_9_  &  (~ i_10_)  &  i_12_  &  (~ i_11_) ) ;
 assign wire19327 = ( wire352 ) | ( wire913  &  n_n281 ) | ( n_n281  &  wire914 ) ;
 assign wire19331 = ( wire5862 ) | ( _6927 ) | ( _6928 ) ;
 assign wire19339 = ( wire5848 ) | ( wire5854 ) | ( _34645 ) ;
 assign wire19345 = ( i_9_  &  i_10_ ) | ( i_9_  &  (~ i_10_)  &  i_11_ ) | ( i_9_  &  (~ i_10_)  &  i_12_  &  (~ i_11_) ) ;
 assign wire19353 = ( i_6_  &  n_n230 ) | ( i_7_  &  i_6_  &  n_n260 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n260 ) | ( i_7_  &  (~ i_6_)  &  n_n230 ) ;
 assign wire19354 = ( (~ i_6_)  &  n_n264 ) | ( (~ i_7_)  &  i_6_  &  n_n264 ) | ( i_7_  &  i_6_  &  n_n284 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n284 ) ;
 assign wire19355 = ( wire5824 ) | ( n_n120  &  wire19353 ) | ( n_n120  &  wire19354 ) ;
 assign wire19363 = ( wire5812 ) | ( wire289  &  n_n118  &  n_n230 ) ;
 assign wire19364 = ( n_n5664 ) | ( n_n5679 ) | ( wire587 ) ;
 assign wire19369 = ( n_n5686 ) | ( wire394 ) | ( n_n151  &  wire937 ) ;
 assign wire19377 = ( n_n54  &  n_n100 ) | ( n_n241  &  n_n103 ) ;
 assign wire19379 = ( wire372 ) | ( wire386 ) ;
 assign wire19383 = ( n_n4  &  n_n95 ) | ( n_n4  &  n_n49 ) | ( n_n4  &  wire71 ) ;
 assign wire19394 = ( n_n228  &  wire902 ) | ( n_n281  &  wire903 ) ;
 assign wire19402 = ( n_n228  &  wire902 ) | ( n_n281  &  wire903 ) ;
 assign wire19422 = ( _6160 ) | ( _6161 ) | ( _35504 ) | ( _35505 ) ;
 assign wire19442 = ( n_n3  &  n_n95 ) | ( n_n3  &  n_n49 ) | ( n_n3  &  wire99 ) ;
 assign wire19443 = ( n_n4  &  n_n12 ) | ( n_n3  &  n_n15 ) ;
 assign wire19447 = ( n_n228  &  n_n4  &  wire902 ) | ( n_n228  &  wire902  &  n_n53 ) ;
 assign wire19452 = ( wire634 ) | ( _6252 ) | ( n_n1  &  wire68 ) ;
 assign wire19453 = ( n_n3791 ) | ( n_n2274 ) | ( n_n639 ) | ( wire19447 ) ;
 assign wire19460 = ( n_n4  &  n_n93 ) | ( n_n94  &  n_n24 ) ;
 assign wire19461 = ( n_n4  &  n_n76 ) | ( n_n4  &  n_n26 ) | ( n_n4  &  n_n30 ) ;
 assign wire19470 = ( n_n5  &  wire70 ) | ( n_n5  &  n_n66 ) | ( n_n5  &  n_n14 ) ;
 assign wire19475 = ( n_n9  &  n_n227 ) | ( n_n9  &  n_n207 ) | ( n_n227  &  n_n59 ) | ( n_n207  &  n_n59 ) ;
 assign wire19478 = ( n_n3803 ) | ( wire5640 ) | ( wire5642 ) ;
 assign wire19499 = ( n_n220  &  wire908  &  n_n53 ) | ( wire908  &  n_n256  &  n_n53 ) ;
 assign wire19502 = ( wire478 ) | ( wire19499 ) | ( _6474 ) ;
 assign wire19515 = ( wire5591 ) | ( wire5592 ) | ( n_n9  &  n_n57 ) ;
 assign wire19516 = ( wire571 ) | ( wire737 ) | ( n_n53  &  wire68 ) ;
 assign wire19519 = ( wire5589 ) | ( wire19516 ) | ( n_n57  &  n_n12 ) ;
 assign wire19520 = ( n_n4381 ) | ( n_n3850 ) | ( wire5577 ) | ( wire19515 ) ;
 assign wire19522 = ( wire869 ) | ( _6408 ) | ( n_n48  &  _35208 ) ;
 assign wire19526 = ( n_n5  &  wire255 ) | ( n_n5  &  wire190 ) ;
 assign wire19528 = ( n_n4770 ) | ( wire19526 ) | ( n_n6  &  wire1747 ) ;
 assign wire19534 = ( n_n4675 ) | ( n_n4676 ) | ( _6058 ) ;
 assign wire19539 = ( n_n57  &  wire70 ) | ( n_n56  &  n_n76 ) ;
 assign wire19541 = ( n_n4924 ) | ( wire788 ) | ( wire5544 ) ;
 assign wire19549 = ( n_n100  &  n_n103 ) | ( n_n94  &  n_n75 ) ;
 assign wire19550 = ( n_n74  &  n_n94 ) | ( n_n94  &  n_n24 ) | ( n_n94  &  wire77 ) ;
 assign wire19559 = ( n_n60  &  n_n100 ) | ( n_n9  &  n_n100 ) | ( wire63  &  n_n100 ) ;
 assign wire19568 = ( wire40  &  n_n100 ) | ( n_n228  &  wire898  &  n_n100 ) ;
 assign wire19571 = ( _5980 ) | ( _5981 ) | ( _5982 ) ;
 assign wire19588 = ( wire19380 ) | ( n_n3661 ) | ( _35648 ) | ( _35724 ) ;
 assign wire19599 = ( wire364 ) | ( wire777 ) | ( wire834 ) ;
 assign wire19609 = ( _35772 ) | ( wire48  &  n_n124 ) ;
 assign wire19617 = ( n_n5678 ) | ( n_n5671 ) | ( wire396  &  wire940 ) ;
 assign wire19619 = ( wire5453 ) | ( wire19613 ) | ( wire19614 ) | ( wire19617 ) ;
 assign wire19620 = ( wire582 ) | ( wire5445 ) | ( n_n106  &  wire941 ) ;
 assign wire19628 = ( i_7_  &  i_6_  &  n_n260  &  n_n116 ) | ( i_7_  &  (~ i_6_)  &  n_n260  &  n_n116 ) ;
 assign wire19631 = ( wire793 ) | ( wire19628 ) ;
 assign wire19632 = ( wire880 ) | ( n_n5672 ) | ( _35855 ) ;
 assign wire19633 = ( n_n139  &  n_n111 ) | ( wire54  &  n_n132 ) ;
 assign wire19636 = ( n_n111  &  n_n121 ) | ( n_n111  &  n_n132 ) | ( n_n111  &  n_n122 ) ;
 assign wire19642 = ( n_n5671 ) | ( wire5412 ) | ( wire5413 ) ;
 assign wire19644 = ( wire5411 ) | ( wire19631 ) | ( wire19632 ) | ( wire19642 ) ;
 assign wire19645 = ( wire5426 ) | ( wire5430 ) | ( wire19633 ) | ( wire19636 ) ;
 assign wire19665 = ( n_n4870 ) | ( _5593 ) | ( n_n6  &  _36101 ) ;
 assign wire19669 = ( n_n220  &  n_n6  &  wire904 ) | ( n_n6  &  n_n256  &  wire904 ) ;
 assign wire19696 = ( n_n3324 ) | ( n_n4381 ) | ( wire5587 ) | ( wire5588 ) ;
 assign wire19701 = ( wire268  &  n_n57 ) | ( n_n57  &  wire198 ) ;
 assign wire19703 = ( n_n4941 ) | ( n_n4942 ) | ( wire762 ) ;
 assign wire19704 = ( wire728 ) | ( wire19701 ) | ( n_n57  &  wire167 ) ;
 assign wire19705 = ( n_n56  &  wire190 ) | ( n_n57  &  wire124 ) ;
 assign wire19706 = ( n_n56  &  wire124 ) | ( n_n57  &  wire212 ) ;
 assign wire19707 = ( n_n56  &  wire212 ) | ( n_n57  &  wire119 ) ;
 assign wire19709 = ( wire19705 ) | ( wire19706 ) ;
 assign wire19710 = ( wire761 ) | ( wire19707 ) | ( n_n56  &  wire198 ) ;
 assign wire19720 = ( n_n57  &  wire180 ) | ( n_n56  &  wire254 ) ;
 assign wire19724 = ( n_n4954 ) | ( n_n4953 ) | ( n_n4955 ) | ( wire671 ) ;
 assign wire19725 = ( wire200  &  n_n57 ) | ( n_n56  &  wire277 ) ;
 assign wire19728 = ( wire729 ) | ( wire19725 ) | ( wire268  &  n_n56 ) ;
 assign wire19730 = ( n_n56  &  wire224 ) | ( n_n56  &  wire180 ) ;
 assign wire19732 = ( n_n4970 ) | ( wire614 ) | ( n_n56  &  wire166 ) ;
 assign wire19735 = ( wire19724 ) | ( wire19728 ) | ( _36064 ) ;
 assign wire19747 = ( n_n4834 ) | ( n_n4839 ) | ( _5552 ) ;
 assign wire19755 = ( wire5238 ) | ( wire5242 ) | ( _36219 ) ;
 assign wire19757 = ( wire19754 ) | ( n_n4858 ) | ( n_n4864 ) | ( _5485 ) ;
 assign wire19759 = ( n_n4807 ) | ( n_n4806 ) | ( wire72  &  n_n5 ) ;
 assign wire19761 = ( n_n4223 ) | ( n_n4224 ) | ( wire19759 ) ;
 assign wire19780 = ( n_n106  &  n_n2 ) | ( n_n2  &  n_n62 ) | ( n_n2  &  wire101 ) ;
 assign wire19791 = ( wire5184 ) | ( wire5709 ) | ( n_n1  &  n_n12 ) ;
 assign wire19807 = ( n_n106  &  n_n2 ) | ( n_n1  &  wire68 ) ;
 assign wire19808 = ( wire19807 ) | ( n_n2  &  wire200 ) | ( n_n2  &  wire112 ) ;
 assign wire19810 = ( wire19808 ) | ( _5381 ) | ( _5389 ) | ( _36298 ) ;
 assign wire19812 = ( wire19798 ) | ( n_n2582 ) | ( wire19810 ) | ( _36289 ) ;
 assign wire19821 = ( n_n2618 ) | ( _5365 ) | ( _36311 ) ;
 assign wire19825 = ( wire758 ) | ( n_n220  &  wire914  &  n_n122 ) ;
 assign wire19826 = ( n_n5678 ) | ( n_n5671 ) | ( wire5144 ) ;
 assign wire19830 = ( wire582 ) | ( wire19826 ) | ( _5341 ) ;
 assign wire19837 = ( n_n5769 ) | ( wire48  &  n_n127 ) ;
 assign wire19842 = ( n_n207  &  _36341 ) | ( wire905  &  n_n207  &  _36337 ) ;
 assign wire19843 = ( n_n9  &  n_n227 ) | ( n_n227  &  n_n59 ) | ( n_n207  &  n_n59 ) ;
 assign wire19854 = ( n_n268  &  wire247 ) | ( n_n265  &  wire277 ) ;
 assign wire19857 = ( n_n265  &  wire268 ) | ( n_n265  &  wire200 ) | ( n_n265  &  wire112 ) ;
 assign wire19859 = ( wire19857 ) | ( _5282 ) | ( _5283 ) ;
 assign wire19862 = ( n_n5796 ) | ( wire914  &  n_n6  &  n_n256 ) ;
 assign wire19867 = ( n_n6  &  wire153 ) | ( n_n6  &  wire57 ) | ( n_n6  &  n_n113 ) ;
 assign wire19868 = ( wire617 ) | ( wire5091 ) | ( n_n5  &  wire255 ) ;
 assign wire19872 = ( n_n4770 ) | ( n_n4773 ) | ( wire19867 ) | ( _36550 ) ;
 assign wire19888 = ( wire541 ) | ( n_n4815 ) | ( n_n4814 ) | ( n_n4816 ) ;
 assign wire19904 = ( n_n4846 ) | ( n_n4852 ) | ( wire5242 ) | ( wire5243 ) ;
 assign wire19906 = ( wire19904 ) | ( _36506 ) ;
 assign wire19916 = ( n_n57  &  n_n11 ) | ( n_n56  &  n_n11 ) | ( n_n57  &  wire113 ) ;
 assign wire19918 = ( wire5589 ) | ( wire5013 ) | ( wire5014 ) | ( wire5590 ) ;
 assign wire19919 = ( n_n4895 ) | ( wire5002 ) | ( wire19916 ) ;
 assign wire19921 = ( wire5011 ) | ( wire5012 ) | ( wire19918 ) | ( wire19919 ) ;
 assign wire19925 = ( wire273  &  n_n56 ) | ( wire268  &  n_n56 ) | ( n_n56  &  wire157 ) ;
 assign wire19926 = ( n_n4941 ) | ( n_n4942 ) | ( wire729 ) ;
 assign wire19927 = ( wire19925 ) | ( wire268  &  n_n57 ) | ( wire200  &  n_n57 ) ;
 assign wire19928 = ( n_n56  &  wire124 ) | ( n_n56  &  wire212 ) ;
 assign wire19938 = ( n_n5796 ) | ( n_n56  &  wire49 ) ;
 assign wire19941 = ( n_n57  &  wire124 ) | ( n_n57  &  wire212 ) ;
 assign wire19943 = ( n_n4926 ) | ( n_n4923 ) | ( wire19938 ) ;
 assign wire19944 = ( n_n4924 ) | ( n_n4922 ) | ( wire19941 ) ;
 assign wire19952 = ( n_n57  &  wire99 ) | ( n_n57  &  wire41 ) ;
 assign wire19958 = ( wire394 ) | ( n_n139  &  wire48 ) | ( wire48  &  n_n132 ) ;
 assign wire19965 = ( n_n5686 ) | ( n_n5693 ) | ( wire609 ) | ( wire4947 ) ;
 assign wire19971 = ( n_n57  &  wire180 ) | ( n_n56  &  wire254 ) ;
 assign wire19973 = ( _36461 ) | ( n_n57  &  wire153 ) | ( n_n57  &  wire166 ) ;
 assign wire19974 = ( wire4939 ) | ( wire19971 ) | ( n_n57  &  wire224 ) ;
 assign wire19977 = ( wire200  &  n_n56 ) | ( wire112  &  n_n56 ) | ( n_n56  &  wire99 ) ;
 assign wire19984 = ( n_n5796 ) | ( n_n6  &  wire75 ) | ( n_n6  &  n_n206 ) ;
 assign wire19986 = ( n_n4806 ) | ( wire19984 ) | ( wire72  &  n_n5 ) ;
 assign wire19987 = ( n_n4808 ) | ( n_n4809 ) | ( wire19986 ) ;
 assign wire19996 = ( i_3_  &  n_n116 ) | ( n_n116  &  n_n155  &  n_n230 ) ;
 assign wire19997 = ( i_7_  &  i_6_  &  n_n260  &  n_n116 ) | ( (~ i_7_)  &  i_6_  &  n_n260  &  n_n116 ) | ( i_7_  &  (~ i_6_)  &  n_n260  &  n_n116 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n260  &  n_n116 ) ;
 assign wire19999 = ( (~ i_7_)  &  i_6_  &  n_n118  &  n_n230 ) | ( i_7_  &  (~ i_6_)  &  n_n118  &  n_n230 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n118  &  n_n230 ) ;
 assign wire20000 = ( i_3_  &  n_n118 ) | ( n_n260  &  n_n118  &  n_n155 ) ;
 assign wire20011 = ( n_n111  &  n_n130 ) | ( n_n111  &  n_n121 ) | ( n_n130  &  wire948 ) ;
 assign wire20015 = ( n_n139  &  n_n110 ) | ( wire48  &  n_n132 ) ;
 assign wire20016 = ( wire4900 ) | ( n_n139  &  wire48 ) ;
 assign wire20017 = ( wire48  &  n_n130 ) | ( n_n110  &  n_n132 ) ;
 assign wire20028 = ( n_n264  &  n_n116  &  n_n155 ) | ( n_n260  &  n_n116  &  n_n155 ) ;
 assign wire20030 = ( wire581 ) | ( wire794 ) ;
 assign wire20031 = ( n_n5685 ) | ( wire4871 ) | ( wire20028 ) ;
 assign wire20038 = ( n_n10  &  n_n100 ) | ( n_n100  &  n_n63 ) | ( n_n100  &  n_n62 ) ;
 assign wire20041 = ( n_n2702 ) | ( wire654 ) | ( _4861 ) ;
 assign wire20042 = ( wire4856 ) | ( wire4869 ) | ( wire4870 ) | ( wire20038 ) ;
 assign wire20045 = ( n_n133  &  n_n94 ) | ( n_n94  &  n_n17 ) | ( n_n94  &  n_n68 ) ;
 assign wire20047 = ( n_n2732 ) | ( n_n2398 ) | ( wire20045 ) ;
 assign wire20048 = ( wire4849 ) | ( n_n100  &  wire1150 ) ;
 assign wire20054 = ( wire4844 ) | ( wire4845 ) | ( _36824 ) ;
 assign wire20055 = ( wire20041 ) | ( wire20042 ) | ( wire20047 ) | ( wire20048 ) ;
 assign wire20066 = ( n_n216  &  n_n94 ) | ( n_n204  &  n_n94 ) | ( n_n94  &  n_n203 ) ;
 assign wire20070 = ( n_n74  &  n_n94 ) | ( n_n94  &  n_n75 ) | ( n_n94  &  n_n24 ) ;
 assign wire20072 = ( n_n707 ) | ( wire4817 ) | ( wire20070 ) ;
 assign wire20081 = ( n_n37  &  n_n100 ) | ( n_n104  &  n_n100 ) | ( n_n100  &  n_n84 ) ;
 assign wire20084 = ( wire4807 ) | ( wire4808 ) ;
 assign wire20088 = ( _4906 ) | ( _4907 ) | ( _4908 ) ;
 assign wire20099 = ( n_n104  &  n_n100 ) | ( n_n110  &  n_n94 ) ;
 assign wire20100 = ( n_n100  &  n_n84 ) | ( n_n94  &  n_n68 ) ;
 assign wire20101 = ( n_n133  &  n_n94 ) | ( n_n16  &  n_n94 ) | ( n_n94  &  n_n22 ) ;
 assign wire20108 = ( n_n10  &  n_n100 ) | ( n_n147  &  n_n94 ) ;
 assign wire20111 = ( wire4766 ) | ( wire20108 ) | ( n_n100  &  n_n63 ) ;
 assign wire20113 = ( n_n2702 ) | ( wire687 ) | ( n_n2671 ) | ( wire20111 ) ;
 assign wire20137 = ( n_n5  &  wire67 ) | ( n_n5  &  wire912  &  n_n258 ) ;
 assign wire20174 = ( n_n6  &  n_n226 ) | ( n_n5  &  wire208 ) ;
 assign wire20186 = ( i_7_  &  i_6_  &  n_n260  &  n_n116 ) | ( (~ i_7_)  &  i_6_  &  n_n260  &  n_n116 ) ;
 assign wire20188 = ( i_7_  &  i_6_  &  n_n116  &  n_n230 ) | ( (~ i_7_)  &  i_6_  &  n_n116  &  n_n230 ) ;
 assign wire20190 = ( n_n5673 ) | ( n_n5675 ) | ( wire20188 ) ;
 assign wire20191 = ( n_n5677 ) | ( wire20186 ) | ( n_n128  &  wire371 ) ;
 assign wire20193 = ( n_n111  &  n_n56 ) | ( n_n56  &  wire453 ) | ( n_n56  &  n_n38 ) ;
 assign wire20203 = ( n_n57  &  n_n32 ) | ( n_n56  &  n_n32 ) | ( n_n57  &  wire85 ) ;
 assign wire20206 = ( wire460 ) | ( n_n4666 ) | ( wire20193 ) | ( wire20203 ) ;
 assign wire20212 = ( wire826 ) | ( n_n54  &  n_n57 ) | ( n_n57  &  n_n99 ) ;
 assign wire20216 = ( n_n4687 ) | ( n_n4686 ) | ( wire4641 ) | ( wire20212 ) ;
 assign wire20227 = ( n_n4923 ) | ( _4769 ) ;
 assign wire20236 = ( n_n5671 ) | ( n_n5659 ) | ( wire4618 ) ;
 assign wire20238 = ( wire4617 ) | ( wire20190 ) | ( wire20191 ) | ( wire20236 ) ;
 assign wire20248 = ( wire912  &  n_n258  &  n_n48 ) | ( wire912  &  n_n256  &  n_n48 ) ;
 assign wire20264 = ( n_n258  &  n_n48  &  wire897 ) | ( n_n258  &  n_n53  &  wire897 ) ;
 assign wire20265 = ( n_n53  &  n_n76 ) | ( n_n53  &  n_n26 ) | ( n_n53  &  n_n78 ) ;
 assign wire20268 = ( wire478 ) | ( wire20265 ) | ( n_n48  &  wire40 ) ;
 assign wire20269 = ( wire20264 ) | ( _4456 ) | ( _4457 ) ;
 assign wire20277 = ( n_n53  &  _37161 ) | ( wire908  &  n_n53  &  _35046 ) ;
 assign wire20278 = ( n_n53  &  n_n10 ) | ( n_n48  &  n_n148 ) ;
 assign wire20279 = ( n_n246  &  n_n48 ) | ( n_n11  &  n_n48 ) | ( n_n48  &  n_n147 ) ;
 assign wire20285 = ( wire911  &  n_n258  &  n_n48 ) | ( n_n258  &  wire899  &  n_n48 ) ;
 assign wire20299 = ( wire571 ) | ( n_n258  &  wire900  &  n_n48 ) ;
 assign wire20307 = ( n_n220  &  wire907 ) | ( wire907  &  n_n256 ) | ( n_n220  &  wire904 ) | ( n_n256  &  wire904 ) ;
 assign wire20323 = ( n_n11  &  n_n48 ) | ( n_n53  &  n_n63 ) ;
 assign wire20324 = ( n_n246  &  n_n48 ) | ( n_n53  &  n_n10 ) ;
 assign wire20325 = ( n_n106  &  n_n53 ) | ( n_n48  &  n_n86 ) ;
 assign wire20334 = ( n_n48  &  _37244 ) | ( wire899  &  n_n48  &  _37091 ) ;
 assign wire20336 = ( n_n53  &  _37247 ) | ( wire899  &  n_n53  &  _37091 ) ;
 assign wire20337 = ( n_n257  &  n_n53 ) | ( n_n145  &  n_n53 ) | ( n_n53  &  n_n144 ) ;
 assign wire20343 = ( n_n70  &  n_n53 ) | ( n_n53  &  n_n107 ) | ( n_n53  &  n_n19 ) ;
 assign wire20346 = ( n_n60  &  n_n53 ) | ( n_n48  &  n_n148 ) ;
 assign wire20347 = ( n_n226  &  n_n53 ) | ( n_n257  &  n_n53 ) | ( n_n108  &  n_n53 ) ;
 assign wire20349 = ( n_n4068 ) | ( wire20347 ) ;
 assign wire20350 = ( wire626 ) | ( n_n1433 ) | ( wire20343 ) | ( wire20346 ) ;
 assign wire20356 = ( n_n6  &  n_n60 ) | ( n_n6  &  n_n9 ) | ( n_n6  &  wire63 ) ;
 assign wire20369 = ( n_n4  &  n_n31 ) | ( n_n10  &  n_n100 ) ;
 assign wire20370 = ( n_n228  &  wire901  &  n_n100 ) | ( n_n279  &  wire901  &  n_n100 ) ;
 assign wire20371 = ( n_n106  &  n_n100 ) | ( n_n100  &  n_n33 ) | ( n_n100  &  n_n81 ) ;
 assign wire20379 = ( n_n6  &  wire75 ) | ( n_n6  &  n_n206 ) | ( n_n6  &  n_n226 ) ;
 assign wire20390 = ( n_n257  &  n_n53 ) | ( n_n1  &  wire68 ) ;
 assign wire20401 = ( n_n4  &  n_n105 ) | ( n_n4  &  n_n108 ) | ( n_n4  &  n_n70 ) ;
 assign wire20404 = ( n_n4  &  _37499 ) | ( n_n4  &  wire906  &  _35394 ) ;
 assign wire20408 = ( _37496 ) | ( n_n4  &  n_n9 ) | ( n_n4  &  _37495 ) ;
 assign wire20409 = ( wire446 ) | ( n_n2982 ) | ( wire20404 ) ;
 assign wire20418 = ( n_n53  &  _37340 ) | ( wire914  &  n_n53  &  _34565 ) ;
 assign wire20419 = ( n_n53  &  _37341 ) | ( wire907  &  n_n53  &  _36833 ) ;
 assign wire20422 = ( n_n3581 ) | ( n_n4160 ) | ( wire20418 ) | ( wire20419 ) ;
 assign wire20424 = ( wire407 ) | ( n_n228  &  wire902  &  n_n53 ) ;
 assign wire20425 = ( n_n145  &  n_n53 ) | ( n_n53  &  n_n7 ) | ( n_n53  &  n_n144 ) ;
 assign wire20434 = ( n_n6  &  n_n104 ) | ( n_n6  &  wire368 ) | ( n_n6  &  n_n88 ) ;
 assign wire20438 = ( n_n6  &  wire78 ) | ( n_n6  &  wire19457 ) | ( n_n6  &  n_n25 ) ;
 assign wire20444 = ( n_n6  &  n_n54 ) | ( n_n53  &  n_n32 ) ;
 assign wire20445 = ( n_n53  &  _37286 ) | ( wire901  &  n_n53  &  _36817 ) ;
 assign wire20449 = ( wire389 ) | ( wire882 ) | ( wire20444 ) | ( wire20445 ) ;
 assign wire20450 = ( wire670 ) | ( n_n3019 ) | ( wire4423 ) ;
 assign wire20455 = ( n_n37  &  n_n53 ) | ( n_n53  &  n_n104 ) | ( n_n53  &  n_n32 ) ;
 assign wire20460 = ( wire571 ) | ( wire4418 ) ;
 assign wire20461 = ( wire407 ) | ( wire579 ) | ( n_n53  &  wire68 ) ;
 assign wire20463 = ( n_n228  &  wire902 ) | ( n_n281  &  wire903 ) ;
 assign wire20474 = ( _4300 ) | ( _4301 ) | ( _4302 ) ;
 assign wire20479 = ( wire478 ) | ( n_n1433 ) | ( wire20344 ) | ( wire20343 ) ;
 assign wire20480 = ( _4263 ) | ( _4264 ) ;
 assign wire20486 = ( n_n57  &  n_n32 ) | ( n_n57  &  n_n81 ) | ( n_n57  &  wire86 ) ;
 assign wire20492 = ( wire95  &  n_n57 ) | ( n_n57  &  n_n108 ) | ( n_n57  &  n_n11 ) ;
 assign wire20499 = ( n_n57  &  n_n95 ) | ( n_n151  &  n_n100 ) ;
 assign wire20506 = ( n_n100  &  wire83 ) | ( wire911  &  n_n258  &  n_n100 ) ;
 assign wire20510 = ( n_n281  &  wire906 ) | ( n_n228  &  wire901 ) ;
 assign wire20519 = ( n_n100  &  n_n103 ) | ( n_n100  &  wire19457 ) | ( n_n100  &  n_n25 ) ;
 assign wire20520 = ( n_n241  &  n_n258  &  wire901 ) | ( n_n241  &  n_n258  &  wire897 ) ;
 assign wire20522 = ( n_n241  &  n_n105 ) | ( n_n54  &  n_n100 ) ;
 assign wire20525 = ( wire559 ) | ( wire20522 ) | ( n_n177  &  n_n200 ) ;
 assign wire20527 = ( wire912  &  n_n258 ) | ( n_n225  &  wire901 ) ;
 assign wire20536 = ( n_n220  &  wire907  &  n_n100 ) | ( wire907  &  n_n256  &  n_n100 ) ;
 assign wire20537 = ( n_n100  &  wire77 ) | ( n_n258  &  wire900  &  n_n100 ) ;
 assign wire20540 = ( n_n3884 ) | ( wire4330 ) | ( wire20536 ) | ( wire20537 ) ;
 assign wire20549 = ( n_n4922 ) | ( n_n4921 ) | ( wire693 ) ;
 assign wire20581 = ( n_n4  &  n_n108 ) | ( n_n4  &  wire44 ) | ( n_n4  &  n_n65 ) ;
 assign wire20590 = ( wire485 ) | ( n_n3731 ) | ( wire4285 ) | ( _37576 ) ;
 assign wire20593 = ( n_n228  &  wire902 ) | ( n_n281  &  wire903 ) ;
 assign wire20600 = ( _37539 ) | ( n_n1  &  wire63 ) | ( n_n1  &  _35356 ) ;
 assign wire20604 = ( n_n1  &  n_n108 ) | ( n_n1  &  wire84 ) | ( n_n1  &  n_n112 ) ;
 assign wire20606 = ( n_n3524 ) | ( wire468 ) | ( wire20604 ) ;
 assign wire20608 = ( n_n4  &  n_n95 ) | ( n_n265  &  n_n62 ) ;
 assign wire20609 = ( n_n4  &  n_n105 ) | ( n_n4  &  n_n47 ) | ( n_n4  &  wire68 ) ;
 assign wire20620 = ( n_n4  &  n_n12 ) | ( n_n4  &  n_n64 ) | ( n_n4  &  n_n13 ) ;
 assign wire20622 = ( n_n4015 ) | ( wire4248 ) | ( wire20620 ) ;
 assign wire20624 = ( n_n2840 ) | ( n_n2839 ) | ( wire20622 ) ;
 assign wire20633 = ( n_n260  &  n_n118  &  n_n155 ) | ( n_n284  &  n_n118  &  n_n155 ) ;
 assign wire20636 = ( n_n5664 ) | ( n_n272  &  wire930 ) | ( n_n272  &  wire1740 ) ;
 assign wire20641 = ( n_n260  &  n_n116  &  n_n155 ) | ( n_n116  &  n_n284  &  n_n155 ) ;
 assign wire20642 = ( n_n264  &  n_n116  &  n_n155 ) | ( n_n116  &  n_n155  &  n_n230 ) ;
 assign wire20643 = ( n_n260  &  n_n116  &  n_n272 ) | ( n_n116  &  n_n272  &  n_n230 ) ;
 assign wire20646 = ( n_n5676 ) | ( wire20641 ) | ( n_n128  &  wire216 ) ;
 assign wire20655 = ( n_n255  &  n_n197 ) | ( n_n241  &  n_n103 ) ;
 assign wire20668 = ( n_n260  &  n_n165  &  n_n272 ) | ( n_n165  &  n_n284  &  n_n272 ) ;
 assign wire20682 = ( n_n4895 ) | ( wire5013 ) | ( wire5014 ) ;
 assign wire20683 = ( n_n4892 ) | ( n_n4898 ) | ( wire5035 ) | ( wire5036 ) ;
 assign wire20686 = ( n_n4210 ) | ( wire878 ) | ( wire20682 ) | ( wire20683 ) ;
 assign wire20689 = ( n_n4870 ) | ( n_n4871 ) | ( wire4183 ) | ( wire5091 ) ;
 assign wire20692 = ( n_n5796 ) | ( n_n56  &  wire49 ) ;
 assign wire20694 = ( n_n57  &  wire190 ) | ( n_n57  &  wire212 ) ;
 assign wire20695 = ( n_n56  &  wire124 ) | ( n_n56  &  wire212 ) ;
 assign wire20696 = ( n_n57  &  wire119 ) | ( n_n56  &  wire119 ) ;
 assign wire20699 = ( n_n4926 ) | ( n_n4929 ) | ( wire20692 ) | ( wire20696 ) ;
 assign wire20701 = ( n_n56  &  wire224 ) | ( n_n56  &  wire180 ) ;
 assign wire20703 = ( _37673 ) | ( n_n57  &  wire99 ) | ( n_n57  &  wire41 ) ;
 assign wire20704 = ( n_n4967 ) | ( wire613 ) | ( wire20701 ) ;
 assign wire20711 = ( n_n132  &  n_n107 ) | ( n_n139  &  wire250 ) ;
 assign wire20714 = ( n_n5796 ) | ( n_n132  &  wire250 ) ;
 assign wire20716 = ( wire4159 ) | ( wire4170 ) | ( wire20711 ) | ( wire20714 ) ;
 assign wire20728 = ( n_n4923 ) | ( n_n4924 ) | ( wire5544 ) ;
 assign wire20737 = ( wire273  &  n_n56 ) | ( n_n56  &  wire157 ) ;
 assign wire20739 = ( n_n4941 ) | ( n_n4942 ) | ( _37689 ) ;
 assign wire20742 = ( n_n4218 ) | ( wire20694 ) | ( wire20695 ) | ( wire20699 ) ;
 assign wire20745 = ( n_n5796 ) | ( n_n6  &  wire75 ) | ( n_n6  &  n_n206 ) ;
 assign wire20746 = ( n_n4806 ) | ( wire20745 ) | ( wire72  &  n_n5 ) ;
 assign wire20748 = ( n_n4223 ) | ( n_n4224 ) | ( wire20746 ) ;
 assign wire20751 = ( n_n4203 ) | ( n_n4206 ) | ( n_n4211 ) | ( wire20686 ) ;
 assign wire20758 = ( n_n94  &  _37738 ) | ( wire911  &  n_n94  &  _36343 ) ;
 assign wire20759 = ( n_n216  &  n_n100 ) | ( n_n94  &  n_n17 ) ;
 assign wire20760 = ( n_n133  &  n_n94 ) | ( n_n16  &  n_n94 ) | ( n_n94  &  n_n67 ) ;
 assign wire20767 = ( n_n241  &  n_n216 ) | ( n_n255  &  n_n197 ) ;
 assign wire20769 = ( wire20755 ) | ( wire20767 ) | ( n_n54  &  n_n100 ) ;
 assign wire20772 = ( wire44  &  n_n100 ) | ( n_n252  &  n_n100 ) | ( n_n15  &  n_n100 ) ;
 assign wire20776 = ( wire118  &  n_n94 ) | ( n_n145  &  n_n94 ) | ( n_n94  &  n_n144 ) ;
 assign wire20779 = ( wire5514 ) | ( wire5515 ) | ( n_n2713 ) | ( wire4100 ) ;
 assign wire20784 = ( n_n57  &  wire82 ) | ( n_n57  &  wire42 ) | ( n_n57  &  n_n223 ) ;
 assign wire20800 = ( n_n4  &  _37915 ) | ( n_n4  &  wire899  &  _37091 ) ;
 assign wire20802 = ( n_n4005 ) | ( wire446 ) | ( wire20800 ) ;
 assign wire20814 = ( wire557 ) | ( n_n3506 ) | ( wire485 ) | ( wire933 ) ;
 assign wire20817 = ( n_n3417 ) | ( _6235 ) | ( _6236 ) | ( _37932 ) ;
 assign wire20820 = ( n_n110  &  n_n53 ) | ( n_n48  &  wire82 ) ;
 assign wire20824 = ( wire4062 ) | ( wire5625 ) | ( wire5626 ) | ( wire20820 ) ;
 assign wire20826 = ( wire764 ) | ( n_n53  &  wire68 ) ;
 assign wire20827 = ( wire579 ) | ( n_n228  &  n_n57  &  wire899 ) ;
 assign wire20831 = ( wire406 ) | ( wire4044 ) | ( n_n95  &  n_n48 ) ;
 assign wire20832 = ( wire309 ) | ( wire4056 ) | ( wire20826 ) | ( wire20827 ) ;
 assign wire20833 = ( n_n1433 ) | ( n_n3587 ) | ( wire5589 ) | ( wire5590 ) ;
 assign wire20842 = ( wire411 ) | ( wire4036 ) | ( n_n5  &  wire255 ) ;
 assign wire20847 = ( n_n70  &  n_n53 ) | ( n_n53  &  n_n107 ) | ( n_n53  &  n_n19 ) ;
 assign wire20851 = ( n_n53  &  _37841 ) | ( wire899  &  n_n53  &  _37091 ) ;
 assign wire20853 = ( n_n4154 ) | ( wire475 ) | ( wire20851 ) ;
 assign wire20854 = ( wire4016 ) | ( wire4520 ) | ( wire20334 ) ;
 assign wire20856 = ( wire5613 ) | ( wire20853 ) | ( wire20854 ) | ( _35030 ) ;
 assign wire20876 = ( wire72  &  n_n5 ) | ( n_n257  &  n_n207 ) ;
 assign wire20883 = ( n_n4  &  n_n93 ) | ( n_n110  &  n_n94 ) ;
 assign wire20894 = ( wire639 ) | ( wire3967 ) | ( wire5656 ) | ( wire5657 ) ;
 assign wire20895 = ( n_n4809 ) | ( wire539 ) | ( wire3968 ) | ( wire20894 ) ;
 assign wire20898 = ( n_n4  &  n_n257 ) | ( n_n53  &  n_n107 ) ;
 assign wire20899 = ( n_n228  &  wire899  &  n_n53 ) | ( wire899  &  n_n256  &  n_n53 ) ;
 assign wire20900 = ( n_n145  &  n_n53 ) | ( n_n53  &  n_n144 ) | ( n_n53  &  n_n71 ) ;
 assign wire20907 = ( n_n4  &  n_n226 ) | ( n_n4  &  n_n145 ) | ( n_n4  &  n_n144 ) ;
 assign wire20908 = ( wire409 ) | ( wire546 ) | ( wire19443 ) | ( wire20907 ) ;
 assign wire20909 = ( wire5681 ) | ( wire19442 ) | ( _37951 ) ;
 assign wire20912 = ( n_n3382 ) | ( n_n3383 ) | ( wire20908 ) | ( wire20909 ) ;
 assign wire20942 = ( _3294 ) | ( _3295 ) ;
 assign wire20952 = ( n_n6  &  _38125 ) | ( n_n6  &  wire899  &  _37091 ) ;
 assign wire20967 = ( n_n1  &  n_n95 ) | ( n_n2  &  wire68 ) ;
 assign wire20981 = ( n_n94  &  n_n41 ) | ( n_n227  &  n_n28 ) ;
 assign wire20982 = ( n_n5  &  n_n145 ) | ( n_n70  &  n_n227 ) ;
 assign wire20988 = ( n_n4  &  n_n9 ) | ( n_n3  &  n_n66 ) ;
 assign wire20989 = ( n_n4  &  n_n61 ) | ( n_n3  &  n_n15 ) ;
 assign wire20993 = ( wire446 ) | ( wire409 ) | ( wire476 ) | ( wire20988 ) ;
 assign wire20994 = ( n_n2982 ) | ( wire20989 ) | ( _3384 ) ;
 assign wire20998 = ( n_n48  &  n_n15 ) | ( n_n53  &  n_n148 ) ;
 assign wire21010 = ( wire457 ) | ( n_n228  &  wire902  &  n_n53 ) ;
 assign wire21017 = ( n_n5  &  n_n41 ) | ( n_n5  &  wire102 ) | ( n_n5  &  n_n113 ) ;
 assign wire21021 = ( n_n6  &  n_n54 ) | ( n_n48  &  n_n148 ) ;
 assign wire21022 = ( n_n220  &  wire914  &  n_n48 ) | ( wire914  &  n_n256  &  n_n48 ) ;
 assign wire21023 = ( n_n5  &  n_n54 ) | ( n_n48  &  n_n147 ) ;
 assign wire21030 = ( n_n5  &  wire67 ) | ( n_n6  &  wire69 ) ;
 assign wire21042 = ( n_n56  &  n_n226 ) | ( n_n57  &  n_n148 ) ;
 assign wire21043 = ( wire3821 ) | ( n_n56  &  wire160 ) ;
 assign wire21049 = ( n_n220  &  wire914  &  n_n48 ) | ( wire914  &  n_n256  &  n_n48 ) ;
 assign wire21051 = ( wire461 ) | ( wire464 ) | ( wire21049 ) ;
 assign wire21057 = ( wire478 ) | ( n_n3587 ) | ( wire20344 ) ;
 assign wire21059 = ( n_n3827 ) | ( n_n1433 ) | ( wire406 ) | ( wire20343 ) ;
 assign wire21061 = ( wire770 ) | ( wire771 ) | ( wire21057 ) | ( wire21059 ) ;
 assign wire21066 = ( wire95  &  n_n57 ) | ( n_n57  &  wire44 ) | ( n_n57  &  n_n11 ) ;
 assign wire21072 = ( n_n56  &  wire88 ) | ( n_n56  &  n_n29 ) | ( n_n56  &  wire49 ) ;
 assign wire21076 = ( n_n57  &  n_n95 ) | ( n_n145  &  n_n94 ) ;
 assign wire21085 = ( n_n94  &  _38050 ) | ( wire914  &  n_n94  &  _37163 ) ;
 assign wire21092 = ( n_n197  &  n_n94 ) | ( n_n100  &  wire83 ) ;
 assign wire21093 = ( wire21092 ) | ( _3472 ) ;
 assign wire21113 = ( n_n54  &  n_n94 ) | ( n_n100  &  wire77 ) ;
 assign wire21114 = ( wire21113 ) | ( _3430 ) ;
 assign wire21120 = ( wire460 ) | ( wire20193 ) | ( _3414 ) | ( _38093 ) ;
 assign wire21125 = ( wire411 ) | ( _3344 ) | ( n_n5  &  n_n197 ) ;
 assign wire21129 = ( n_n3118 ) | ( n_n3117 ) | ( wire21125 ) | ( _38151 ) ;
 assign wire21143 = ( n_n4  &  n_n108 ) | ( n_n3  &  n_n15 ) ;
 assign wire21146 = ( n_n3506 ) | ( n_n3229 ) | ( wire742 ) | ( wire21143 ) ;
 assign wire21151 = ( n_n3727 ) | ( wire3736 ) | ( n_n4  &  n_n9 ) ;
 assign wire21153 = ( n_n3140 ) | ( n_n3138 ) | ( wire21151 ) ;
 assign wire21157 = ( wire54  &  n_n122 ) | ( n_n111  &  n_n122 ) | ( n_n110  &  n_n122 ) ;
 assign wire21159 = ( i_7_  &  i_6_  &  n_n260  &  n_n116 ) | ( (~ i_7_)  &  i_6_  &  n_n260  &  n_n116 ) | ( i_7_  &  (~ i_6_)  &  n_n260  &  n_n116 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n260  &  n_n116 ) ;
 assign wire21160 = ( n_n5682 ) | ( wire21159 ) | ( n_n111  &  n_n121 ) ;
 assign wire21163 = ( n_n4489 ) | ( wire3733 ) | ( wire21157 ) | ( wire21160 ) ;
 assign wire21164 = ( n_n5769 ) | ( wire48  &  n_n132 ) ;
 assign wire21165 = ( wire364 ) | ( wire48  &  n_n124 ) | ( wire48  &  n_n122 ) ;
 assign wire21169 = ( wire535 ) | ( n_n260  &  n_n118  &  n_n155 ) ;
 assign wire21170 = ( wire777 ) | ( n_n5675 ) | ( wire4928 ) | ( wire19999 ) ;
 assign wire21173 = ( wire879 ) | ( n_n2772 ) | ( wire21169 ) | ( wire21170 ) ;
 assign wire21175 = ( wire394 ) | ( n_n139  &  n_n281  &  wire911 ) ;
 assign wire21180 = ( n_n4  &  n_n108 ) | ( n_n48  &  n_n148 ) ;
 assign wire21183 = ( wire640 ) | ( wire455 ) | ( wire485 ) ;
 assign wire21195 = ( n_n4  &  _38302 ) | ( n_n4  &  wire900  &  _35425 ) ;
 assign wire21196 = ( n_n3  &  _38305 ) | ( n_n3  &  wire898  &  _35396 ) ;
 assign wire21197 = ( n_n3  &  n_n252 ) | ( n_n3  &  n_n14 ) | ( n_n3  &  wire83 ) ;
 assign wire21206 = ( n_n216  &  n_n3 ) | ( n_n4  &  n_n197 ) ;
 assign wire21208 = ( wire333 ) | ( n_n2986 ) | ( wire21206 ) ;
 assign wire21225 = ( n_n4  &  n_n31 ) | ( n_n4  &  n_n76 ) | ( n_n4  &  n_n26 ) ;
 assign wire21233 = ( wire476 ) | ( _3211 ) | ( n_n4  &  _38263 ) ;
 assign wire21238 = ( n_n4  &  _38313 ) | ( n_n4  &  wire908  &  _35046 ) ;
 assign wire21248 = ( n_n257  &  n_n53 ) | ( n_n268  &  wire56 ) ;
 assign wire21252 = ( n_n4  &  _38335 ) | ( wire905  &  n_n4  &  _36337 ) ;
 assign wire21253 = ( n_n4  &  n_n145 ) | ( n_n3  &  n_n14 ) ;
 assign wire21260 = ( n_n4  &  _38339 ) | ( n_n4  &  wire899  &  _37091 ) ;
 assign wire21261 = ( n_n4  &  n_n8 ) | ( n_n4  &  n_n61 ) | ( n_n4  &  n_n144 ) ;
 assign wire21263 = ( wire557 ) | ( wire21260 ) | ( wire21261 ) ;
 assign wire21268 = ( n_n268  &  n_n148 ) | ( n_n265  &  n_n62 ) ;
 assign wire21269 = ( n_n106  &  n_n265 ) | ( n_n4  &  n_n54 ) ;
 assign wire21271 = ( wire913  &  n_n281 ) | ( n_n220  &  wire914 ) ;
 assign wire21288 = ( n_n896 ) | ( _38371 ) ;
 assign wire21298 = ( n_n54  &  n_n57 ) | ( n_n177  &  n_n112 ) ;
 assign wire21299 = ( n_n189  &  n_n109 ) | ( n_n177  &  n_n35 ) ;
 assign wire21329 = ( wire95  &  n_n57 ) | ( n_n57  &  n_n11 ) | ( n_n57  &  n_n148 ) ;
 assign wire21337 = ( n_n1584 ) | ( _2992 ) | ( _2993 ) ;
 assign wire21356 = ( wire635 ) | ( wire3550 ) | ( wire3584 ) | ( wire3585 ) ;
 assign wire21372 = ( n_n4  &  _38725 ) | ( n_n4  &  _38726 ) | ( n_n4  &  _38727 ) ;
 assign wire21385 = ( n_n110  &  n_n268 ) | ( n_n265  &  n_n32 ) ;
 assign wire21394 = ( wire476 ) | ( _2719 ) | ( _2720 ) ;
 assign wire21403 = ( n_n1  &  n_n145 ) | ( n_n1  &  wire1030 ) | ( n_n2  &  wire1030 ) ;
 assign wire21404 = ( n_n268  &  wire264 ) | ( n_n2  &  wire1031 ) ;
 assign wire21408 = ( wire21403 ) | ( wire21404 ) | ( n_n12  &  wire135 ) ;
 assign wire21409 = ( wire3499 ) | ( wire3500 ) ;
 assign wire21415 = ( _2716 ) | ( _38673 ) | ( n_n1  &  wire1102 ) ;
 assign wire21426 = ( n_n4  &  n_n12 ) | ( n_n3  &  n_n66 ) ;
 assign wire21427 = ( n_n4  &  _38740 ) | ( n_n4  &  wire899  &  _34575 ) ;
 assign wire21428 = ( n_n4  &  n_n145 ) | ( n_n4  &  n_n76 ) | ( n_n4  &  n_n26 ) ;
 assign wire21434 = ( n_n281  &  wire902  &  n_n53 ) | ( n_n281  &  wire899  &  n_n53 ) ;
 assign wire21435 = ( n_n2  &  wire78 ) | ( n_n281  &  wire907  &  n_n2 ) ;
 assign wire21438 = ( n_n2274 ) | ( wire3469 ) | ( wire21434 ) ;
 assign wire21448 = ( n_n57  &  n_n95 ) | ( n_n56  &  n_n42 ) ;
 assign wire21455 = ( n_n12  &  n_n100 ) | ( n_n100  &  n_n66 ) | ( n_n12  &  n_n94 ) ;
 assign wire21459 = ( n_n281  &  wire907  &  n_n100 ) | ( n_n281  &  wire908  &  n_n100 ) ;
 assign wire21466 = ( n_n111  &  n_n56 ) | ( n_n57  &  n_n32 ) | ( n_n56  &  n_n32 ) ;
 assign wire21467 = ( n_n57  &  n_n81 ) | ( n_n57  &  wire86 ) | ( n_n57  &  wire1383 ) ;
 assign wire21474 = ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire897 ) | ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  wire897 ) ;
 assign wire21478 = ( n_n94  &  _38614 ) | ( wire903  &  n_n94  &  _35626 ) ;
 assign wire21479 = ( wire21478 ) | ( n_n100  &  wire1413 ) ;
 assign wire21486 = ( n_n57  &  n_n76 ) | ( n_n57  &  n_n26 ) | ( n_n57  &  wire80 ) ;
 assign wire21487 = ( n_n110  &  n_n57 ) | ( n_n57  &  wire19738 ) | ( n_n57  &  n_n67 ) ;
 assign wire21488 = ( n_n110  &  n_n56 ) | ( n_n57  &  n_n108 ) ;
 assign wire21490 = ( n_n56  &  n_n108 ) | ( n_n57  &  n_n148 ) ;
 assign wire21491 = ( n_n106  &  n_n57 ) | ( n_n106  &  n_n56 ) | ( n_n57  &  wire1096 ) ;
 assign wire21493 = ( n_n4916 ) | ( wire3409 ) | ( wire21488 ) | ( wire21491 ) ;
 assign wire21494 = ( wire3402 ) | ( wire3413 ) | ( wire21487 ) | ( wire21490 ) ;
 assign wire21497 = ( n_n186  &  n_n53 ) | ( n_n7  &  wire191 ) ;
 assign wire21499 = ( wire3393 ) | ( wire3400 ) | ( wire3401 ) | ( wire21497 ) ;
 assign wire21500 = ( n_n56  &  n_n76 ) | ( n_n57  &  n_n22 ) ;
 assign wire21501 = ( n_n56  &  wire369 ) | ( n_n220  &  n_n56  &  wire903 ) ;
 assign wire21505 = ( n_n4920 ) | ( n_n4924 ) | ( wire693 ) | ( wire21500 ) ;
 assign wire21506 = ( wire3382 ) | ( wire3416 ) | ( wire21486 ) | ( wire21501 ) ;
 assign wire21521 = ( n_n281  &  wire914  &  n_n4 ) | ( n_n281  &  n_n4  &  wire908 ) ;
 assign wire21522 = ( n_n281  &  wire905  &  n_n4 ) | ( n_n281  &  n_n4  &  wire903 ) ;
 assign wire21525 = ( wire21521 ) | ( wire21522 ) | ( _38713 ) ;
 assign wire21530 = ( n_n281  &  n_n6  &  wire905 ) | ( n_n281  &  n_n6  &  wire908 ) ;
 assign wire21531 = ( n_n60  &  n_n5 ) | ( n_n6  &  wire985 ) | ( n_n5  &  wire985 ) ;
 assign wire21544 = ( n_n110  &  n_n94 ) | ( n_n4  &  n_n30 ) ;
 assign wire21545 = ( wire907  &  n_n279  &  n_n100 ) | ( n_n279  &  wire901  &  n_n100 ) ;
 assign wire21546 = ( n_n106  &  n_n100 ) | ( n_n100  &  n_n33 ) | ( n_n100  &  n_n81 ) ;
 assign wire21569 = ( n_n145  &  n_n48 ) | ( n_n53  &  n_n280 ) ;
 assign wire21614 = ( n_n151  &  n_n4 ) | ( n_n151  &  n_n3 ) | ( n_n3  &  n_n145 ) ;
 assign wire21626 = ( i_7_  &  i_6_  &  n_n284  &  n_n118 ) | ( (~ i_7_)  &  i_6_  &  n_n284  &  n_n118 ) | ( i_7_  &  (~ i_6_)  &  n_n284  &  n_n118 ) ;
 assign wire21627 = ( i_7_  &  i_6_  &  n_n116  &  n_n284 ) | ( (~ i_7_)  &  i_6_  &  n_n116  &  n_n284 ) | ( i_7_  &  (~ i_6_)  &  n_n116  &  n_n284 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n116  &  n_n284 ) ;
 assign wire21628 = ( n_n5769 ) | ( n_n5660 ) | ( n_n151  &  n_n126 ) ;
 assign wire21633 = ( n_n4  &  n_n29 ) | ( n_n4  &  n_n80 ) | ( n_n4  &  wire61 ) ;
 assign wire21647 = ( n_n78 ) | ( wire236 ) | ( wire424 ) | ( wire230 ) ;
 assign wire21651 = ( n_n1  &  n_n64 ) | ( n_n2  &  n_n64 ) | ( n_n1  &  wire1451 ) ;
 assign wire21655 = ( n_n2  &  wire1772 ) | ( n_n1  &  wire1771 ) | ( n_n2  &  wire1771 ) ;
 assign wire21662 = ( n_n110  &  n_n268 ) | ( n_n265  &  n_n62 ) ;
 assign wire21663 = ( n_n3  &  n_n47 ) | ( n_n268  &  n_n147 ) ;
 assign wire21670 = ( wire690 ) | ( wire3178 ) | ( n_n4  &  n_n47 ) ;
 assign wire21671 = ( wire3179 ) | ( wire3213 ) | ( wire3214 ) ;
 assign wire21681 = ( n_n4  &  _39053 ) | ( n_n4  &  wire902  &  _35049 ) ;
 assign wire21694 = ( n_n227  &  n_n28 ) | ( n_n94  &  n_n199 ) ;
 assign wire21695 = ( n_n227  &  wire143 ) | ( n_n207  &  wire1794 ) ;
 assign wire21709 = ( n_n1752 ) | ( _2235 ) | ( _2236 ) | ( _39091 ) ;
 assign wire21715 = ( i_15_  &  n_n242  &  n_n222 ) | ( (~ i_15_)  &  n_n242  &  n_n222 ) | ( i_15_  &  n_n222  &  n_n270 ) | ( (~ i_15_)  &  n_n222  &  n_n270 ) ;
 assign wire21716 = ( n_n220  &  wire905  &  n_n57 ) | ( n_n220  &  n_n57  &  wire903 ) ;
 assign wire21721 = ( n_n56  &  n_n108 ) | ( n_n57  &  wire1198 ) ;
 assign wire21726 = ( n_n57  &  wire1249 ) | ( n_n57  &  wire1248 ) | ( n_n56  &  wire1248 ) ;
 assign wire21732 = ( n_n220  &  wire914  &  n_n57 ) | ( n_n220  &  wire907  &  n_n57 ) ;
 assign wire21733 = ( n_n56  &  n_n32 ) | ( n_n57  &  wire158 ) ;
 assign wire21735 = ( wire200  &  n_n57 ) | ( wire273  &  n_n56 ) ;
 assign wire21737 = ( wire21732 ) | ( wire21735 ) | ( wire200  &  n_n56 ) ;
 assign wire21741 = ( n_n56  &  n_n95 ) | ( n_n57  &  wire429 ) ;
 assign wire21742 = ( wire273  &  n_n57 ) | ( n_n56  &  wire99 ) ;
 assign wire21743 = ( n_n57  &  n_n99 ) | ( n_n8  &  n_n94 ) ;
 assign wire21744 = ( n_n57  &  n_n52 ) | ( wire168  &  wire1195 ) ;
 assign wire21751 = ( n_n147  &  n_n94 ) | ( n_n100  &  n_n64 ) | ( n_n94  &  n_n64 ) ;
 assign wire21752 = ( wire3072 ) | ( wire21743 ) | ( wire21744 ) | ( wire21751 ) ;
 assign wire21753 = ( n_n100  &  wire1597 ) | ( n_n94  &  wire1596 ) ;
 assign wire21756 = ( n_n281  &  wire911  &  n_n94 ) | ( wire911  &  n_n256  &  n_n94 ) ;
 assign wire21757 = ( n_n110  &  n_n94 ) | ( n_n94  &  n_n203 ) | ( n_n94  &  n_n68 ) ;
 assign wire21759 = ( wire3056 ) | ( wire21756 ) | ( wire21757 ) ;
 assign wire21760 = ( wire3065 ) | ( n_n100  &  wire1599 ) | ( n_n100  &  wire1730 ) ;
 assign wire21761 = ( n_n57  &  n_n95 ) | ( n_n56  &  n_n42 ) ;
 assign wire21762 = ( n_n57  &  wire494 ) | ( n_n220  &  n_n57  &  wire906 ) ;
 assign wire21764 = ( n_n57  &  wire99 ) | ( n_n57  &  wire180 ) ;
 assign wire21780 = ( n_n53  &  _39283 ) | ( wire907  &  n_n53  &  _36212 ) ;
 assign wire21781 = ( n_n48  &  _39286 ) | ( n_n48  &  n_n247  &  _36683 ) ;
 assign wire21790 = ( n_n6  &  n_n95 ) | ( n_n5  &  n_n47 ) ;
 assign wire21811 = ( n_n6  &  wire1290 ) | ( n_n6  &  wire1289 ) | ( n_n5  &  wire1289 ) ;
 assign wire21815 = ( wire164  &  n_n150 ) | ( n_n207  &  wire425 ) ;
 assign wire21844 = ( n_n53  &  _39113 ) | ( wire899  &  n_n53  &  _37042 ) ;
 assign wire21845 = ( n_n53  &  n_n107 ) | ( n_n53  &  n_n20 ) | ( n_n53  &  wire1803 ) ;
 assign wire21849 = ( n_n111  &  n_n48 ) | ( n_n53  &  n_n80 ) ;
 assign wire21850 = ( n_n281  &  wire912  &  n_n48 ) | ( wire912  &  n_n256  &  n_n48 ) ;
 assign wire21853 = ( wire2942 ) | ( wire2943 ) | ( wire21849 ) | ( wire21850 ) ;
 assign wire21859 = ( i_7_  &  i_6_  &  n_n260  &  n_n118 ) | ( (~ i_7_)  &  i_6_  &  n_n260  &  n_n118 ) | ( i_7_  &  (~ i_6_)  &  n_n260  &  n_n118 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n260  &  n_n118 ) ;
 assign wire21860 = ( i_7_  &  i_6_  &  n_n260  &  n_n116 ) | ( (~ i_7_)  &  i_6_  &  n_n260  &  n_n116 ) | ( i_7_  &  (~ i_6_)  &  n_n260  &  n_n116 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n260  &  n_n116 ) ;
 assign wire21861 = ( wire21859 ) | ( n_n142  &  wire1593 ) ;
 assign wire21862 = ( wire503 ) | ( wire21860 ) | ( wire48  &  n_n152 ) ;
 assign wire21872 = ( wire912  &  n_n225  &  n_n94 ) | ( wire912  &  n_n256  &  n_n94 ) ;
 assign wire21884 = ( n_n4  &  n_n108 ) | ( n_n4  &  n_n107 ) | ( n_n4  &  n_n221 ) ;
 assign wire21902 = ( wire3228 ) | ( wire21633 ) | ( _39382 ) ;
 assign wire21910 = ( wire333 ) | ( wire485 ) | ( _39450 ) ;
 assign wire21912 = ( n_n4  &  n_n252 ) | ( n_n3  &  wire83 ) ;
 assign wire21918 = ( n_n4  &  _39425 ) | ( wire905  &  n_n4  &  _36337 ) ;
 assign wire21920 = ( wire2874 ) | ( wire21918 ) | ( n_n3  &  wire1112 ) ;
 assign wire21922 = ( n_n3  &  _39432 ) | ( n_n3  &  wire904  &  _35391 ) ;
 assign wire21923 = ( n_n4  &  n_n64 ) | ( n_n3  &  n_n64 ) | ( n_n4  &  n_n13 ) | ( n_n3  &  n_n13 ) ;
 assign wire21925 = ( wire2864 ) | ( wire21922 ) | ( wire21923 ) ;
 assign wire21926 = ( n_n1320 ) | ( wire2883 ) | ( wire2885 ) | ( wire21912 ) ;
 assign wire21927 = ( n_n1157 ) | ( wire21920 ) | ( wire21925 ) ;
 assign wire21928 = ( wire2888 ) | ( wire2889 ) | ( wire21910 ) | ( wire21926 ) ;
 assign wire21933 = ( n_n4  &  n_n31 ) | ( n_n4  &  n_n26 ) | ( n_n4  &  n_n80 ) ;
 assign wire21948 = ( wire519 ) | ( wire2845 ) | ( _39495 ) ;
 assign wire21950 = ( n_n1108 ) | ( wire21941 ) | ( wire21948 ) | ( _39486 ) ;
 assign wire21956 = ( n_n1412 ) | ( _1195 ) | ( _1196 ) ;
 assign wire21962 = ( _1194 ) | ( n_n1  &  wire245 ) | ( n_n1  &  n_n39 ) ;
 assign wire21968 = ( n_n3768 ) | ( n_n3770 ) | ( n_n2  &  wire1424 ) ;
 assign wire21969 = ( wire21968 ) | ( _1215 ) | ( _1216 ) ;
 assign wire21970 = ( wire2839 ) | ( wire2842 ) | ( wire21956 ) | ( wire21962 ) ;
 assign wire21973 = ( n_n2  &  n_n257 ) | ( n_n268  &  wire56 ) ;
 assign wire21977 = ( n_n253  &  _39961 ) | ( n_n253  &  _39962 ) ;
 assign wire21981 = ( n_n3523 ) | ( n_n2  &  wire1514 ) ;
 assign wire21982 = ( i_14_  &  i_13_  &  i_12_  &  wire905 ) | ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire905 ) | ( i_14_  &  i_13_  &  (~ i_12_)  &  wire905 ) | ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  wire905 ) | ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire905 ) ;
 assign wire21987 = ( n_n3255 ) | ( n_n1  &  wire100 ) | ( n_n1  &  wire21982 ) ;
 assign wire21988 = ( n_n1  &  n_n10 ) | ( n_n2  &  n_n10 ) | ( n_n2  &  n_n62 ) ;
 assign wire21991 = ( wire2813 ) | ( wire2814 ) | ( wire2830 ) | ( wire2831 ) ;
 assign wire21992 = ( wire2827 ) | ( wire21973 ) | ( wire21988 ) | ( wire21991 ) ;
 assign wire21993 = ( wire2822 ) | ( wire2825 ) | ( wire21981 ) | ( wire21987 ) ;
 assign wire22002 = ( n_n220  &  wire914 ) | ( wire914  &  n_n256 ) | ( n_n220  &  wire897 ) ;
 assign wire22005 = ( n_n268  &  n_n240 ) | ( n_n265  &  n_n10 ) ;
 assign wire22010 = ( n_n4  &  n_n105 ) | ( n_n4  &  n_n47 ) | ( n_n4  &  n_n46 ) ;
 assign wire22012 = ( n_n1359 ) | ( n_n1363 ) | ( wire22010 ) ;
 assign wire22035 = ( n_n220  &  wire899  &  n_n53 ) | ( n_n281  &  wire899  &  n_n53 ) ;
 assign wire22039 = ( n_n1  &  wire41 ) | ( n_n2  &  wire1171 ) ;
 assign wire22047 = ( n_n4  &  _39839 ) | ( n_n4  &  wire900  &  _35425 ) ;
 assign wire22048 = ( n_n258  &  wire899  &  n_n53 ) | ( n_n222  &  wire899  &  n_n53 ) ;
 assign wire22050 = ( n_n53  &  n_n31 ) | ( n_n53  &  wire42 ) | ( n_n53  &  n_n80 ) ;
 assign wire22052 = ( n_n53  &  wire61 ) | ( n_n53  &  wire140 ) | ( n_n53  &  n_n27 ) ;
 assign wire22070 = ( n_n147  &  n_n94 ) | ( n_n100  &  n_n81 ) ;
 assign wire22071 = ( n_n104  &  n_n100 ) | ( n_n110  &  n_n94 ) ;
 assign wire22081 = ( n_n227  &  n_n28 ) | ( n_n94  &  n_n203 ) ;
 assign wire22082 = ( n_n279  &  wire903  &  n_n94 ) | ( n_n222  &  wire903  &  n_n94 ) ;
 assign wire22083 = ( n_n257  &  n_n227 ) | ( n_n207  &  wire232 ) ;
 assign wire22084 = ( wire40  &  n_n94 ) | ( n_n74  &  n_n94 ) | ( n_n94  &  n_n24 ) ;
 assign wire22090 = ( n_n4  &  _39878 ) | ( n_n4  &  wire906  &  _35716 ) ;
 assign wire22093 = ( n_n1359 ) | ( wire333 ) | ( wire455 ) | ( wire22090 ) ;
 assign wire22097 = ( wire2708 ) | ( wire2709 ) ;
 assign wire22101 = ( n_n1217 ) | ( wire22097 ) | ( _39906 ) | ( _39908 ) ;
 assign wire22117 = ( n_n4846 ) | ( n_n4852 ) | ( n_n1490 ) ;
 assign wire22124 = ( n_n6  &  n_n54 ) | ( n_n53  &  n_n10 ) ;
 assign wire22125 = ( n_n220  &  wire914  &  n_n48 ) | ( wire914  &  n_n256  &  n_n48 ) ;
 assign wire22126 = ( n_n246  &  n_n48 ) | ( n_n48  &  n_n135 ) | ( n_n48  &  n_n86 ) ;
 assign wire22140 = ( n_n37  &  n_n53 ) | ( n_n48  &  wire223 ) ;
 assign wire22154 = ( n_n53  &  n_n197 ) | ( n_n53  &  n_n107 ) | ( n_n53  &  n_n221 ) ;
 assign wire22160 = ( n_n48  &  wire82 ) | ( n_n228  &  wire905  &  n_n48 ) ;
 assign wire22164 = ( n_n220  &  wire905 ) | ( wire907  &  n_n258 ) ;
 assign wire22174 = ( n_n3827 ) | ( n_n53  &  wire124 ) | ( n_n53  &  wire212 ) ;
 assign wire22181 = ( n_n110  &  n_n94 ) | ( n_n133  &  n_n94 ) | ( n_n94  &  n_n203 ) ;
 assign wire22208 = ( n_n267  &  _39758 ) | ( n_n267  &  _39759 ) ;
 assign wire22217 = ( n_n57  &  n_n50 ) | ( n_n94  &  n_n150 ) ;
 assign wire22255 = ( n_n253  &  _39529 ) | ( n_n253  &  _39530 ) ;
 assign wire22262 = ( wire407 ) | ( wire457 ) | ( wire75  &  n_n57 ) ;
 assign wire22273 = ( n_n267  &  _39555 ) | ( n_n267  &  _39556 ) ;
 assign wire22282 = ( n_n281  &  wire902  &  n_n53 ) | ( wire902  &  n_n258  &  n_n53 ) ;
 assign wire22302 = ( wire2495 ) | ( _39578 ) | ( _39580 ) ;
 assign wire22308 = ( n_n1597 ) | ( n_n1598 ) | ( wire704 ) ;
 assign wire22312 = ( n_n111  &  n_n56 ) | ( n_n57  &  wire49 ) ;
 assign wire22314 = ( wire762 ) | ( n_n1591 ) | ( wire22312 ) ;
 assign wire22317 = ( n_n56  &  wire49 ) | ( n_n57  &  n_n22 ) ;
 assign wire22322 = ( wire2486 ) | ( wire2491 ) | ( wire22308 ) | ( wire22314 ) ;
 assign wire22326 = ( wire2521 ) | ( wire22277 ) | ( _39571 ) | ( _39582 ) ;
 assign wire22327 = ( n_n1095 ) | ( _39645 ) | ( _39646 ) | ( _39664 ) ;
 assign wire22328 = ( n_n1097 ) | ( n_n1102 ) | ( n_n1101 ) | ( n_n1103 ) ;
 assign wire22330 = ( wire21969 ) | ( wire21970 ) | ( wire21992 ) | ( wire21993 ) ;
 assign wire22332 = ( n_n1092 ) | ( n_n1093 ) | ( wire22101 ) | ( wire22330 ) ;
 assign wire22337 = ( n_n4  &  n_n70 ) | ( n_n4  &  n_n197 ) | ( n_n4  &  n_n21 ) ;
 assign wire22346 = ( n_n4  &  _40413 ) | ( n_n4  &  wire906  &  _35716 ) ;
 assign wire22356 = ( wire642 ) | ( n_n3  &  wire1217 ) ;
 assign wire22366 = ( wire907  &  n_n258 ) | ( n_n258  &  wire904 ) ;
 assign wire22369 = ( wire907  &  n_n258  &  n_n100 ) | ( wire911  &  n_n258  &  n_n100 ) ;
 assign wire22370 = ( n_n100  &  n_n13 ) | ( n_n94  &  n_n13 ) | ( n_n100  &  wire1066 ) ;
 assign wire22378 = ( n_n54  &  n_n57 ) | ( n_n61  &  n_n94 ) ;
 assign wire22379 = ( n_n257  &  n_n100 ) | ( n_n257  &  n_n94 ) | ( n_n100  &  n_n236 ) ;
 assign wire22380 = ( n_n240  &  wire168 ) | ( n_n57  &  wire486 ) ;
 assign wire22389 = ( n_n197  &  n_n100 ) | ( n_n216  &  n_n94 ) ;
 assign wire22395 = ( wire911  &  n_n258  &  n_n48 ) | ( wire911  &  n_n258  &  n_n53 ) ;
 assign wire22399 = ( n_n48  &  n_n197 ) | ( n_n53  &  n_n197 ) | ( n_n53  &  wire123 ) ;
 assign wire22443 = ( n_n48  &  n_n31 ) | ( n_n53  &  n_n26 ) ;
 assign wire22449 = ( wire112  &  n_n53 ) | ( n_n258  &  wire901  &  n_n53 ) ;
 assign wire22456 = ( n_n56  &  wire1677 ) | ( n_n57  &  wire1676 ) | ( n_n56  &  wire1676 ) ;
 assign wire22461 = ( n_n48  &  n_n104 ) | ( n_n53  &  n_n41 ) ;
 assign wire22489 = ( i_7_  &  i_6_  &  n_n118  &  n_n230 ) | ( (~ i_7_)  &  i_6_  &  n_n118  &  n_n230 ) | ( i_7_  &  (~ i_6_)  &  n_n118  &  n_n230 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n118  &  n_n230 ) ;
 assign wire22490 = ( i_7_  &  i_6_  &  n_n116  &  n_n230 ) | ( (~ i_7_)  &  i_6_  &  n_n116  &  n_n230 ) | ( i_7_  &  (~ i_6_)  &  n_n116  &  n_n230 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n116  &  n_n230 ) ;
 assign wire22491 = ( wire22489 ) | ( n_n136  &  wire1307 ) ;
 assign wire22492 = ( wire394 ) | ( wire22490 ) | ( n_n139  &  wire48 ) ;
 assign wire22502 = ( wire688 ) | ( wire2269 ) | ( _40385 ) ;
 assign wire22511 = ( wire2264 ) | ( wire2267 ) | ( wire2268 ) ;
 assign wire22518 = ( wire2263 ) | ( n_n2  &  wire1311 ) | ( n_n2  &  wire1733 ) ;
 assign wire22523 = ( i_15_  &  n_n258  &  n_n267 ) | ( i_15_  &  n_n256  &  n_n267 ) | ( (~ i_15_)  &  n_n256  &  n_n267 ) ;
 assign wire22532 = ( n_n268  &  n_n240 ) | ( n_n3  &  wire408 ) ;
 assign wire22538 = ( n_n1  &  n_n236 ) | ( n_n1  &  wire1673 ) | ( n_n2  &  wire1673 ) ;
 assign wire22539 = ( n_n1  &  n_n240 ) | ( n_n2  &  n_n240 ) | ( n_n2  &  wire403 ) ;
 assign wire22541 = ( n_n1  &  wire1357 ) | ( n_n1  &  wire1355 ) | ( n_n2  &  wire1355 ) ;
 assign wire22543 = ( wire2225 ) | ( wire22538 ) | ( wire22539 ) | ( wire22541 ) ;
 assign wire22551 = ( n_n246  &  n_n94 ) | ( n_n257  &  n_n207 ) ;
 assign wire22552 = ( n_n4  &  n_n26 ) | ( n_n104  &  n_n100 ) ;
 assign wire22566 = ( n_n6  &  n_n240 ) | ( n_n103  &  n_n207 ) ;
 assign wire22567 = ( n_n5  &  n_n257 ) | ( n_n227  &  wire276 ) ;
 assign wire22570 = ( n_n6  &  wire1680 ) | ( n_n6  &  wire1679 ) | ( n_n5  &  wire1679 ) ;
 assign wire22571 = ( n_n207  &  wire292 ) | ( n_n5  &  wire1682 ) ;
 assign wire22574 = ( n_n4  &  n_n258  &  wire906 ) | ( n_n4  &  n_n258  &  wire900 ) ;
 assign wire22575 = ( n_n4  &  _40232 ) | ( n_n4  &  wire908  &  _35046 ) ;
 assign wire22576 = ( n_n4  &  n_n70 ) | ( n_n3  &  n_n49 ) ;
 assign wire22578 = ( wire22574 ) | ( wire22575 ) | ( wire22576 ) ;
 assign wire22590 = ( n_n3  &  n_n61 ) | ( n_n4  &  n_n257 ) | ( n_n3  &  n_n257 ) ;
 assign wire22593 = ( n_n380 ) | ( n_n381 ) | ( wire2176 ) | ( wire22590 ) ;
 assign wire22596 = ( n_n4  &  wire88 ) | ( n_n4  &  n_n80 ) | ( n_n4  &  wire114 ) ;
 assign wire22600 = ( n_n216  &  n_n3 ) | ( n_n4  &  n_n197 ) ;
 assign wire22606 = ( wire911  &  n_n258  &  n_n94 ) | ( n_n258  &  wire899  &  n_n94 ) ;
 assign wire22618 = ( n_n100  &  wire1121 ) | ( n_n94  &  wire1120 ) ;
 assign wire22633 = ( wire571 ) | ( wire737 ) | ( n_n105  &  n_n48 ) ;
 assign wire22635 = ( wire5591 ) | ( wire5592 ) | ( n_n9  &  n_n56 ) ;
 assign wire22636 = ( n_n57  &  n_n226 ) | ( n_n56  &  n_n226 ) | ( n_n57  &  wire1717 ) | ( n_n56  &  wire1717 ) ;
 assign wire22637 = ( n_n57  &  n_n65 ) | ( n_n56  &  n_n65 ) | ( n_n57  &  n_n11 ) ;
 assign wire22638 = ( n_n57  &  wire1753 ) | ( n_n56  &  wire1752 ) ;
 assign wire22639 = ( wire22635 ) | ( wire22636 ) | ( wire22637 ) ;
 assign wire22640 = ( wire2122 ) | ( wire22633 ) | ( wire22638 ) ;
 assign wire22642 = ( n_n56  &  n_n179 ) | ( n_n56  &  wire55 ) | ( n_n56  &  wire190 ) ;
 assign wire22643 = ( n_n57  &  wire190 ) | ( n_n57  &  wire198 ) ;
 assign wire22651 = ( n_n100  &  n_n103 ) | ( n_n94  &  n_n39 ) ;
 assign wire22652 = ( n_n31  &  n_n100 ) | ( n_n94  &  n_n103 ) ;
 assign wire22658 = ( n_n94  &  n_n41 ) | ( n_n100  &  n_n36 ) ;
 assign wire22659 = ( n_n37  &  n_n100 ) | ( n_n104  &  n_n100 ) | ( n_n100  &  n_n84 ) ;
 assign wire22665 = ( n_n105  &  n_n100 ) | ( n_n54  &  n_n94 ) ;
 assign wire22667 = ( n_n3884 ) | ( wire22665 ) | ( n_n94  &  wire139 ) ;
 assign wire22668 = ( wire776 ) | ( wire2072 ) ;
 assign wire22672 = ( n_n6  &  wire120 ) | ( n_n6  &  wire19457 ) | ( n_n6  &  n_n25 ) ;
 assign wire22680 = ( n_n6  &  n_n228  &  wire899 ) | ( n_n6  &  n_n228  &  wire897 ) ;
 assign wire22681 = ( n_n6  &  n_n206 ) | ( n_n206  &  n_n5 ) | ( n_n5  &  wire1253 ) ;
 assign wire22683 = ( n_n6  &  wire1640 ) | ( n_n6  &  wire1638 ) | ( n_n5  &  wire1638 ) ;
 assign wire22684 = ( n_n227  &  wire275 ) | ( n_n5  &  wire1639 ) ;
 assign wire22689 = ( n_n6  &  wire114 ) | ( n_n6  &  n_n258  &  wire897 ) ;
 assign wire22692 = ( wire22672 ) | ( n_n5  &  wire1641 ) | ( n_n5  &  wire1918 ) ;
 assign wire22695 = ( wire88  &  n_n48 ) | ( n_n48  &  n_n31 ) | ( n_n48  &  n_n80 ) ;
 assign wire22698 = ( n_n216  &  n_n48 ) | ( n_n216  &  n_n53 ) | ( n_n53  &  n_n197 ) ;
 assign wire22700 = ( wire2034 ) | ( wire2035 ) ;
 assign wire22701 = ( n_n4073 ) | ( wire2041 ) | ( wire22695 ) | ( wire22698 ) ;
 assign wire22703 = ( n_n48  &  n_n103 ) | ( n_n53  &  n_n103 ) | ( n_n53  &  wire114 ) ;
 assign wire22704 = ( n_n53  &  n_n104 ) | ( n_n48  &  n_n41 ) ;
 assign wire22708 = ( n_n4094 ) | ( n_n4090 ) | ( wire2023 ) | ( wire22704 ) ;
 assign wire22709 = ( wire483 ) | ( wire2022 ) | ( wire2030 ) | ( wire22703 ) ;
 assign wire22712 = ( wire912  &  n_n258  &  n_n53 ) | ( n_n258  &  wire900  &  n_n53 ) ;
 assign wire22720 = ( n_n6  &  n_n54 ) | ( n_n53  &  n_n63 ) ;
 assign wire22732 = ( n_n48  &  n_n197 ) | ( n_n48  &  wire1063 ) | ( n_n53  &  wire1063 ) ;
 assign wire22742 = ( n_n4644 ) | ( wire1977 ) | ( n_n5  &  n_n54 ) ;
 assign wire22780 = ( n_n1  &  n_n59 ) | ( n_n2  &  n_n59 ) | ( n_n1  &  wire1606 ) ;
 assign wire22786 = ( n_n4  &  _40548 ) | ( n_n4  &  wire902  &  _35056 ) ;
 assign wire22787 = ( n_n228  &  n_n4  &  wire899 ) | ( n_n228  &  n_n4  &  wire900 ) ;
 assign wire22788 = ( n_n4  &  n_n197 ) | ( n_n3  &  n_n15 ) ;
 assign wire22801 = ( n_n204  &  n_n94 ) | ( n_n100  &  n_n84 ) ;
 assign wire22805 = ( n_n4  &  n_n31 ) | ( n_n94  &  n_n39 ) ;
 assign wire22806 = ( n_n11  &  n_n94 ) | ( n_n100  &  n_n63 ) ;
 assign wire22820 = ( n_n785 ) | ( wire529 ) | ( _40671 ) | ( _40672 ) ;
 assign wire22837 = ( n_n4  &  n_n65 ) | ( n_n3  &  n_n15 ) ;
 assign wire22843 = ( wire238 ) | ( n_n4  &  wire126 ) | ( n_n4  &  n_n31 ) ;
 assign wire22844 = ( wire2170 ) | ( wire2173 ) | ( wire2174 ) | ( wire22596 ) ;
 assign _61 = ( n_n208  &  n_n284  &  n_n285  &  wire1837 ) ;
 assign _92 = ( n_n3  &  wire88 ) | ( n_n3  &  wire20149 ) | ( n_n3  &  _40812 ) ;
 assign _140 = ( n_n5  &  wire469 ) | ( n_n5  &  wire128 ) | ( n_n5  &  _143 ) ;
 assign _143 = ( i_14_  &  i_13_  &  (~ i_12_)  &  wire899 ) ;
 assign _231 = ( n_n57  &  wire60 ) | ( n_n57  &  wire227 ) | ( n_n57  &  _237 ) ;
 assign _235 = ( n_n56  &  wire60 ) | ( n_n56  &  wire227 ) | ( n_n56  &  _237 ) ;
 assign _237 = ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire911 ) ;
 assign _290 = ( n_n94  &  wire469 ) | ( n_n94  &  wire128 ) | ( n_n94  &  _40678 ) ;
 assign _339 = ( n_n265  &  wire901  &  _36817 ) ;
 assign _350 = ( n_n284  &  n_n285  &  n_n266  &  wire85 ) ;
 assign _358 = ( n_n2  &  wire60 ) | ( n_n2  &  wire198 ) | ( n_n2  &  _361 ) ;
 assign _361 = ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire911 ) ;
 assign _367 = ( n_n2  &  wire254 ) | ( n_n2  &  wire301 ) | ( n_n2  &  wire335 ) ;
 assign _370 = ( n_n1  &  wire55 ) | ( n_n1  &  wire304 ) | ( n_n1  &  _373 ) ;
 assign _373 = ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire912 ) ;
 assign _379 = ( n_n1  &  wire301 ) | ( n_n1  &  wire277 ) | ( n_n1  &  wire275 ) ;
 assign _380 = ( n_n1  &  wire190 ) | ( n_n1  &  wire198 ) ;
 assign _382 = ( n_n2  &  wire55 ) | ( n_n2  &  wire190 ) | ( n_n2  &  _385 ) ;
 assign _385 = ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire912 ) ;
 assign _399 = ( n_n2  &  wire126 ) | ( n_n2  &  wire89 ) | ( n_n2  &  _40584 ) ;
 assign _455 = ( n_n5  &  wire89 ) | ( n_n5  &  wire96 ) | ( n_n5  &  _40536 ) ;
 assign _492 = ( wire912  &  n_n48  &  _36184 ) ;
 assign _506 = ( n_n264  &  n_n273  &  n_n285  &  wire301 ) ;
 assign _560 = ( n_n48  &  wire96 ) | ( n_n48  &  wire134 ) | ( n_n48  &  _562 ) ;
 assign _561 = ( n_n48  &  wire19577 ) | ( n_n48  &  wire139 ) | ( n_n48  &  _567 ) ;
 assign _562 = ( i_14_  &  i_13_  &  (~ i_12_)  &  wire898 ) ;
 assign _567 = ( i_14_  &  i_13_  &  i_12_  &  wire906 ) ;
 assign _605 = ( n_n4  &  wire65 ) | ( n_n4  &  wire47 ) | ( n_n4  &  _40420 ) ;
 assign _608 = ( n_n3  &  wire320 ) | ( n_n3  &  wire22335 ) | ( n_n3  &  _40418 ) ;
 assign _614 = ( n_n4  &  wire245 ) | ( n_n4  &  wire22341 ) | ( n_n4  &  _40408 ) ;
 assign _617 = ( n_n3  &  wire22341 ) | ( n_n3  &  wire47 ) | ( n_n3  &  _40405 ) ;
 assign _632 = ( n_n4  &  wire514 ) | ( n_n4  &  wire232 ) | ( n_n4  &  _635 ) ;
 assign _635 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire911 ) ;
 assign _654 = ( n_n139  &  wire54 ) | ( n_n139  &  _40371 ) ;
 assign _655 = ( n_n139  &  wire103 ) | ( n_n139  &  n_n220  &  wire914 ) ;
 assign _675 = ( wire41  &  n_n100 ) | ( n_n100  &  n_n41 ) | ( n_n100  &  _40345 ) ;
 assign _696 = ( n_n57  &  wire53 ) | ( n_n57  &  wire405 ) | ( n_n57  &  _699 ) ;
 assign _699 = ( i_14_  &  (~ i_13_)  &  i_12_  &  wire897 ) ;
 assign _702 = ( n_n57  &  wire233 ) | ( n_n57  &  wire444 ) | ( n_n57  &  _710 ) ;
 assign _703 = ( n_n57  &  wire57 ) | ( n_n57  &  wire414 ) | ( n_n57  &  _713 ) ;
 assign _705 = ( n_n56  &  wire233 ) | ( n_n56  &  wire444 ) | ( n_n56  &  _710 ) ;
 assign _706 = ( n_n56  &  wire57 ) | ( n_n56  &  wire414 ) | ( n_n56  &  _713 ) ;
 assign _710 = ( i_14_  &  i_13_  &  (~ i_12_)  &  wire907 ) ;
 assign _713 = ( i_14_  &  (~ i_13_)  &  i_12_  &  wire912 ) ;
 assign _716 = ( wire906  &  wire191  &  _35394 ) ;
 assign _719 = ( n_n56  &  wire42 ) | ( n_n56  &  _40311 ) ;
 assign _720 = ( n_n56  &  wire52 ) | ( n_n56  &  wire441 ) | ( n_n56  &  _728 ) ;
 assign _721 = ( n_n56  &  wire292 ) | ( n_n258  &  n_n56  &  wire904 ) ;
 assign _725 = ( n_n57  &  wire52 ) | ( n_n57  &  wire441 ) | ( n_n57  &  _728 ) ;
 assign _726 = ( n_n57  &  wire292 ) | ( n_n258  &  n_n57  &  wire904 ) ;
 assign _727 = ( wire914  &  n_n57  &  _37163 ) ;
 assign _728 = ( i_14_  &  (~ i_13_)  &  i_12_  &  wire911 ) ;
 assign _774 = ( wire902  &  n_n53  &  _35622 ) ;
 assign _788 = ( n_n5  &  wire65 ) | ( n_n5  &  wire22335 ) | ( n_n5  &  _40272 ) ;
 assign _793 = ( n_n6  &  wire306 ) | ( n_n6  &  wire22335 ) | ( n_n6  &  _796 ) ;
 assign _796 = ( i_14_  &  i_13_  &  (~ i_12_)  &  wire903 ) ;
 assign _801 = ( n_n6  &  wire65 ) | ( n_n6  &  wire276 ) | ( n_n6  &  _40266 ) ;
 assign _808 = ( n_n6  &  wire351 ) | ( n_n6  &  wire233 ) | ( n_n6  &  _40259 ) ;
 assign _817 = ( n_n5  &  wire22340 ) | ( n_n5  &  wire47 ) | ( n_n5  &  _40250 ) ;
 assign _822 = ( n_n5  &  wire143 ) | ( n_n5  &  wire1649 ) | ( n_n5  &  _40246 ) ;
 assign _830 = ( n_n6  &  wire514 ) | ( n_n6  &  wire232 ) | ( n_n6  &  _40239 ) ;
 assign _833 = ( n_n5  &  wire514 ) | ( n_n5  &  wire232 ) | ( n_n5  &  _40239 ) ;
 assign _834 = ( n_n285  &  n_n230  &  n_n263  &  wire306 ) ;
 assign _848 = ( n_n4  &  wire906  &  n_n256 ) ;
 assign _897 = ( n_n6  &  wire408 ) | ( n_n6  &  wire22341 ) | ( n_n6  &  _40195 ) ;
 assign _899 = ( n_n5  &  wire408 ) | ( n_n5  &  wire22341 ) | ( n_n5  &  _40195 ) ;
 assign _900 = ( n_n285  &  n_n230  &  n_n263  &  wire357 ) ;
 assign _945 = ( n_n260  &  n_n285  &  n_n263  &  wire140 ) ;
 assign _946 = ( n_n260  &  n_n285  &  n_n263  &  wire1069 ) ;
 assign _995 = ( n_n94  &  wire52 ) | ( n_n94  &  wire22366 ) | ( n_n94  &  _998 ) ;
 assign _998 = ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire913 ) ;
 assign _1010 = ( n_n268  &  wire53 ) | ( n_n268  &  wire52 ) | ( n_n268  &  _40103 ) ;
 assign _1051 = ( n_n265  &  wire233 ) | ( n_n265  &  wire414 ) | ( n_n265  &  _40078 ) ;
 assign _1054 = ( n_n4  &  wire357 ) | ( n_n4  &  wire22340 ) | ( n_n4  &  _40072 ) ;
 assign _1064 = ( n_n268  &  wire57 ) | ( n_n268  &  wire444 ) | ( n_n268  &  _1067 ) ;
 assign _1067 = ( i_14_  &  (~ i_13_)  &  i_12_  &  wire912 ) ;
 assign _1102 = ( n_n1  &  wire57 ) | ( n_n1  &  wire229 ) | ( n_n1  &  _40037 ) ;
 assign _1166 = ( n_n2  &  wire343 ) | ( n_n2  &  wire431 ) ;
 assign _1167 = ( n_n2  &  wire62 ) | ( n_n2  &  wire65 ) | ( n_n2  &  _39957 ) ;
 assign _1168 = ( n_n2  &  wire84 ) | ( n_n2  &  _39959 ) ;
 assign _1194 = ( n_n1  &  wire67 ) | ( n_n1  &  wire347 ) | ( n_n1  &  _39937 ) ;
 assign _1195 = ( n_n2  &  wire245 ) | ( n_n2  &  wire912  &  n_n225 ) ;
 assign _1196 = ( n_n2  &  wire67 ) | ( n_n2  &  wire347 ) | ( n_n2  &  _39934 ) ;
 assign _1203 = ( n_n2  &  wire85 ) | ( n_n2  &  wire437 ) | ( n_n2  &  _1206 ) ;
 assign _1204 = ( n_n2  &  wire41 ) | ( n_n2  &  wire47 ) | ( n_n2  &  _1209 ) ;
 assign _1205 = ( n_n2  &  wire99 ) | ( n_n2  &  _39929 ) ;
 assign _1206 = ( i_14_  &  i_13_  &  i_12_  &  wire907 ) ;
 assign _1209 = ( (~ i_14_)  &  i_13_  &  i_12_  &  wire901 ) ;
 assign _1215 = ( n_n1  &  wire346 ) | ( n_n1  &  wire431 ) ;
 assign _1216 = ( n_n1  &  wire40 ) | ( n_n1  &  _39925 ) ;
 assign _1248 = ( n_n6  &  wire73 ) | ( n_n6  &  wire52 ) | ( n_n6  &  _39893 ) ;
 assign _1251 = ( n_n5  &  wire83 ) | ( n_n5  &  wire274 ) | ( n_n5  &  _1254 ) ;
 assign _1254 = ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  wire899 ) ;
 assign _1261 = ( n_n5  &  wire60 ) | ( n_n5  &  wire325 ) | ( n_n5  &  _1263 ) ;
 assign _1262 = ( n_n5  &  wire165 ) | ( n_n5  &  wire514 ) | ( n_n5  &  _1266 ) ;
 assign _1263 = ( i_14_  &  i_13_  &  i_12_  &  wire913 ) ;
 assign _1266 = ( (~ i_14_)  &  i_13_  &  i_12_  &  wire911 ) ;
 assign _1292 = ( n_n227  &  wire143 ) | ( n_n227  &  wire306 ) | ( n_n227  &  _39861 ) ;
 assign _1305 = ( n_n2  &  wire19385 ) | ( n_n2  &  n_n256  &  wire900 ) ;
 assign _1306 = ( n_n2  &  wire51 ) | ( n_n2  &  wire448 ) | ( n_n2  &  _39848 ) ;
 assign _1338 = ( n_n94  &  wire77 ) | ( n_n94  &  wire311 ) | ( n_n94  &  _1340 ) ;
 assign _1340 = ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  wire898 ) ;
 assign _1346 = ( wire55  &  n_n100 ) | ( n_n100  &  wire81 ) | ( n_n100  &  _1349 ) ;
 assign _1349 = ( i_14_  &  i_13_  &  i_12_  &  wire914 ) ;
 assign _1354 = ( wire19578  &  n_n94 ) | ( n_n94  &  wire300 ) | ( n_n94  &  _1357 ) ;
 assign _1357 = ( i_14_  &  i_13_  &  (~ i_12_)  &  wire906 ) ;
 assign _1360 = ( n_n100  &  wire807 ) | ( n_n100  &  wire311 ) | ( n_n100  &  _1363 ) ;
 assign _1363 = ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire904 ) ;
 assign _1372 = ( n_n258  &  wire898  &  n_n100 ) ;
 assign _1394 = ( n_n56  &  wire19578 ) | ( n_n56  &  wire81 ) | ( n_n56  &  _39772 ) ;
 assign _1427 = ( n_n100  &  wire56 ) | ( n_n100  &  wire345 ) | ( n_n100  &  _1430 ) ;
 assign _1428 = ( n_n100  &  wire104 ) | ( n_n100  &  wire274 ) | ( n_n100  &  _1433 ) ;
 assign _1429 = ( wire66  &  n_n100 ) | ( n_n100  &  _39740 ) ;
 assign _1430 = ( i_14_  &  i_13_  &  i_12_  &  wire903 ) ;
 assign _1433 = ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire903 ) ;
 assign _1473 = ( n_n48  &  wire56 ) | ( n_n48  &  wire104 ) | ( n_n48  &  _39690 ) ;
 assign _1497 = ( n_n48  &  wire52 ) | ( n_n48  &  wire247 ) | ( n_n48  &  _39670 ) ;
 assign _1498 = ( wire66  &  n_n53 ) | ( n_n53  &  wire343 ) | ( n_n53  &  _39674 ) ;
 assign _1509 = ( n_n57  &  wire78 ) | ( n_n57  &  wire342 ) | ( n_n57  &  _1512 ) ;
 assign _1510 = ( n_n57  &  wire64 ) | ( n_n57  &  wire102 ) | ( n_n57  &  _39657 ) ;
 assign _1512 = ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  wire901 ) ;
 assign _1515 = ( n_n56  &  wire102 ) | ( n_n56  &  wire342 ) | ( n_n56  &  _1518 ) ;
 assign _1516 = ( n_n56  &  wire55 ) | ( n_n56  &  wire19407 ) | ( n_n56  &  _39653 ) ;
 assign _1518 = ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire914 ) ;
 assign _1526 = ( n_n57  &  wire56 ) | ( n_n57  &  wire345 ) | ( n_n57  &  _1528 ) ;
 assign _1527 = ( n_n57  &  wire104 ) | ( n_n57  &  wire274 ) | ( n_n57  &  _1531 ) ;
 assign _1528 = ( i_14_  &  i_13_  &  i_12_  &  wire903 ) ;
 assign _1531 = ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire903 ) ;
 assign _1534 = ( n_n5  &  wire81 ) | ( n_n5  &  wire311 ) | ( n_n5  &  _1537 ) ;
 assign _1535 = ( n_n5  &  wire19578 ) | ( n_n5  &  wire300 ) | ( n_n5  &  _1540 ) ;
 assign _1537 = ( i_14_  &  i_13_  &  i_12_  &  wire906 ) ;
 assign _1540 = ( i_14_  &  i_13_  &  (~ i_12_)  &  wire906 ) ;
 assign _1580 = ( n_n285  &  n_n230  &  n_n263  &  wire998 ) ;
 assign _1583 = ( n_n6  &  wire56 ) | ( n_n6  &  wire104 ) | ( n_n6  &  _39601 ) ;
 assign _1584 = ( n_n285  &  n_n230  &  n_n261  &  wire345 ) ;
 assign _1588 = ( wire914  &  n_n6  &  _36202 ) ;
 assign _1591 = ( wire112  &  n_n5 ) | ( n_n5  &  wire77 ) | ( n_n5  &  _1593 ) ;
 assign _1592 = ( wire200  &  n_n5 ) | ( n_n5  &  wire807 ) | ( n_n5  &  _1596 ) ;
 assign _1593 = ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  wire898 ) ;
 assign _1596 = ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire904 ) ;
 assign _1599 = ( n_n6  &  wire55 ) | ( n_n6  &  wire87 ) | ( n_n6  &  _1602 ) ;
 assign _1602 = ( i_14_  &  i_13_  &  i_12_  &  wire914 ) ;
 assign _1614 = ( n_n6  &  wire78 ) | ( n_n6  &  wire433 ) | ( n_n6  &  _1617 ) ;
 assign _1617 = ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  wire901 ) ;
 assign _1626 = ( n_n48  &  wire68 ) | ( n_n48  &  wire19575 ) | ( n_n48  &  _39574 ) ;
 assign _1652 = ( n_n56  &  wire514 ) | ( n_n56  &  wire325 ) | ( n_n56  &  _1655 ) ;
 assign _1655 = ( (~ i_14_)  &  i_13_  &  i_12_  &  wire911 ) ;
 assign _1673 = ( n_n53  &  wire19575 ) | ( n_n53  &  wire22255 ) | ( n_n53  &  _1676 ) ;
 assign _1676 = ( (~ i_14_)  &  i_13_  &  i_12_  &  wire898 ) ;
 assign _1683 = ( wire273  &  n_n53 ) | ( n_n53  &  wire57 ) | ( n_n53  &  _39526 ) ;
 assign _1686 = ( wire64  &  n_n48 ) | ( n_n48  &  wire78 ) | ( n_n48  &  _39514 ) ;
 assign _1718 = ( n_n3  &  wire49 ) | ( n_n3  &  wire212 ) | ( n_n3  &  _1720 ) ;
 assign _1719 = ( n_n3  &  wire65 ) | ( n_n3  &  wire124 ) | ( n_n3  &  _1723 ) ;
 assign _1720 = ( i_14_  &  i_13_  &  i_12_  &  wire908 ) ;
 assign _1723 = ( (~ i_14_)  &  i_13_  &  i_12_  &  wire902 ) ;
 assign _1729 = ( n_n3  &  wire85 ) | ( n_n3  &  wire437 ) | ( n_n3  &  _1731 ) ;
 assign _1730 = ( n_n3  &  wire47 ) | ( n_n3  &  _39479 ) ;
 assign _1731 = ( i_14_  &  i_13_  &  i_12_  &  wire907 ) ;
 assign _1737 = ( n_n208  &  n_n284  &  n_n285  &  wire1491 ) ;
 assign _1743 = ( n_n3  &  wire67 ) | ( n_n3  &  wire245 ) | ( n_n3  &  _39461 ) ;
 assign _1744 = ( n_n229  &  n_n284  &  n_n285  &  wire347 ) ;
 assign _1760 = ( n_n3  &  wire84 ) | ( n_n3  &  wire62 ) | ( n_n3  &  _39441 ) ;
 assign _1796 = ( n_n3  &  wire51 ) | ( n_n3  &  wire19385 ) | ( n_n3  &  _39412 ) ;
 assign _1797 = ( n_n229  &  n_n284  &  n_n285  &  wire448 ) ;
 assign _1801 = ( n_n208  &  n_n284  &  n_n285  &  wire300 ) ;
 assign _1807 = ( n_n265  &  wire85 ) | ( n_n265  &  wire47 ) | ( n_n265  &  _39398 ) ;
 assign _1815 = ( n_n268  &  wire40 ) | ( n_n268  &  wire343 ) | ( n_n268  &  _1817 ) ;
 assign _1816 = ( n_n268  &  wire84 ) | ( n_n268  &  wire62 ) | ( n_n268  &  _39396 ) ;
 assign _1817 = ( i_14_  &  (~ i_13_)  &  i_12_  &  wire911 ) ;
 assign _1832 = ( n_n268  &  wire57 ) | ( n_n268  &  wire22002 ) | ( n_n268  &  _1835 ) ;
 assign _1835 = ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire914 ) ;
 assign _1843 = ( n_n4  &  wire154 ) | ( n_n4  &  wire64 ) | ( n_n4  &  _39379 ) ;
 assign _1853 = ( n_n3  &  wire104 ) | ( n_n3  &  wire228 ) | ( n_n3  &  _39375 ) ;
 assign _1861 = ( n_n3  &  wire143 ) | ( n_n3  &  _39369 ) ;
 assign _1889 = ( n_n3  &  wire84 ) | ( n_n3  &  _1895 ) | ( n_n3  &  _1896 ) ;
 assign _1892 = ( n_n4  &  wire84 ) | ( n_n4  &  _1895 ) | ( n_n4  &  _1896 ) ;
 assign _1895 = ( i_14_  &  i_13_  &  (~ i_12_)  &  _39347 ) ;
 assign _1896 = ( i_14_  &  i_13_  &  (~ i_12_)  &  _39348 ) ;
 assign _1898 = ( n_n6  &  wire64 ) | ( n_n6  &  wire61 ) | ( n_n6  &  _39338 ) ;
 assign _1903 = ( n_n5  &  wire102 ) | ( n_n5  &  wire263 ) | ( n_n5  &  _1906 ) ;
 assign _1906 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire912 ) ;
 assign _1909 = ( n_n5  &  wire104 ) | ( n_n5  &  wire228 ) | ( n_n5  &  _39334 ) ;
 assign _1934 = ( n_n5  &  wire143 ) | ( n_n5  &  wire375 ) | ( n_n5  &  _39322 ) ;
 assign _1952 = ( n_n5  &  wire84 ) | ( n_n5  &  n_n69 ) | ( n_n5  &  wire230 ) ;
 assign _1966 = ( n_n5  &  wire226 ) | ( n_n5  &  wire21668 ) | ( n_n5  &  _39296 ) ;
 assign _1967 = ( n_n5  &  wire807 ) | ( n_n5  &  wire270 ) | ( n_n5  &  _1968 ) ;
 assign _1968 = ( i_14_  &  i_13_  &  (~ i_12_)  &  wire904 ) ;
 assign _1997 = ( n_n48  &  wire143 ) | ( n_n48  &  wire195 ) | ( n_n48  &  _39275 ) ;
 assign _1998 = ( n_n48  &  wire84 ) | ( n_n48  &  n_n69 ) | ( n_n48  &  wire375 ) ;
 assign _2137 = ( n_n94  &  wire362 ) | ( n_n94  &  wire361 ) ;
 assign _2138 = ( n_n94  &  wire59 ) | ( n_n94  &  wire243 ) | ( n_n94  &  _2140 ) ;
 assign _2139 = ( n_n94  &  wire226 ) | ( wire898  &  n_n256  &  n_n94 ) ;
 assign _2140 = ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  wire906 ) ;
 assign _2145 = ( n_n100  &  wire87 ) | ( n_n100  &  wire428 ) | ( n_n100  &  _2147 ) ;
 assign _2146 = ( n_n100  &  wire59 ) | ( n_n100  &  wire243 ) | ( n_n100  &  _2150 ) ;
 assign _2147 = ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  wire914 ) ;
 assign _2150 = ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  wire906 ) ;
 assign _2215 = ( n_n48  &  wire104 ) | ( n_n48  &  wire228 ) | ( n_n48  &  _39109 ) ;
 assign _2220 = ( n_n264  &  n_n273  &  n_n285  &  wire1594 ) ;
 assign _2223 = ( n_n48  &  wire226 ) | ( n_n48  &  wire21668 ) | ( n_n48  &  _39100 ) ;
 assign _2224 = ( n_n48  &  wire807 ) | ( n_n48  &  wire270 ) | ( n_n48  &  _2225 ) ;
 assign _2225 = ( i_14_  &  i_13_  &  (~ i_12_)  &  wire904 ) ;
 assign _2230 = ( n_n53  &  wire807 ) | ( n_n53  &  wire226 ) | ( n_n53  &  _39097 ) ;
 assign _2235 = ( n_n2  &  wire59 ) | ( n_n2  &  wire243 ) | ( n_n2  &  _2237 ) ;
 assign _2236 = ( n_n2  &  wire154 ) | ( n_n2  &  wire64 ) | ( n_n2  &  _2240 ) ;
 assign _2237 = ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  wire906 ) ;
 assign _2240 = ( i_14_  &  i_13_  &  (~ i_12_)  &  wire907 ) ;
 assign _2306 = ( n_n2  &  wire226 ) | ( n_n2  &  wire362 ) | ( n_n2  &  _2308 ) ;
 assign _2307 = ( n_n2  &  wire154 ) | ( n_n2  &  wire361 ) | ( n_n2  &  _2314 ) ;
 assign _2308 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire898 ) ;
 assign _2314 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire901 ) ;
 assign _2337 = ( n_n1  &  wire154 ) | ( n_n1  &  wire74 ) | ( n_n1  &  _39007 ) ;
 assign _2346 = ( n_n2  &  wire74 ) | ( n_n2  &  wire87 ) | ( n_n2  &  _38986 ) ;
 assign _2347 = ( n_n260  &  n_n285  &  n_n283  &  wire428 ) ;
 assign _2348 = ( n_n260  &  n_n285  &  n_n283  &  wire424 ) ;
 assign _2403 = ( n_n284  &  n_n285  &  n_n271  &  wire1696 ) ;
 assign _2404 = ( n_n284  &  n_n285  &  n_n271  &  wire212 ) ;
 assign _2412 = ( n_n4  &  wire807 ) | ( n_n4  &  wire226 ) | ( n_n4  &  _38943 ) ;
 assign _2448 = ( wire103  &  n_n127 ) | ( n_n127  &  _38907 ) ;
 assign _2449 = ( wire54  &  n_n127 ) | ( n_n220  &  wire914  &  n_n127 ) ;
 assign _2458 = ( n_n48  &  wire80 ) | ( n_n48  &  _38892 ) ;
 assign _2459 = ( n_n48  &  wire40 ) | ( n_n48  &  wire21367 ) | ( n_n48  &  _2463 ) ;
 assign _2463 = ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  wire897 ) ;
 assign _2474 = ( n_n279  &  wire905  &  n_n53 ) ;
 assign _2475 = ( wire48  &  n_n53 ) | ( n_n53  &  wire62 ) | ( n_n53  &  _38877 ) ;
 assign _2476 = ( n_n279  &  wire899  &  n_n48 ) ;
 assign _2477 = ( wire48  &  n_n48 ) | ( n_n48  &  wire62 ) | ( n_n48  &  _38877 ) ;
 assign _2478 = ( wire79  &  n_n48 ) | ( n_n48  &  wire83 ) | ( n_n48  &  _38874 ) ;
 assign _2483 = ( wire54  &  n_n53 ) | ( n_n53  &  wire21596 ) | ( n_n53  &  _38870 ) ;
 assign _2486 = ( n_n48  &  wire77 ) | ( n_n48  &  wire86 ) | ( n_n48  &  _38867 ) ;
 assign _2487 = ( n_n48  &  wire71 ) | ( n_n48  &  wire78 ) | ( n_n48  &  _2488 ) ;
 assign _2488 = ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire904 ) ;
 assign _2498 = ( wire54  &  n_n6 ) | ( n_n6  &  wire21389 ) | ( n_n6  &  _38855 ) ;
 assign _2503 = ( n_n5  &  wire71 ) | ( n_n5  &  _38853 ) ;
 assign _2517 = ( wire54  &  n_n5 ) | ( n_n5  &  wire86 ) | ( n_n5  &  _38844 ) ;
 assign _2557 = ( n_n5  &  _38804 ) | ( n_n5  &  _38805 ) ;
 assign _2558 = ( n_n5  &  wire80 ) | ( n_n5  &  _38806 ) ;
 assign _2611 = ( wire48  &  n_n6 ) | ( n_n6  &  wire62 ) | ( n_n6  &  _38772 ) ;
 assign _2630 = ( n_n2  &  wire153 ) | ( n_n2  &  wire255 ) | ( n_n2  &  wire436 ) ;
 assign _2633 = ( n_n4  &  wire79 ) | ( n_n4  &  wire80 ) | ( n_n4  &  _38741 ) ;
 assign _2656 = ( n_n3  &  _38722 ) | ( n_n3  &  _38723 ) ;
 assign _2657 = ( n_n3  &  wire80 ) | ( n_n3  &  _38724 ) ;
 assign _2677 = ( wire48  &  n_n4 ) | ( n_n4  &  wire62 ) | ( n_n4  &  _38699 ) ;
 assign _2711 = ( n_n1  &  wire119 ) | ( n_n1  &  wire281 ) | ( n_n1  &  wire858 ) ;
 assign _2716 = ( n_n2  &  wire268 ) | ( n_n2  &  wire119 ) | ( n_n2  &  wire858 ) ;
 assign _2719 = ( n_n3  &  wire71 ) | ( n_n3  &  _38666 ) ;
 assign _2720 = ( n_n3  &  wire21389 ) | ( n_n281  &  n_n3  &  wire900 ) ;
 assign _2727 = ( wire54  &  n_n3 ) | ( n_n3  &  _38665 ) ;
 assign _2728 = ( n_n3  &  wire78 ) | ( n_n3  &  wire86 ) | ( n_n3  &  _38663 ) ;
 assign _2732 = ( n_n4  &  wire78 ) | ( n_n4  &  wire86 ) | ( n_n4  &  _38663 ) ;
 assign _2733 = ( n_n208  &  n_n284  &  n_n285  &  wire67 ) ;
 assign _2741 = ( wire54  &  n_n4 ) | ( n_n4  &  wire71 ) | ( n_n4  &  _38656 ) ;
 assign _2760 = ( n_n268  &  wire19738 ) | ( n_n268  &  wire19408 ) | ( n_n268  &  _38643 ) ;
 assign _2761 = ( n_n284  &  n_n285  &  n_n271  &  wire21383 ) ;
 assign _2766 = ( n_n268  &  wire453 ) | ( n_n268  &  wire21379 ) | ( n_n268  &  _38640 ) ;
 assign _2793 = ( n_n94  &  wire327 ) | ( n_n94  &  wire235 ) | ( n_n94  &  wire21474 ) ;
 assign _2854 = ( n_n53  &  _38550 ) | ( n_n53  &  _38551 ) ;
 assign _2888 = ( n_n56  &  wire453 ) | ( n_n56  &  wire329 ) | ( n_n56  &  _2891 ) ;
 assign _2891 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire914 ) ;
 assign _2946 = ( n_n228  &  n_n57  &  wire899 ) ;
 assign _2959 = ( n_n56  &  wire73 ) | ( n_n56  &  wire469 ) | ( n_n56  &  _38452 ) ;
 assign _2960 = ( n_n56  &  wire79 ) | ( n_n56  &  wire83 ) | ( n_n56  &  _2962 ) ;
 assign _2961 = ( n_n56  &  wire66 ) | ( wire905  &  n_n56  &  n_n222 ) ;
 assign _2962 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire899 ) ;
 assign _2965 = ( n_n57  &  wire199 ) | ( n_n57  &  wire113 ) | ( n_n57  &  _38448 ) ;
 assign _2976 = ( wire95  &  n_n56 ) | ( n_n56  &  wire101 ) | ( n_n56  &  _2979 ) ;
 assign _2979 = ( i_14_  &  i_13_  &  i_12_  &  wire912 ) ;
 assign _2982 = ( n_n57  &  wire514 ) | ( n_n57  &  wire20155 ) | ( n_n57  &  _38437 ) ;
 assign _2983 = ( n_n57  &  wire20149 ) | ( n_n57  &  _38439 ) ;
 assign _2984 = ( n_n56  &  wire514 ) | ( n_n56  &  wire20155 ) | ( n_n56  &  _38437 ) ;
 assign _2985 = ( n_n56  &  wire20149 ) | ( n_n56  &  _38439 ) ;
 assign _2992 = ( n_n56  &  wire88 ) | ( n_n56  &  wire80 ) | ( n_n56  &  _38430 ) ;
 assign _2993 = ( n_n56  &  wire65 ) | ( n_n56  &  _38432 ) ;
 assign _3000 = ( n_n57  &  wire469 ) | ( n_n57  &  wire74 ) | ( n_n57  &  _38426 ) ;
 assign _3001 = ( n_n57  &  wire79 ) | ( n_n57  &  wire40 ) | ( n_n57  &  _3003 ) ;
 assign _3002 = ( n_n57  &  wire66 ) | ( wire905  &  n_n57  &  n_n222 ) ;
 assign _3003 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire899 ) ;
 assign _3006 = ( n_n57  &  wire86 ) | ( n_n57  &  wire47 ) | ( n_n57  &  _38421 ) ;
 assign _3007 = ( n_n57  &  wire88 ) | ( n_n57  &  wire89 ) | ( n_n57  &  _38423 ) ;
 assign _3008 = ( n_n57  &  wire78 ) | ( wire902  &  n_n258  &  n_n57 ) ;
 assign _3011 = ( n_n56  &  wire67 ) | ( n_n56  &  n_n41 ) | ( n_n56  &  _38418 ) ;
 assign _3012 = ( n_n56  &  wire102 ) | ( n_n56  &  wire87 ) | ( n_n56  &  _38419 ) ;
 assign _3013 = ( n_n56  &  wire104 ) | ( n_n56  &  wire74 ) | ( n_n56  &  _38413 ) ;
 assign _3014 = ( n_n56  &  wire40 ) | ( n_n56  &  wire19457 ) | ( n_n56  &  _3016 ) ;
 assign _3016 = ( i_14_  &  i_13_  &  (~ i_12_)  &  wire897 ) ;
 assign _3021 = ( n_n57  &  wire80 ) | ( n_n57  &  wire19457 ) | ( n_n57  &  _38409 ) ;
 assign _3022 = ( n_n57  &  wire65 ) | ( n_n57  &  _38411 ) ;
 assign _3023 = ( n_n57  &  wire104 ) | ( n_n279  &  n_n57  &  wire903 ) ;
 assign _3027 = ( n_n57  &  _38403 ) | ( n_n57  &  _38404 ) ;
 assign _3028 = ( n_n57  &  wire19578 ) | ( n_n57  &  _38405 ) ;
 assign _3035 = ( n_n56  &  wire59 ) | ( n_n56  &  wire19575 ) | ( n_n56  &  _38399 ) ;
 assign _3036 = ( n_n56  &  wire51 ) | ( n_n56  &  wire71 ) | ( n_n56  &  _3038 ) ;
 assign _3037 = ( n_n56  &  wire96 ) | ( n_n56  &  wire898  &  n_n222 ) ;
 assign _3038 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire898 ) ;
 assign _3041 = ( n_n57  &  wire67 ) | ( n_n57  &  n_n41 ) | ( n_n57  &  _38394 ) ;
 assign _3042 = ( n_n57  &  wire102 ) | ( n_n57  &  wire87 ) | ( n_n57  &  _38395 ) ;
 assign _3043 = ( n_n56  &  wire86 ) | ( n_n56  &  wire47 ) | ( n_n56  &  _38390 ) ;
 assign _3044 = ( n_n56  &  wire89 ) | ( n_n56  &  _38392 ) ;
 assign _3058 = ( n_n56  &  wire19578 ) | ( n_n56  &  _38380 ) ;
 assign _3064 = ( n_n57  &  wire71 ) | ( n_n57  &  wire96 ) | ( n_n57  &  _3067 ) ;
 assign _3067 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire898 ) ;
 assign _3070 = ( (~ i_14_)  &  i_13_  &  i_12_  &  wire898 ) ;
 assign _3077 = ( n_n3  &  _38368 ) | ( n_n3  &  _38369 ) ;
 assign _3078 = ( n_n3  &  wire19578 ) | ( n_n3  &  _38370 ) ;
 assign _3082 = ( n_n4  &  wire71 ) | ( n_n4  &  wire19575 ) | ( n_n4  &  _38365 ) ;
 assign _3094 = ( n_n268  &  wire57 ) | ( n_n268  &  wire20107 ) | ( n_n268  &  _38355 ) ;
 assign _3095 = ( n_n268  &  wire453 ) | ( n_n268  &  wire245 ) | ( n_n268  &  _38357 ) ;
 assign _3096 = ( n_n268  &  wire50 ) | ( n_n268  &  wire21271 ) ;
 assign _3101 = ( n_n265  &  wire89 ) | ( n_n265  &  wire86 ) | ( n_n265  &  _38348 ) ;
 assign _3102 = ( n_n265  &  wire64 ) | ( n_n265  &  wire85 ) | ( n_n265  &  _3103 ) ;
 assign _3103 = ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire907 ) ;
 assign _3106 = ( n_n268  &  wire84 ) | ( n_n268  &  wire52 ) | ( n_n268  &  _38345 ) ;
 assign _3107 = ( n_n268  &  wire19738 ) | ( n_n268  &  wire60 ) | ( n_n268  &  _3108 ) ;
 assign _3108 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire913 ) ;
 assign _3124 = ( n_n268  &  wire19407 ) | ( n_n268  &  wire53 ) | ( n_n268  &  _38328 ) ;
 assign _3132 = ( wire905  &  n_n4  &  n_n256 ) ;
 assign _3173 = ( n_n3  &  wire66 ) | ( n_n3  &  wire20155 ) | ( n_n3  &  _38289 ) ;
 assign _3174 = ( n_n3  &  wire79 ) | ( n_n3  &  wire469 ) | ( n_n3  &  _38291 ) ;
 assign _3175 = ( n_n3  &  wire62 ) | ( n_n258  &  n_n3  &  wire899 ) ;
 assign _3178 = ( n_n4  &  wire62 ) | ( n_n4  &  wire20155 ) | ( n_n4  &  _38285 ) ;
 assign _3179 = ( n_n4  &  wire514 ) | ( n_n4  &  wire20149 ) | ( n_n4  &  _38287 ) ;
 assign _3180 = ( n_n4  &  wire19457 ) | ( n_n4  &  wire74 ) | ( n_n4  &  _38274 ) ;
 assign _3181 = ( n_n4  &  wire104 ) | ( n_n279  &  n_n4  &  wire903 ) ;
 assign _3182 = ( n_n208  &  n_n284  &  n_n285  &  wire40 ) ;
 assign _3187 = ( n_n3  &  wire80 ) | ( n_n3  &  wire20149 ) | ( n_n3  &  _38277 ) ;
 assign _3188 = ( n_n3  &  wire69 ) | ( n_n3  &  wire65 ) | ( n_n3  &  _3190 ) ;
 assign _3189 = ( n_n3  &  wire514 ) | ( wire911  &  n_n3  &  n_n225 ) ;
 assign _3190 = ( (~ i_14_)  &  i_13_  &  i_12_  &  wire902 ) ;
 assign _3195 = ( n_n3  &  wire88 ) | ( n_n3  &  _38273 ) ;
 assign _3196 = ( n_n3  &  wire19457 ) | ( n_n3  &  wire74 ) | ( n_n3  &  _38274 ) ;
 assign _3197 = ( n_n3  &  wire104 ) | ( n_n279  &  n_n3  &  wire903 ) ;
 assign _3206 = ( n_n4  &  wire102 ) | ( n_n4  &  wire368 ) | ( n_n4  &  _38266 ) ;
 assign _3211 = ( n_n3  &  wire71 ) | ( n_n3  &  wire19575 ) | ( n_n3  &  _38118 ) ;
 assign _3216 = ( n_n4  &  wire87 ) | ( n_n4  &  _38260 ) ;
 assign _3217 = ( n_n4  &  wire86 ) | ( n_n4  &  wire47 ) | ( n_n4  &  _38256 ) ;
 assign _3218 = ( n_n4  &  wire89 ) | ( n_n4  &  _38258 ) ;
 assign _3222 = ( n_n3  &  wire86 ) | ( n_n3  &  wire47 ) | ( n_n3  &  _38256 ) ;
 assign _3223 = ( n_n3  &  wire89 ) | ( n_n3  &  _38258 ) ;
 assign _3235 = ( n_n3  &  wire67 ) | ( n_n3  &  n_n103 ) | ( n_n3  &  _38248 ) ;
 assign _3236 = ( n_n3  &  wire102 ) | ( n_n3  &  wire87 ) | ( n_n3  &  _38249 ) ;
 assign _3260 = ( wire48  &  n_n127 ) | ( wire54  &  n_n127 ) | ( n_n127  &  _38211 ) ;
 assign _3263 = ( wire54  &  n_n132 ) | ( wire54  &  _3271 ) | ( n_n132  &  _38208 ) | ( _3271  &  _38208 ) ;
 assign _3271 = ( n_n229  &  n_n165  &  n_n284 ) ;
 assign _3294 = ( n_n2  &  wire44 ) | ( n_n2  &  wire160 ) | ( n_n2  &  _38187 ) ;
 assign _3295 = ( n_n1  &  wire95 ) | ( n_n1  &  wire44 ) | ( n_n1  &  _38189 ) ;
 assign _3296 = ( n_n2  &  wire66 ) | ( n_n2  &  wire42 ) | ( n_n2  &  _36256 ) ;
 assign _3300 = ( n_n3  &  wire96 ) | ( n_n3  &  wire807 ) | ( n_n3  &  _35454 ) ;
 assign _3311 = ( n_n2  &  wire72 ) | ( n_n2  &  wire184 ) | ( n_n2  &  _3314 ) ;
 assign _3314 = ( i_14_  &  (~ i_13_)  &  i_12_  &  wire905 ) ;
 assign _3319 = ( n_n3  &  wire66 ) | ( n_n3  &  wire79 ) | ( n_n3  &  _38167 ) ;
 assign _3320 = ( n_n3  &  wire42 ) | ( n_n3  &  _38169 ) ;
 assign _3324 = ( n_n4  &  wire453 ) | ( n_n4  &  wire55 ) | ( n_n4  &  _3330 ) ;
 assign _3327 = ( n_n3  &  wire453 ) | ( n_n3  &  wire55 ) | ( n_n3  &  _3330 ) ;
 assign _3328 = ( n_n3  &  wire57 ) | ( n_n279  &  wire912  &  n_n3 ) ;
 assign _3329 = ( n_n3  &  wire245 ) | ( wire912  &  n_n3  &  n_n225 ) ;
 assign _3330 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire914 ) ;
 assign _3333 = ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire912 ) ;
 assign _3343 = ( n_n3  &  wire88 ) | ( n_n3  &  wire80 ) | ( n_n3  &  _38157 ) ;
 assign _3344 = ( n_n5  &  wire66 ) | ( n_n5  &  wire469 ) | ( n_n5  &  _37064 ) ;
 assign _3358 = ( wire49  &  n_n227 ) | ( n_n227  &  wire143 ) | ( n_n227  &  _38138 ) ;
 assign _3384 = ( n_n3  &  wire71 ) | ( n_n3  &  wire19575 ) | ( n_n3  &  _38118 ) ;
 assign _3396 = ( n_n2  &  wire96 ) | ( n_n2  &  wire807 ) | ( n_n2  &  _35352 ) ;
 assign _3400 = ( n_n2  &  wire80 ) | ( n_n2  &  wire61 ) | ( n_n2  &  _35370 ) ;
 assign _3408 = ( n_n2  &  wire453 ) | ( n_n2  &  wire55 ) | ( n_n2  &  _3411 ) ;
 assign _3411 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire914 ) ;
 assign _3414 = ( wire914  &  n_n57  &  _34952 ) ;
 assign _3423 = ( n_n56  &  wire66 ) | ( n_n56  &  wire79 ) | ( n_n56  &  _36518 ) ;
 assign _3424 = ( n_n56  &  wire44 ) | ( n_n56  &  _38083 ) ;
 assign _3430 = ( n_n94  &  wire96 ) | ( n_n94  &  wire19575 ) | ( n_n94  &  _35700 ) ;
 assign _3443 = ( wire80  &  n_n100 ) | ( n_n100  &  wire69 ) | ( n_n100  &  _3446 ) ;
 assign _3444 = ( wire88  &  n_n100 ) | ( n_n100  &  wire65 ) | ( n_n100  &  _35652 ) ;
 assign _3446 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire902 ) ;
 assign _3449 = ( wire67  &  n_n94 ) | ( n_n94  &  wire65 ) | ( n_n94  &  _3452 ) ;
 assign _3452 = ( (~ i_14_)  &  i_13_  &  i_12_  &  wire902 ) ;
 assign _3472 = ( wire66  &  n_n94 ) | ( n_n94  &  wire469 ) | ( n_n94  &  _37753 ) ;
 assign _3498 = ( wire44  &  n_n48 ) | ( wire79  &  n_n48 ) | ( n_n48  &  _38020 ) ;
 assign _3503 = ( wire66  &  n_n48 ) | ( n_n48  &  wire42 ) | ( n_n48  &  _37834 ) ;
 assign _3512 = ( wire912  &  n_n256  &  n_n48 ) ;
 assign _3529 = ( n_n48  &  wire96 ) | ( n_n48  &  wire807 ) | ( n_n48  &  _35178 ) ;
 assign _3547 = ( n_n5  &  wire80 ) | ( n_n5  &  wire65 ) | ( n_n5  &  _37037 ) ;
 assign _3550 = ( n_n5  &  wire96 ) | ( n_n5  &  wire19575 ) | ( n_n5  &  _37027 ) ;
 assign _3566 = ( wire48  &  n_n132 ) | ( wire103  &  n_n132 ) | ( n_n132  &  _37969 ) ;
 assign _3567 = ( wire54  &  n_n132 ) | ( n_n220  &  wire914  &  n_n132 ) ;
 assign _3570 = ( n_n264  &  n_n229  &  n_n165  &  _37961 ) ;
 assign _3589 = ( n_n1  &  wire96 ) | ( n_n1  &  wire807 ) | ( n_n1  &  _35428 ) ;
 assign _3597 = ( n_n268  &  wire210 ) | ( n_n268  &  wire130 ) | ( n_n268  &  _3599 ) ;
 assign _3598 = ( n_n268  &  wire60 ) | ( n_n268  &  wire52 ) | ( n_n268  &  _37922 ) ;
 assign _3599 = ( i_14_  &  i_13_  &  i_12_  &  wire911 ) ;
 assign _3602 = ( n_n2  &  wire72 ) | ( n_n2  &  _37919 ) ;
 assign _3628 = ( n_n3  &  wire60 ) | ( n_n3  &  wire52 ) | ( n_n3  &  _37905 ) ;
 assign _3629 = ( n_n3  &  wire19738 ) | ( n_n3  &  wire84 ) | ( n_n3  &  _37907 ) ;
 assign _3636 = ( n_n3  &  wire66 ) | ( n_n3  &  wire42 ) | ( n_n3  &  _37899 ) ;
 assign _3674 = ( n_n1  &  wire66 ) | ( n_n1  &  wire79 ) | ( n_n1  &  _36265 ) ;
 assign _3675 = ( n_n1  &  wire42 ) | ( n_n1  &  _37860 ) ;
 assign _3679 = ( n_n2  &  wire71 ) | ( n_n2  &  _37859 ) ;
 assign _3680 = ( n_n2  &  wire96 ) | ( n_n2  &  wire807 ) | ( n_n2  &  _35352 ) ;
 assign _3692 = ( n_n2  &  wire19738 ) | ( n_n2  &  wire42 ) | ( n_n2  &  _37849 ) ;
 assign _3695 = ( n_n2  &  wire84 ) | ( n_n2  &  wire52 ) | ( n_n2  &  _36270 ) ;
 assign _3708 = ( wire66  &  n_n48 ) | ( n_n48  &  wire42 ) | ( n_n48  &  _37834 ) ;
 assign _3718 = ( n_n48  &  wire84 ) | ( n_n48  &  _37830 ) ;
 assign _3719 = ( wire19738  &  n_n48 ) | ( n_n48  &  wire52 ) | ( n_n48  &  _37828 ) ;
 assign _3723 = ( wire19738  &  n_n53 ) | ( n_n53  &  wire52 ) | ( n_n53  &  _37828 ) ;
 assign _3724 = ( n_n264  &  n_n273  &  n_n285  &  wire60 ) ;
 assign _3786 = ( wire66  &  n_n94 ) | ( n_n94  &  wire469 ) | ( n_n94  &  _37753 ) ;
 assign _3787 = ( n_n100  &  wire514 ) | ( n_n100  &  wire20155 ) | ( n_n100  &  _37755 ) ;
 assign _3833 = ( n_n5  &  wire64 ) | ( n_n5  &  wire89 ) | ( n_n5  &  _36116 ) ;
 assign _3834 = ( n_n285  &  n_n230  &  n_n263  &  wire99 ) ;
 assign _3852 = ( n_n285  &  n_n266  &  n_n230  &  wire140 ) ;
 assign _3878 = ( n_n56  &  wire66 ) | ( n_n56  &  wire79 ) | ( n_n56  &  _36518 ) ;
 assign _3896 = ( n_n260  &  n_n285  &  n_n271  &  wire950 ) ;
 assign _3920 = ( (~ i_7_)  &  (~ i_6_)  &  n_n264  &  n_n118 ) ;
 assign _3973 = ( n_n4  &  wire88 ) | ( n_n4  &  wire61 ) | ( n_n4  &  _37568 ) ;
 assign _3979 = ( n_n4  &  wire70 ) | ( n_n4  &  wire19738 ) | ( n_n4  &  _37562 ) ;
 assign _3980 = ( n_n4  &  wire42 ) | ( n_n279  &  n_n4  &  wire899 ) ;
 assign _3988 = ( n_n4  &  wire60 ) | ( n_n4  &  wire84 ) | ( n_n4  &  _3991 ) ;
 assign _3991 = ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire913 ) ;
 assign _4005 = ( n_n1  &  wire118 ) | ( n_n1  &  wire50 ) | ( n_n1  &  _37535 ) ;
 assign _4006 = ( wire75  &  n_n1 ) | ( n_n1  &  wire20593 ) | ( n_n1  &  _4008 ) ;
 assign _4007 = ( n_n1  &  wire72 ) | ( n_n1  &  wire113 ) ;
 assign _4008 = ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  wire913 ) ;
 assign _4013 = ( n_n1  &  wire70 ) | ( n_n1  &  wire73 ) | ( n_n1  &  _37530 ) ;
 assign _4014 = ( n_n1  &  wire95 ) | ( n_n1  &  wire101 ) | ( n_n1  &  _37532 ) ;
 assign _4015 = ( n_n1  &  wire44 ) | ( n_n228  &  n_n1  &  wire900 ) ;
 assign _4018 = ( n_n4  &  wire76 ) | ( n_n4  &  wire19385 ) | ( n_n4  &  _35456 ) ;
 assign _4028 = ( n_n4  &  wire96 ) | ( n_n4  &  wire807 ) | ( n_n4  &  _37525 ) ;
 assign _4031 = ( n_n1  &  wire53 ) | ( n_n1  &  _37516 ) ;
 assign _4032 = ( n_n1  &  wire82 ) | ( n_n1  &  wire19408 ) | ( n_n1  &  _37517 ) ;
 assign _4039 = ( n_n1  &  wire96 ) | ( n_n1  &  wire807 ) | ( n_n1  &  _35428 ) ;
 assign _4040 = ( n_n1  &  wire71 ) | ( n_n1  &  n_n256  &  wire904 ) ;
 assign _4041 = ( n_n1  &  wire76 ) | ( n_n1  &  n_n279  &  wire900 ) ;
 assign _4044 = ( n_n1  &  wire55 ) | ( n_n1  &  wire19385 ) | ( n_n1  &  _37509 ) ;
 assign _4045 = ( n_n1  &  wire57 ) | ( n_n1  &  wire19384 ) | ( n_n1  &  _37511 ) ;
 assign _4046 = ( n_n1  &  wire81 ) | ( n_n220  &  n_n1  &  wire904 ) ;
 assign _4139 = ( wire56  &  n_n207 ) | ( n_n207  &  wire20362 ) | ( n_n207  &  _37445 ) ;
 assign _4147 = ( n_n6  &  wire62 ) | ( n_n6  &  wire20155 ) | ( n_n6  &  _37433 ) ;
 assign _4148 = ( n_n6  &  wire44 ) | ( n_n6  &  wire514 ) | ( n_n6  &  _37435 ) ;
 assign _4149 = ( n_n6  &  wire66 ) | ( n_n6  &  wire469 ) | ( n_n6  &  _37047 ) ;
 assign _4155 = ( n_n57  &  wire82 ) | ( n_n57  &  wire53 ) | ( n_n57  &  _37424 ) ;
 assign _4156 = ( n_n57  &  wire19407 ) | ( n_n57  &  _37426 ) ;
 assign _4160 = ( n_n220  &  n_n57  &  wire908 ) ;
 assign _4161 = ( n_n57  &  wire80 ) | ( n_n57  &  wire61 ) | ( n_n57  &  _35563 ) ;
 assign _4165 = ( n_n57  &  wire70 ) | ( n_n57  &  wire44 ) | ( n_n57  &  _37416 ) ;
 assign _4166 = ( n_n57  &  wire73 ) | ( n_n57  &  wire60 ) | ( n_n57  &  _4167 ) ;
 assign _4167 = ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  wire906 ) ;
 assign _4170 = ( n_n57  &  wire64 ) | ( n_n57  &  wire89 ) | ( n_n57  &  _36876 ) ;
 assign _4177 = ( n_n57  &  wire245 ) | ( n_n57  &  wire57 ) | ( n_n57  &  _37409 ) ;
 assign _4180 = ( n_n100  &  wire104 ) | ( n_n100  &  wire74 ) | ( n_n100  &  _35635 ) ;
 assign _4189 = ( i_14_  &  (~ i_13_)  &  i_12_  &  wire899 ) ;
 assign _4209 = ( wire71  &  n_n100 ) | ( n_n100  &  wire19575 ) | ( n_n100  &  _35712 ) ;
 assign _4210 = ( n_n100  &  wire96 ) | ( wire898  &  n_n222  &  n_n100 ) ;
 assign _4219 = ( n_n100  &  wire59 ) | ( n_n100  &  wire86 ) | ( n_n100  &  _37382 ) ;
 assign _4220 = ( n_n100  &  wire368 ) | ( n_n100  &  n_n88 ) | ( n_n100  &  wire20527 ) ;
 assign _4221 = ( wire51  &  n_n100 ) | ( wire907  &  n_n222  &  n_n100 ) ;
 assign _4226 = ( n_n100  &  wire87 ) | ( n_n100  &  _37380 ) ;
 assign _4249 = ( n_n100  &  wire514 ) | ( n_n100  &  wire20155 ) | ( n_n100  &  _37361 ) ;
 assign _4252 = ( wire66  &  n_n100 ) | ( wire79  &  n_n100 ) | ( n_n100  &  _37358 ) ;
 assign _4260 = ( n_n57  &  wire19385 ) | ( n_n57  &  wire19384 ) | ( n_n57  &  _35572 ) ;
 assign _4263 = ( n_n53  &  wire19407 ) | ( n_n53  &  wire19408 ) | ( n_n53  &  _35125 ) ;
 assign _4264 = ( n_n53  &  wire56 ) | ( n_n53  &  wire53 ) | ( n_n53  &  _37346 ) ;
 assign _4271 = ( wire70  &  n_n53 ) | ( wire44  &  n_n53 ) | ( n_n53  &  _37333 ) ;
 assign _4272 = ( wire73  &  n_n53 ) | ( n_n53  &  wire52 ) | ( n_n53  &  _37335 ) ;
 assign _4273 = ( wire19738  &  n_n53 ) | ( wire60  &  n_n53 ) | ( n_n53  &  _4274 ) ;
 assign _4274 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire913 ) ;
 assign _4277 = ( wire64  &  n_n53 ) | ( n_n53  &  wire89 ) | ( n_n53  &  _37300 ) ;
 assign _4295 = ( n_n53  &  wire55 ) | ( n_n53  &  wire57 ) | ( n_n53  &  _37314 ) ;
 assign _4296 = ( n_n53  &  _37316 ) | ( n_n53  &  _37317 ) ;
 assign _4297 = ( n_n53  &  wire81 ) | ( n_n220  &  wire904  &  n_n53 ) ;
 assign _4300 = ( n_n53  &  wire96 ) | ( n_n53  &  wire807 ) | ( n_n53  &  _35148 ) ;
 assign _4301 = ( n_n53  &  wire19385 ) | ( n_n256  &  wire900  &  n_n53 ) ;
 assign _4302 = ( n_n53  &  wire71 ) | ( n_n256  &  wire904  &  n_n53 ) ;
 assign _4310 = ( wire118  &  n_n57 ) | ( n_n57  &  wire50 ) | ( n_n57  &  _37304 ) ;
 assign _4311 = ( n_n57  &  wire101 ) | ( n_n57  &  wire20463 ) | ( n_n57  &  _4313 ) ;
 assign _4312 = ( wire72  &  n_n57 ) | ( n_n57  &  wire113 ) ;
 assign _4313 = ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  wire914 ) ;
 assign _4318 = ( wire64  &  n_n53 ) | ( n_n53  &  wire89 ) | ( n_n53  &  _37300 ) ;
 assign _4324 = ( n_n53  &  wire453 ) | ( n_n53  &  _37297 ) ;
 assign _4342 = ( n_n6  &  wire96 ) | ( n_n6  &  wire19575 ) | ( n_n6  &  _36964 ) ;
 assign _4348 = ( n_n6  &  wire104 ) | ( n_n6  &  wire74 ) | ( n_n6  &  _37072 ) ;
 assign _4349 = ( n_n6  &  wire88 ) | ( n_n6  &  _37280 ) ;
 assign _4357 = ( n_n6  &  wire89 ) | ( n_n6  &  wire47 ) | ( n_n6  &  _37000 ) ;
 assign _4362 = ( n_n6  &  wire59 ) | ( n_n6  &  wire86 ) | ( n_n6  &  _37273 ) ;
 assign _4365 = ( n_n53  &  _37226 ) | ( n_n53  &  _37227 ) ;
 assign _4366 = ( n_n53  &  wire19578 ) | ( n_n53  &  _37228 ) ;
 assign _4370 = ( n_n48  &  wire96 ) | ( n_n48  &  wire59 ) | ( n_n48  &  _37222 ) ;
 assign _4371 = ( n_n48  &  wire71 ) | ( n_n48  &  wire19575 ) | ( n_n48  &  _37224 ) ;
 assign _4376 = ( n_n48  &  wire86 ) | ( n_n48  &  wire20307 ) | ( n_n48  &  _4378 ) ;
 assign _4377 = ( n_n48  &  wire89 ) | ( n_n48  &  wire47 ) | ( n_n48  &  _37215 ) ;
 assign _4378 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire901 ) ;
 assign _4385 = ( n_n53  &  wire102 ) | ( n_n53  &  wire87 ) | ( n_n53  &  _37209 ) ;
 assign _4390 = ( n_n48  &  wire19578 ) | ( n_n48  &  wire19577 ) | ( n_n48  &  _37204 ) ;
 assign _4401 = ( n_n53  &  wire71 ) | ( n_n53  &  wire19575 ) | ( n_n53  &  _37189 ) ;
 assign _4412 = ( wire44  &  n_n48 ) | ( n_n48  &  wire469 ) | ( n_n48  &  _37178 ) ;
 assign _4413 = ( wire79  &  n_n48 ) | ( n_n48  &  _37180 ) ;
 assign _4414 = ( wire66  &  n_n48 ) | ( wire905  &  n_n222  &  n_n48 ) ;
 assign _4426 = ( n_n48  &  wire514 ) | ( n_n48  &  wire20149 ) | ( n_n48  &  _37168 ) ;
 assign _4429 = ( n_n53  &  wire514 ) | ( n_n53  &  wire20149 ) | ( n_n53  &  _37168 ) ;
 assign _4432 = ( (~ i_14_)  &  i_13_  &  i_12_  &  wire913 ) ;
 assign _4456 = ( n_n53  &  wire19457 ) | ( n_n53  &  wire104 ) | ( n_n53  &  _37148 ) ;
 assign _4457 = ( n_n53  &  wire65 ) | ( wire902  &  n_n225  &  n_n53 ) ;
 assign _4469 = ( n_n48  &  wire19457 ) | ( n_n48  &  wire74 ) | ( n_n48  &  _37141 ) ;
 assign _4485 = ( n_n48  &  wire80 ) | ( n_n48  &  wire65 ) | ( n_n48  &  _37128 ) ;
 assign _4514 = ( wire88  &  n_n53 ) | ( n_n53  &  wire61 ) | ( n_n53  &  _35213 ) ;
 assign _4559 = ( n_n5  &  n_n259  &  _34638 ) | ( n_n5  &  n_n259  &  _34639 ) ;
 assign _4567 = ( n_n5  &  wire73 ) | ( n_n5  &  wire44 ) | ( n_n5  &  _37097 ) ;
 assign _4574 = ( n_n6  &  wire95 ) | ( n_n6  &  wire256 ) | ( n_n6  &  _4577 ) ;
 assign _4577 = ( i_14_  &  i_13_  &  i_12_  &  wire912 ) ;
 assign _4582 = ( n_n6  &  wire113 ) | ( n_n6  &  wire50 ) | ( n_n6  &  _37087 ) ;
 assign _4585 = ( n_n5  &  wire95 ) | ( n_n5  &  wire50 ) | ( n_n5  &  _37084 ) ;
 assign _4596 = ( n_n6  &  wire104 ) | ( n_n6  &  wire74 ) | ( n_n6  &  _37072 ) ;
 assign _4599 = ( n_n5  &  wire40 ) | ( n_n5  &  wire104 ) | ( n_n5  &  _37068 ) ;
 assign _4600 = ( n_n5  &  wire19457 ) | ( n_n5  &  wire74 ) | ( n_n5  &  _37070 ) ;
 assign _4605 = ( n_n5  &  wire66 ) | ( n_n5  &  wire469 ) | ( n_n5  &  _37064 ) ;
 assign _4609 = ( n_n6  &  wire20149 ) | ( n_n6  &  _37063 ) ;
 assign _4610 = ( n_n6  &  wire514 ) | ( n_n6  &  wire20155 ) | ( n_n6  &  _37057 ) ;
 assign _4614 = ( n_n5  &  wire514 ) | ( n_n5  &  wire20155 ) | ( n_n5  &  _37057 ) ;
 assign _4615 = ( n_n285  &  n_n230  &  n_n263  &  wire62 ) ;
 assign _4622 = ( n_n6  &  wire66 ) | ( n_n6  &  wire469 ) | ( n_n6  &  _37047 ) ;
 assign _4631 = ( n_n5  &  wire80 ) | ( n_n5  &  wire65 ) | ( n_n5  &  _37037 ) ;
 assign _4635 = ( n_n5  &  wire88 ) | ( n_n5  &  _37032 ) ;
 assign _4643 = ( n_n5  &  wire96 ) | ( n_n5  &  wire19575 ) | ( n_n5  &  _37027 ) ;
 assign _4653 = ( n_n6  &  wire19578 ) | ( n_n6  &  wire19577 ) | ( n_n6  &  _37024 ) ;
 assign _4675 = ( n_n6  &  wire88 ) | ( n_n6  &  _37003 ) ;
 assign _4681 = ( n_n6  &  wire89 ) | ( n_n6  &  wire47 ) | ( n_n6  &  _37000 ) ;
 assign _4687 = ( n_n5  &  wire86 ) | ( n_n5  &  wire47 ) | ( n_n5  &  _36993 ) ;
 assign _4688 = ( n_n5  &  wire89 ) | ( n_n5  &  _36995 ) ;
 assign _4694 = ( n_n6  &  wire102 ) | ( n_n6  &  wire87 ) | ( n_n6  &  _36982 ) ;
 assign _4701 = ( n_n5  &  wire51 ) | ( n_n5  &  wire59 ) | ( n_n5  &  _36967 ) ;
 assign _4702 = ( n_n5  &  wire19578 ) | ( n_n5  &  wire19577 ) | ( n_n5  &  _36969 ) ;
 assign _4706 = ( n_n6  &  wire96 ) | ( n_n6  &  wire19575 ) | ( n_n6  &  _36964 ) ;
 assign _4769 = ( n_n56  &  wire66 ) | ( n_n56  &  wire79 ) | ( n_n56  &  _36518 ) ;
 assign _4771 = ( n_n285  &  n_n266  &  n_n230  &  wire44 ) ;
 assign _4775 = ( n_n56  &  wire84 ) | ( n_n56  &  wire52 ) | ( n_n56  &  _36895 ) ;
 assign _4777 = ( n_n56  &  wire76 ) | ( n_n56  &  wire19385 ) | ( n_n56  &  _36890 ) ;
 assign _4778 = ( n_n56  &  wire19384 ) | ( n_n281  &  n_n56  &  wire900 ) ;
 assign _4782 = ( n_n57  &  wire19385 ) | ( n_n57  &  wire19384 ) | ( n_n57  &  _35572 ) ;
 assign _4792 = ( n_n56  &  wire245 ) | ( n_n56  &  wire55 ) | ( n_n56  &  _4795 ) ;
 assign _4795 = ( (~ i_14_)  &  i_13_  &  i_12_  &  wire912 ) ;
 assign _4798 = ( n_n57  &  wire64 ) | ( n_n57  &  wire89 ) | ( n_n57  &  _36876 ) ;
 assign _4799 = ( n_n56  &  wire64 ) | ( n_n56  &  wire86 ) | ( n_n56  &  _36878 ) ;
 assign _4811 = ( n_n57  &  wire245 ) | ( n_n57  &  wire55 ) | ( n_n57  &  _4814 ) ;
 assign _4814 = ( (~ i_14_)  &  i_13_  &  i_12_  &  wire912 ) ;
 assign _4861 = ( wire118  &  n_n100 ) | ( wire132  &  n_n100 ) | ( n_n100  &  _36826 ) ;
 assign _4868 = ( wire70  &  n_n100 ) | ( n_n100  &  wire184 ) | ( n_n100  &  _36821 ) ;
 assign _4878 = ( wire113  &  n_n94 ) | ( n_n94  &  wire281 ) | ( n_n94  &  _4881 ) ;
 assign _4881 = ( i_14_  &  (~ i_13_)  &  i_12_  &  wire907 ) ;
 assign _4901 = ( n_n260  &  n_n285  &  n_n263  &  wire130 ) ;
 assign _4906 = ( wire153  &  n_n100 ) | ( wire57  &  n_n100 ) | ( n_n100  &  _4909 ) ;
 assign _4907 = ( wire166  &  n_n100 ) | ( wire180  &  n_n100 ) ;
 assign _4908 = ( wire55  &  n_n100 ) | ( n_n279  &  wire912  &  n_n100 ) ;
 assign _4909 = ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire914 ) ;
 assign _4920 = ( n_n260  &  n_n285  &  wire112  &  n_n263 ) ;
 assign _4943 = ( wire224  &  n_n100 ) | ( wire99  &  n_n100 ) | ( wire41  &  n_n100 ) ;
 assign _4944 = ( wire254  &  n_n100 ) | ( n_n100  &  wire255 ) ;
 assign _4977 = ( n_n260  &  n_n285  &  n_n263  &  wire1194 ) ;
 assign _5028 = ( wire913  &  n_n121  &  _35748 ) ;
 assign _5079 = ( i_7_  &  i_6_  &  n_n264  &  n_n120 ) ;
 assign _5101 = ( n_n5  &  wire64 ) | ( n_n5  &  wire89 ) | ( n_n5  &  _36116 ) ;
 assign _5118 = ( n_n56  &  wire66 ) | ( n_n56  &  wire79 ) | ( n_n56  &  _36518 ) ;
 assign _5119 = ( n_n56  &  wire42 ) | ( n_n279  &  n_n56  &  wire899 ) ;
 assign _5135 = ( n_n56  &  n_n259  &  _35950 ) | ( n_n56  &  n_n259  &  _35951 ) ;
 assign _5145 = ( n_n285  &  n_n271  &  n_n230  &  wire132 ) ;
 assign _5150 = ( n_n6  &  wire19407 ) | ( n_n6  &  wire19408 ) | ( n_n6  &  _36193 ) ;
 assign _5153 = ( n_n5  &  wire453 ) | ( n_n5  &  wire245 ) | ( n_n5  &  _36203 ) ;
 assign _5158 = ( n_n6  &  wire88 ) | ( n_n6  &  wire61 ) | ( n_n6  &  _36205 ) ;
 assign _5164 = ( n_n5  &  wire61 ) | ( n_n5  &  wire52 ) | ( n_n5  &  _36489 ) ;
 assign _5165 = ( n_n5  &  wire88 ) | ( n_n5  &  wire80 ) | ( n_n5  &  _36491 ) ;
 assign _5173 = ( n_n5  &  wire19738 ) | ( n_n5  &  wire84 ) | ( n_n5  &  _36476 ) ;
 assign _5174 = ( n_n5  &  wire66 ) | ( n_n5  &  wire899  &  n_n256 ) ;
 assign _5179 = ( n_n6  &  wire84 ) | ( n_n6  &  wire52 ) | ( n_n6  &  _36161 ) ;
 assign _5183 = ( n_n5  &  wire79 ) | ( n_n5  &  wire101 ) | ( n_n5  &  _36467 ) ;
 assign _5218 = ( wire48  &  n_n152 ) | ( n_n152  &  wire103 ) | ( n_n152  &  _36430 ) ;
 assign _5219 = ( n_n152  &  wire54 ) | ( n_n152  &  n_n220  &  wire914 ) ;
 assign _5225 = ( i_7_  &  (~ i_6_)  &  n_n260  &  n_n165 ) ;
 assign _5227 = ( wire54  &  n_n130 ) | ( wire103  &  n_n130 ) | ( n_n130  &  _5241 ) ;
 assign _5230 = ( wire54  &  n_n132 ) | ( wire54  &  _5239 ) | ( n_n132  &  _36421 ) | ( _5239  &  _36421 ) ;
 assign _5231 = ( wire103  &  n_n132 ) | ( wire103  &  _5239 ) | ( n_n132  &  _5355 ) | ( _5239  &  _5355 ) ;
 assign _5239 = ( n_n260  &  n_n229  &  n_n165 ) ;
 assign _5241 = ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  wire913 ) ;
 assign _5244 = ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  wire905 ) ;
 assign _5274 = ( n_n56  &  wire84 ) | ( n_n56  &  wire52 ) | ( n_n56  &  _36396 ) ;
 assign _5282 = ( n_n268  &  wire50 ) | ( n_n268  &  wire157 ) | ( n_n268  &  _5288 ) ;
 assign _5283 = ( n_n268  &  wire130 ) | ( wire911  &  n_n228  &  n_n268 ) ;
 assign _5288 = ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  wire903 ) ;
 assign _5302 = ( n_n268  &  wire55 ) | ( n_n268  &  wire57 ) | ( n_n268  &  _36383 ) ;
 assign _5303 = ( n_n284  &  n_n285  &  n_n271  &  wire273 ) ;
 assign _5309 = ( n_n268  &  wire210 ) | ( n_n268  &  wire190 ) | ( n_n268  &  wire119 ) ;
 assign _5310 = ( n_n268  &  wire60 ) | ( n_n268  &  wire52 ) | ( n_n268  &  _36377 ) ;
 assign _5341 = ( n_n121  &  wire419 ) | ( n_n121  &  wire19604 ) | ( n_n121  &  _36331 ) ;
 assign _5346 = ( wire54  &  n_n127 ) | ( n_n127  &  _36317 ) ;
 assign _5347 = ( wire103  &  n_n127 ) | ( n_n220  &  wire914  &  n_n127 ) ;
 assign _5355 = ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  wire914 ) ;
 assign _5357 = ( wire54  &  n_n124 ) | ( wire103  &  n_n124 ) | ( n_n124  &  _35745 ) ;
 assign _5359 = ( wire54  &  n_n122 ) | ( wire103  &  n_n122 ) | ( n_n122  &  _5362 ) ;
 assign _5362 = ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  wire913 ) ;
 assign _5365 = ( wire75  &  n_n1 ) | ( n_n1  &  wire72 ) | ( n_n1  &  _36308 ) ;
 assign _5376 = ( n_n2  &  wire118 ) | ( n_n2  &  wire63 ) | ( n_n2  &  _36304 ) ;
 assign _5377 = ( wire75  &  n_n2 ) | ( n_n2  &  wire72 ) | ( n_n2  &  _5378 ) ;
 assign _5378 = ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  wire913 ) ;
 assign _5381 = ( n_n260  &  n_n285  &  n_n283  &  wire1627 ) ;
 assign _5389 = ( n_n1  &  wire96 ) | ( n_n1  &  wire807 ) | ( n_n1  &  _35428 ) ;
 assign _5392 = ( n_n2  &  wire96 ) | ( n_n2  &  wire807 ) | ( n_n2  &  _35352 ) ;
 assign _5399 = ( n_n2  &  wire89 ) | ( n_n2  &  wire71 ) | ( n_n2  &  _36291 ) ;
 assign _5405 = ( n_n2  &  _36285 ) | ( n_n2  &  _36286 ) ;
 assign _5408 = ( n_n1  &  wire19385 ) | ( n_n1  &  wire19384 ) | ( n_n1  &  _35377 ) ;
 assign _5422 = ( n_n1  &  wire73 ) | ( n_n1  &  wire63 ) | ( n_n1  &  _36275 ) ;
 assign _5425 = ( n_n2  &  wire84 ) | ( n_n2  &  wire52 ) | ( n_n2  &  _36270 ) ;
 assign _5426 = ( n_n2  &  wire19738 ) | ( wire913  &  n_n2  &  n_n256 ) ;
 assign _5435 = ( n_n1  &  wire66 ) | ( n_n1  &  wire79 ) | ( n_n1  &  _36265 ) ;
 assign _5446 = ( n_n2  &  wire66 ) | ( n_n2  &  wire42 ) | ( n_n2  &  _36256 ) ;
 assign _5457 = ( n_n2  &  wire57 ) | ( n_n2  &  wire86 ) | ( n_n2  &  _36245 ) ;
 assign _5458 = ( n_n2  &  wire64 ) | ( n_n2  &  wire55 ) | ( n_n2  &  _5459 ) ;
 assign _5459 = ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire907 ) ;
 assign _5462 = ( n_n1  &  wire64 ) | ( n_n1  &  wire86 ) | ( n_n1  &  _36242 ) ;
 assign _5470 = ( n_n2  &  wire80 ) | ( n_n2  &  wire61 ) | ( n_n2  &  _35370 ) ;
 assign _5480 = ( n_n5  &  wire453 ) | ( n_n5  &  wire245 ) | ( n_n5  &  _36203 ) ;
 assign _5481 = ( n_n6  &  wire88 ) | ( n_n6  &  wire61 ) | ( n_n6  &  _36205 ) ;
 assign _5485 = ( n_n5  &  wire57 ) | ( n_n5  &  wire86 ) | ( n_n5  &  _36224 ) ;
 assign _5501 = ( n_n6  &  wire19407 ) | ( n_n6  &  wire19408 ) | ( n_n6  &  _36193 ) ;
 assign _5502 = ( n_n6  &  wire42 ) | ( n_n6  &  wire53 ) | ( n_n6  &  _36195 ) ;
 assign _5503 = ( n_n5  &  wire88 ) | ( n_n5  &  wire80 ) | ( n_n5  &  _36190 ) ;
 assign _5552 = ( n_n6  &  wire84 ) | ( n_n6  &  wire52 ) | ( n_n6  &  _36161 ) ;
 assign _5559 = ( n_n5  &  wire19738 ) | ( n_n5  &  wire84 ) | ( n_n5  &  _36157 ) ;
 assign _5578 = ( n_n5  &  wire73 ) | ( n_n5  &  wire79 ) | ( n_n5  &  _36140 ) ;
 assign _5593 = ( n_n5  &  wire64 ) | ( n_n5  &  wire89 ) | ( n_n5  &  _36116 ) ;
 assign _5604 = ( n_n6  &  wire245 ) | ( n_n6  &  wire57 ) | ( n_n6  &  _36096 ) ;
 assign _5617 = ( n_n5  &  wire68 ) | ( n_n5  &  wire96 ) | ( n_n5  &  _5620 ) ;
 assign _5618 = ( n_n5  &  _36085 ) | ( n_n5  &  _36086 ) ;
 assign _5619 = ( n_n5  &  wire19385 ) | ( n_n5  &  n_n256  &  wire900 ) ;
 assign _5620 = ( i_14_  &  i_13_  &  (~ i_12_)  &  wire904 ) ;
 assign _5624 = ( n_n6  &  wire19385 ) | ( n_n6  &  n_n256  &  wire900 ) ;
 assign _5751 = ( n_n56  &  wire52 ) | ( n_n56  &  wire167 ) | ( n_n56  &  _5753 ) ;
 assign _5752 = ( n_n56  &  wire60 ) | ( n_n56  &  wire140 ) | ( n_n56  &  _5756 ) ;
 assign _5753 = ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire913 ) ;
 assign _5756 = ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire911 ) ;
 assign _5776 = ( n_n57  &  wire60 ) | ( n_n57  &  wire52 ) | ( n_n57  &  _35941 ) ;
 assign _5783 = ( n_n56  &  wire123 ) | ( n_n56  &  wire247 ) | ( n_n56  &  wire227 ) ;
 assign _5807 = ( n_n56  &  wire113 ) | ( n_n56  &  wire281 ) | ( n_n56  &  _5810 ) ;
 assign _5810 = ( i_14_  &  (~ i_13_)  &  i_12_  &  wire907 ) ;
 assign _5820 = ( n_n57  &  wire70 ) | ( n_n57  &  wire184 ) | ( n_n57  &  _5823 ) ;
 assign _5823 = ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  wire898 ) ;
 assign _5889 = ( n_n127  &  wire250 ) | ( n_n127  &  wire19604 ) | ( n_n127  &  _35763 ) ;
 assign _5900 = ( wire54  &  n_n124 ) | ( wire103  &  n_n124 ) | ( n_n124  &  _35745 ) ;
 assign _5901 = ( wire48  &  n_n124 ) | ( n_n124  &  _35749 ) ;
 assign _5905 = ( n_n165  &  n_n208  &  n_n284  &  wire939 ) ;
 assign _5910 = ( i_7_  &  i_6_  &  n_n264  &  n_n118 ) | ( (~ i_7_)  &  i_6_  &  n_n264  &  n_n118 ) | ( i_7_  &  (~ i_6_)  &  n_n264  &  n_n118 ) ;
 assign _5922 = ( wire71  &  n_n100 ) | ( n_n100  &  wire19575 ) | ( n_n100  &  _35712 ) ;
 assign _5925 = ( n_n100  &  wire19578 ) | ( n_n100  &  wire59 ) | ( n_n100  &  _35706 ) ;
 assign _5932 = ( n_n94  &  wire96 ) | ( n_n94  &  wire19575 ) | ( n_n94  &  _35700 ) ;
 assign _5940 = ( wire51  &  n_n94 ) | ( wire71  &  n_n94 ) | ( n_n94  &  _5943 ) ;
 assign _5943 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire898 ) ;
 assign _5967 = ( wire902  &  n_n258  &  n_n100 ) ;
 assign _5968 = ( wire88  &  n_n100 ) | ( n_n100  &  wire65 ) | ( n_n100  &  _35652 ) ;
 assign _5980 = ( n_n100  &  wire104 ) | ( n_n100  &  wire74 ) | ( n_n100  &  _35635 ) ;
 assign _5981 = ( wire44  &  n_n100 ) | ( n_n258  &  wire904  &  n_n100 ) ;
 assign _5982 = ( n_n100  &  wire19457 ) | ( n_n222  &  n_n100  &  wire897 ) ;
 assign _5993 = ( n_n94  &  wire69 ) | ( n_n94  &  wire65 ) | ( n_n94  &  _5996 ) ;
 assign _5996 = ( (~ i_14_)  &  i_13_  &  i_12_  &  wire902 ) ;
 assign _6010 = ( n_n56  &  wire76 ) | ( n_n56  &  wire19385 ) | ( n_n56  &  _35603 ) ;
 assign _6034 = ( wire44  &  n_n94 ) | ( wire63  &  n_n94 ) | ( n_n94  &  _35592 ) ;
 assign _6055 = ( n_n56  &  wire19407 ) | ( n_n56  &  wire53 ) | ( n_n56  &  _35577 ) ;
 assign _6058 = ( n_n57  &  wire19385 ) | ( n_n57  &  wire19384 ) | ( n_n57  &  _35572 ) ;
 assign _6069 = ( n_n57  &  wire19407 ) | ( n_n57  &  _35567 ) ;
 assign _6070 = ( n_n57  &  wire53 ) | ( n_n279  &  n_n57  &  wire897 ) ;
 assign _6077 = ( n_n57  &  wire80 ) | ( n_n57  &  wire61 ) | ( n_n57  &  _35563 ) ;
 assign _6157 = ( n_n4  &  wire70 ) | ( n_n4  &  wire19408 ) | ( n_n4  &  _35502 ) ;
 assign _6160 = ( n_n3  &  _35498 ) | ( n_n3  &  _35499 ) ;
 assign _6161 = ( n_n3  &  wire88 ) | ( n_n3  &  wire80 ) | ( n_n3  &  _35500 ) ;
 assign _6176 = ( n_n3  &  wire53 ) | ( n_n3  &  wire19408 ) | ( n_n3  &  _35485 ) ;
 assign _6177 = ( n_n3  &  wire19407 ) | ( n_n3  &  _35487 ) ;
 assign _6189 = ( n_n3  &  wire50 ) | ( n_n3  &  wire19402 ) | ( n_n3  &  _6192 ) ;
 assign _6192 = ( i_14_  &  i_13_  &  i_12_  &  wire897 ) ;
 assign _6205 = ( n_n2  &  wire50 ) | ( n_n2  &  wire19394 ) | ( n_n2  &  _6208 ) ;
 assign _6208 = ( i_14_  &  i_13_  &  i_12_  &  wire897 ) ;
 assign _6220 = ( n_n3  &  wire96 ) | ( n_n3  &  wire807 ) | ( n_n3  &  _35454 ) ;
 assign _6221 = ( n_n4  &  wire76 ) | ( n_n4  &  wire19385 ) | ( n_n4  &  _35456 ) ;
 assign _6235 = ( n_n4  &  wire96 ) | ( n_n4  &  wire807 ) | ( n_n4  &  _35446 ) ;
 assign _6236 = ( n_n208  &  n_n284  &  n_n285  &  wire68 ) ;
 assign _6237 = ( n_n3  &  wire19384 ) | ( n_n3  &  _35444 ) ;
 assign _6238 = ( n_n3  &  wire19385 ) | ( n_n3  &  n_n256  &  wire900 ) ;
 assign _6252 = ( n_n1  &  wire96 ) | ( n_n1  &  wire807 ) | ( n_n1  &  _35428 ) ;
 assign _6280 = ( n_n2  &  _35381 ) | ( n_n2  &  _35382 ) ;
 assign _6287 = ( n_n1  &  wire19385 ) | ( n_n1  &  wire19384 ) | ( n_n1  &  _35377 ) ;
 assign _6294 = ( n_n2  &  wire80 ) | ( n_n2  &  wire61 ) | ( n_n2  &  _35370 ) ;
 assign _6298 = ( n_n2  &  wire19407 ) | ( n_n2  &  wire53 ) | ( n_n2  &  _35366 ) ;
 assign _6301 = ( n_n2  &  wire903  &  _35101 ) ;
 assign _6319 = ( n_n2  &  wire96 ) | ( n_n2  &  wire807 ) | ( n_n2  &  _35352 ) ;
 assign _6363 = ( n_n5  &  wire124 ) | ( n_n5  &  wire212 ) | ( n_n5  &  wire119 ) ;
 assign _6387 = ( n_n285  &  n_n230  &  n_n263  &  wire166 ) ;
 assign _6408 = ( wire88  &  n_n53 ) | ( n_n53  &  wire61 ) | ( n_n53  &  _35213 ) ;
 assign _6443 = ( n_n48  &  wire96 ) | ( n_n48  &  wire807 ) | ( n_n48  &  _35178 ) ;
 assign _6447 = ( n_n48  &  wire19385 ) | ( n_n48  &  wire19384 ) | ( n_n48  &  _35172 ) ;
 assign _6448 = ( n_n48  &  wire76 ) | ( n_n48  &  _35174 ) ;
 assign _6461 = ( n_n53  &  wire96 ) | ( n_n53  &  wire807 ) | ( n_n53  &  _35148 ) ;
 assign _6474 = ( n_n53  &  wire19407 ) | ( n_n53  &  wire19408 ) | ( n_n53  &  _35125 ) ;
 assign _6483 = ( n_n48  &  wire53 ) | ( n_n48  &  wire19408 ) | ( n_n48  &  _35112 ) ;
 assign _6484 = ( n_n48  &  wire19407 ) | ( n_n48  &  _35116 ) ;
 assign _6540 = ( wire63  &  n_n48 ) | ( n_n48  &  wire50 ) | ( n_n48  &  _35040 ) ;
 assign _6592 = ( (~ i_9_)  &  (~ i_10_) ) ;
 assign _6597 = ( n_n139  &  wire54 ) | ( n_n139  &  wire103 ) | ( n_n139  &  _34957 ) ;
 assign _6700 = ( n_n152  &  wire326 ) | ( n_n152  &  wire19244 ) | ( n_n152  &  _6703 ) ;
 assign _6703 = ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  wire911 ) ;
 assign _6706 = ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  wire914 ) ;
 assign _6708 = ( n_n284  &  _6730  &  _34827 ) | ( n_n284  &  _34827  &  _34834 ) ;
 assign _6730 = ( n_n283  &  n_n282  &  wire152 ) | ( n_n283  &  n_n282  &  _34642 ) ;
 assign _6812 = ( n_n152  &  wire19239 ) | ( n_n152  &  wire214 ) | ( n_n152  &  _34720 ) ;
 assign _6813 = ( n_n152  &  wire19237 ) | ( n_n152  &  _34722 ) ;
 assign _6821 = ( n_n136  &  wire321 ) | ( n_n136  &  _34715 ) ;
 assign _6822 = ( n_n136  &  wire331 ) | ( n_n136  &  wire19233 ) | ( n_n136  &  _6827 ) ;
 assign _6824 = ( (~ i_9_)  &  (~ i_10_) ) ;
 assign _6827 = ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  wire911 ) ;
 assign _6830 = ( n_n139  &  wire19239 ) | ( n_n139  &  wire19238 ) | ( n_n139  &  _34708 ) ;
 assign _6836 = ( n_n142  &  wire321 ) | ( n_n142  &  _34703 ) ;
 assign _6837 = ( n_n142  &  wire331 ) | ( n_n142  &  wire19233 ) | ( n_n142  &  _6843 ) ;
 assign _6838 = ( (~ i_9_)  &  (~ i_10_) ) ;
 assign _6843 = ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  wire911 ) ;
 assign _6848 = ( wire896  &  _6857 ) | ( wire896  &  _6858 ) | ( wire896  &  _6859 ) ;
 assign _6849 = ( n_n273  &  n_n230  &  _34695 ) ;
 assign _6857 = ( wire196  &  _34696 ) | ( n_n247  &  wire152  &  _34696 ) ;
 assign _6858 = ( _34697  &  _34698 ) | ( n_n281  &  wire912  &  _34698 ) ;
 assign _6859 = ( i_7_  &  (~ i_8_)  &  (~ i_6_) ) ;
 assign _6865 = ( n_n132  &  wire19244 ) | ( n_n132  &  wire19255 ) | ( n_n132  &  _6868 ) ;
 assign _6866 = ( n_n132  &  wire19253 ) | ( n_n279  &  n_n132  &  wire912 ) ;
 assign _6868 = ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  wire911 ) ;
 assign _6927 = ( n_n128  &  wire397 ) | ( n_n128  &  wire19307 ) | ( n_n128  &  _6930 ) ;
 assign _6928 = ( n_n128  &  wire130 ) | ( wire911  &  n_n279  &  n_n128 ) ;
 assign _6930 = ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  wire914 ) ;
 assign _6970 = ( n_n127  &  wire184 ) | ( n_n127  &  wire130 ) | ( n_n127  &  _34583 ) ;
 assign _6977 = ( n_n124  &  wire19238 ) | ( n_n124  &  wire19237 ) | ( n_n124  &  _34567 ) ;
 assign _6984 = ( n_n122  &  wire19253 ) | ( n_n122  &  wire19311 ) | ( n_n122  &  _34551 ) ;
 assign _6995 = ( n_n121  &  wire397 ) | ( n_n121  &  wire19307 ) | ( n_n121  &  _6998 ) ;
 assign _6996 = ( n_n121  &  wire19237 ) | ( n_n121  &  _34535 ) ;
 assign _6997 = ( n_n121  &  wire130 ) | ( wire911  &  n_n279  &  n_n121 ) ;
 assign _6998 = ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  wire914 ) ;
 assign _34535 = ( wire328 ) | ( n_n220  &  wire912 ) ;
 assign _34536 = ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  i_15_ ) ;
 assign _34537 = ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  (~ i_15_) ) ;
 assign _34544 = ( i_14_  &  (~ i_13_)  &  (~ i_12_) ) ;
 assign _34546 = ( (~ i_14_)  &  i_13_  &  (~ i_12_) ) ;
 assign _34548 = ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  i_15_ ) ;
 assign _34549 = ( i_14_  &  i_13_  &  (~ i_12_) ) ;
 assign _34551 = ( wire912  &  _34544 ) | ( wire911  &  _34546 ) ;
 assign _34558 = ( (~ i_9_)  &  i_10_  &  i_11_ ) | ( i_9_  &  (~ i_10_)  &  i_11_ ) | ( (~ i_9_)  &  i_10_  &  i_12_  &  (~ i_11_) ) | ( i_9_  &  (~ i_10_)  &  i_12_  &  (~ i_11_) ) ;
 assign _34559 = ( wire5874 ) | ( _6984 ) | ( n_n122  &  wire19313 ) ;
 assign _34563 = ( (~ i_14_)  &  i_13_  &  (~ i_12_) ) ;
 assign _34565 = ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_) ) ;
 assign _34567 = ( wire912  &  _34563 ) | ( wire914  &  _34565 ) ;
 assign _34575 = ( i_14_  &  (~ i_13_)  &  (~ i_12_) ) ;
 assign _34576 = ( n_n124  &  wire19239 ) | ( n_n124  &  wire899  &  _34575 ) ;
 assign _34580 = ( i_14_  &  (~ i_13_)  &  (~ i_12_) ) ;
 assign _34581 = ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  i_15_ ) ;
 assign _34582 = ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  (~ i_15_) ) ;
 assign _34583 = ( wire196 ) | ( wire911  &  _34580 ) ;
 assign _34585 = ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  i_15_ ) ;
 assign _34586 = ( n_n127  &  wire397 ) | ( n_n127  &  wire19334 ) ;
 assign _34594 = ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  i_15_ ) ;
 assign _34606 = ( _6970 ) | ( _6977 ) | ( _34576 ) | ( _34586 ) ;
 assign _34625 = ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  i_15_ ) ;
 assign _34626 = ( i_14_  &  i_13_  &  (~ i_12_) ) ;
 assign _34627 = ( wire911  &  _34546 ) | ( wire899  &  _34575 ) ;
 assign _34637 = ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  i_15_ ) ;
 assign _34638 = ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  i_15_ ) ;
 assign _34639 = ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  (~ i_15_) ) ;
 assign _34642 = ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  i_15_ ) ;
 assign _34644 = ( n_n165  &  n_n273  &  n_n284 ) ;
 assign _34645 = ( wire5850 ) | ( wire384  &  _34644 ) ;
 assign _34685 = ( wire5875 ) | ( n_n5009 ) | ( wire19355 ) | ( _34559 ) ;
 assign _34687 = ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  wire905 ) ;
 assign _34692 = ( i_9_  &  i_10_  &  i_11_ ) | ( i_9_  &  (~ i_10_)  &  i_11_ ) | ( i_9_  &  i_10_  &  i_12_  &  (~ i_11_) ) | ( i_9_  &  (~ i_10_)  &  i_12_  &  (~ i_11_) ) ;
 assign _34695 = ( i_1_  &  (~ i_2_)  &  (~ i_0_) ) ;
 assign _34696 = ( i_7_  &  i_8_  &  (~ i_6_) ) ;
 assign _34697 = ( (~ i_9_) ) | ( i_9_  &  i_10_ ) ;
 assign _34698 = ( i_7_  &  i_8_  &  (~ i_6_) ) ;
 assign _34702 = ( (~ i_12_)  &  i_13_ ) ;
 assign _34703 = ( wire215 ) | ( _6838 ) | ( n_n242  &  _34702 ) ;
 assign _34708 = ( wire914  &  _34565 ) | ( wire899  &  _34575 ) ;
 assign _34710 = ( n_n253 ) | ( n_n220  &  wire912 ) ;
 assign _34711 = ( n_n139  &  wire435 ) | ( n_n139  &  wire19237 ) | ( n_n139  &  _34710 ) ;
 assign _34713 = ( n_n165  &  n_n283  &  n_n230 ) ;
 assign _34715 = ( wire215 ) | ( _6824 ) | ( n_n242  &  _34702 ) ;
 assign _34720 = ( n_n143 ) | ( wire899  &  _34575 ) ;
 assign _34722 = ( n_n253 ) | ( n_n220  &  wire912 ) ;
 assign _34724 = ( _6830 ) | ( _6836 ) | ( _6837 ) | ( _34711 ) ;
 assign _34730 = ( i_14_  &  (~ i_13_)  &  i_12_  &  (~ i_15_) ) ;
 assign _34738 = ( (~ i_9_)  &  i_10_  &  (~ i_11_) ) ;
 assign _34748 = ( i_9_  &  (~ i_10_)  &  i_11_ ) ;
 assign _34780 = ( i_9_  &  i_10_  &  (~ i_11_) ) ;
 assign _34797 = ( i_5_  &  i_6_  &  (~ i_3_)  &  (~ i_4_) ) ;
 assign _34819 = ( (~ i_9_)  &  i_5_  &  (~ i_3_)  &  (~ i_4_) ) ;
 assign _34822 = ( i_9_  &  i_5_  &  (~ i_3_)  &  (~ i_4_) ) ;
 assign _34827 = ( (~ i_1_)  &  (~ i_2_)  &  (~ i_0_) ) ;
 assign _34834 = ( i_7_  &  (~ i_6_) ) | ( (~ i_7_)  &  i_8_  &  (~ i_6_) ) | ( (~ i_7_)  &  (~ i_8_)  &  (~ i_6_)  &  wire19205 ) ;
 assign _34842 = ( wire5988 ) | ( n_n152  &  wire19238 ) | ( n_n152  &  _6706 ) ;
 assign _34843 = ( i_9_  &  (~ i_7_)  &  i_8_  &  (~ i_6_) ) ;
 assign _34860 = ( i_5_  &  i_3_  &  (~ i_4_) ) ;
 assign _34908 = ( i_9_  &  (~ i_10_)  &  i_11_ ) ;
 assign _34910 = ( i_9_  &  (~ i_10_)  &  (~ i_11_) ) ;
 assign _34914 = ( i_9_  &  i_10_  &  (~ i_11_) ) ;
 assign _34919 = ( (~ i_9_)  &  (~ i_10_)  &  i_11_ ) ;
 assign _34942 = ( wire19359 ) | ( wire19260 ) | ( wire19261 ) | ( wire19263 ) ;
 assign _34949 = ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  i_15_ ) ;
 assign _34950 = ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  (~ i_15_) ) ;
 assign _34952 = ( (~ i_14_)  &  i_13_  &  (~ i_12_) ) ;
 assign _34953 = ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  i_15_ ) ;
 assign _34954 = ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  (~ i_15_) ) ;
 assign _34956 = ( (~ i_14_)  &  i_13_  &  (~ i_12_) ) ;
 assign _34957 = ( wire914  &  _34952 ) | ( wire905  &  _34956 ) ;
 assign _34985 = ( i_5_  &  (~ i_3_)  &  i_4_ ) ;
 assign _34990 = ( (~ i_5_)  &  (~ i_3_)  &  i_4_ ) ;
 assign _35004 = ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_) ) ;
 assign _35011 = ( wire19373 ) | ( wire19374 ) | ( wire19365 ) | ( _6597 ) ;
 assign _35013 = ( i_14_  &  (~ i_13_)  &  i_12_  &  wire898 ) ;
 assign _35014 = ( i_14_  &  i_13_  &  (~ i_12_)  &  wire898 ) ;
 assign _35030 = ( n_n6  &  wire99 ) | ( n_n6  &  _35013 ) | ( n_n6  &  _35014 ) ;
 assign _35033 = ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_) ) ;
 assign _35034 = ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  i_15_ ) ;
 assign _35035 = ( i_14_  &  (~ i_13_)  &  i_12_  &  (~ i_15_) ) ;
 assign _35036 = ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  i_15_ ) ;
 assign _35037 = ( i_14_  &  (~ i_13_)  &  i_12_  &  (~ i_15_) ) ;
 assign _35039 = ( i_14_  &  i_13_  &  i_12_ ) ;
 assign _35040 = ( wire908  &  _35033 ) | ( wire897  &  _35039 ) ;
 assign _35042 = ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  i_15_ ) ;
 assign _35043 = ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  (~ i_15_) ) ;
 assign _35044 = ( wire44  &  n_n48 ) | ( n_n48  &  wire19491 ) ;
 assign _35046 = ( i_14_  &  (~ i_13_)  &  i_12_ ) ;
 assign _35049 = ( (~ i_14_)  &  i_13_  &  (~ i_12_) ) ;
 assign _35051 = ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  i_15_ ) ;
 assign _35052 = ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  (~ i_15_) ) ;
 assign _35053 = ( i_14_  &  (~ i_13_)  &  i_12_  &  (~ i_15_) ) ;
 assign _35054 = ( i_14_  &  i_13_  &  i_12_  &  i_15_ ) ;
 assign _35056 = ( i_14_  &  i_13_  &  i_12_ ) ;
 assign _35058 = ( wire5613 ) | ( _6540 ) | ( _35030 ) | ( _35044 ) ;
 assign _35064 = ( i_14_  &  i_13_  &  i_12_  &  (~ i_15_) ) ;
 assign _35065 = ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  i_15_ ) ;
 assign _35071 = ( i_14_  &  i_13_  &  (~ i_12_) ) ;
 assign _35074 = ( i_14_  &  i_13_  &  i_12_ ) ;
 assign _35076 = ( (~ i_14_)  &  i_13_  &  i_12_  &  (~ i_15_) ) ;
 assign _35077 = ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  i_15_ ) ;
 assign _35079 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_ ) ;
 assign _35084 = ( i_14_  &  (~ i_13_)  &  i_12_  &  (~ i_15_) ) ;
 assign _35085 = ( i_14_  &  i_13_  &  i_12_  &  i_15_ ) ;
 assign _35086 = ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  i_15_ ) ;
 assign _35087 = ( i_14_  &  (~ i_13_)  &  i_12_  &  (~ i_15_) ) ;
 assign _35091 = ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_) ) ;
 assign _35097 = ( i_14_  &  i_13_  &  (~ i_12_) ) ;
 assign _35099 = ( i_14_  &  (~ i_13_)  &  i_12_ ) ;
 assign _35101 = ( (~ i_14_)  &  i_13_  &  (~ i_12_) ) ;
 assign _35103 = ( i_14_  &  (~ i_13_)  &  (~ i_12_) ) ;
 assign _35109 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_ ) ;
 assign _35110 = ( (~ i_14_)  &  i_13_  &  i_12_  &  (~ i_15_) ) ;
 assign _35111 = ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  i_15_ ) ;
 assign _35112 = ( wire897  &  _35103 ) | ( wire903  &  _35109 ) ;
 assign _35114 = ( (~ i_14_)  &  i_13_  &  i_12_  &  i_15_ ) ;
 assign _35115 = ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  (~ i_15_) ) ;
 assign _35116 = ( i_14_  &  (~ i_13_)  &  i_12_  &  wire897 ) | ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire897 ) | ( i_14_  &  i_13_  &  (~ i_12_)  &  wire897 ) ;
 assign _35118 = ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  wire902 ) ;
 assign _35120 = ( (~ i_14_)  &  i_13_  &  i_12_ ) ;
 assign _35124 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_ ) ;
 assign _35125 = ( wire903  &  _35109 ) | ( wire897  &  _35124 ) ;
 assign _35129 = ( n_n1542 ) | ( wire5596 ) | ( _6483 ) | ( _6484 ) ;
 assign _35131 = ( wire19495 ) | ( wire19502 ) | ( _35058 ) | ( _35129 ) ;
 assign _35137 = ( (~ i_14_)  &  i_13_  &  (~ i_12_) ) ;
 assign _35139 = ( i_14_  &  (~ i_13_)  &  (~ i_12_) ) ;
 assign _35141 = ( i_14_  &  i_13_  &  (~ i_12_) ) ;
 assign _35142 = ( i_14_  &  i_13_  &  i_12_  &  (~ i_15_) ) ;
 assign _35143 = ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  i_15_ ) ;
 assign _35148 = ( i_14_  &  i_13_  &  (~ i_12_)  &  wire904 ) | ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire904 ) ;
 assign _35150 = ( (~ i_14_)  &  i_13_  &  i_12_  &  (~ i_15_) ) ;
 assign _35151 = ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  i_15_ ) ;
 assign _35153 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_ ) ;
 assign _35154 = ( n_n53  &  wire71 ) | ( wire904  &  n_n53  &  _35153 ) ;
 assign _35160 = ( i_14_  &  (~ i_13_)  &  (~ i_12_) ) ;
 assign _35163 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_ ) ;
 assign _35164 = ( (~ i_14_)  &  i_13_  &  i_12_  &  i_15_ ) ;
 assign _35165 = ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  (~ i_15_) ) ;
 assign _35167 = ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_) ) ;
 assign _35172 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire900 ) | ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  wire900 ) ;
 assign _35174 = ( n_n220  &  wire906 ) | ( wire900  &  _35160 ) ;
 assign _35176 = ( _6447 ) | ( _6448 ) | ( _6461 ) | ( _35154 ) ;
 assign _35178 = ( i_14_  &  i_13_  &  (~ i_12_)  &  wire904 ) | ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire904 ) ;
 assign _35186 = ( (~ i_14_)  &  i_13_  &  (~ i_12_) ) ;
 assign _35190 = ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_) ) ;
 assign _35208 = ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  wire904 ) ;
 assign _35212 = ( i_14_  &  (~ i_13_)  &  (~ i_12_) ) ;
 assign _35213 = ( i_14_  &  i_13_  &  (~ i_12_)  &  wire908 ) | ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire908 ) ;
 assign _35218 = ( wire662 ) | ( wire5564 ) | ( wire5565 ) | ( _6443 ) ;
 assign _35219 = ( n_n3843 ) | ( wire5569 ) | ( _35176 ) | ( _35218 ) ;
 assign _35235 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire904 ) ;
 assign _35236 = ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  wire904 ) ;
 assign _35255 = ( n_n285  &  n_n230  &  n_n261 ) ;
 assign _35257 = ( wire674 ) | ( wire224  &  _35255 ) ;
 assign _35258 = ( wire389 ) | ( wire708 ) | ( wire19485 ) | ( _6387 ) ;
 assign _35290 = ( n_n285  &  n_n230  &  n_n261 ) ;
 assign _35306 = ( n_n5  &  wire140 ) | ( n_n5  &  wire198 ) ;
 assign _35339 = ( _6363 ) | ( _35306 ) | ( wire1552  &  _35290 ) ;
 assign _35341 = ( wire19530 ) | ( wire19523 ) | ( _35219 ) ;
 assign _35343 = ( i_14_  &  i_13_  &  i_12_  &  wire900 ) ;
 assign _35346 = ( n_n1  &  wire73 ) | ( n_n1  &  wire44 ) | ( n_n1  &  _35343 ) ;
 assign _35352 = ( i_14_  &  i_13_  &  (~ i_12_)  &  wire904 ) | ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire904 ) ;
 assign _35354 = ( wire395 ) | ( wire496 ) ;
 assign _35356 = ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  wire908 ) ;
 assign _35357 = ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  wire908 ) ;
 assign _35358 = ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  wire906 ) ;
 assign _35359 = ( n_n2  &  _35357 ) | ( n_n1  &  _35358 ) ;
 assign _35366 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire897 ) | ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire897 ) ;
 assign _35368 = ( n_n2  &  wire19408 ) | ( n_n2  &  wire903  &  _35109 ) ;
 assign _35370 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire908 ) | ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire908 ) ;
 assign _35372 = ( wire5725 ) | ( wire5726 ) | ( _6298 ) | ( _35368 ) ;
 assign _35376 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire900 ) ;
 assign _35377 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire900 ) | ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  wire900 ) ;
 assign _35379 = ( n_n1  &  wire71 ) | ( n_n1  &  wire904  &  _35153 ) ;
 assign _35381 = ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire900 ) | ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  wire900 ) ;
 assign _35382 = ( i_14_  &  i_13_  &  i_12_  &  wire906 ) | ( (~ i_14_)  &  i_13_  &  i_12_  &  wire906 ) | ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire906 ) | ( i_14_  &  i_13_  &  (~ i_12_)  &  wire906 ) ;
 assign _35384 = ( n_n3782 ) | ( n_n2  &  wire19385 ) | ( n_n2  &  _35376 ) ;
 assign _35389 = ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  wire898 ) ;
 assign _35391 = ( i_14_  &  (~ i_13_)  &  i_12_ ) ;
 assign _35392 = ( i_14_  &  i_13_  &  i_12_  &  wire900 ) ;
 assign _35394 = ( i_14_  &  (~ i_13_)  &  i_12_ ) ;
 assign _35396 = ( i_14_  &  i_13_  &  i_12_ ) ;
 assign _35400 = ( n_n229  &  n_n284  &  n_n285 ) ;
 assign _35412 = ( n_n229  &  n_n284  &  n_n285 ) ;
 assign _35414 = ( wire254  &  _35400 ) | ( wire1786  &  _35412 ) ;
 assign _35418 = ( i_14_  &  (~ i_13_)  &  (~ i_12_) ) ;
 assign _35420 = ( i_14_  &  i_13_  &  (~ i_12_) ) ;
 assign _35422 = ( i_14_  &  (~ i_13_)  &  i_12_ ) ;
 assign _35425 = ( (~ i_14_)  &  i_13_  &  (~ i_12_) ) ;
 assign _35427 = ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_) ) ;
 assign _35428 = ( i_14_  &  i_13_  &  (~ i_12_)  &  wire904 ) | ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire904 ) ;
 assign _35444 = ( n_n220  &  wire906 ) | ( wire900  &  _35167 ) ;
 assign _35446 = ( i_14_  &  i_13_  &  (~ i_12_)  &  wire904 ) | ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire904 ) ;
 assign _35454 = ( i_14_  &  i_13_  &  (~ i_12_)  &  wire904 ) | ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire904 ) ;
 assign _35456 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire900 ) | ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire900 ) ;
 assign _35464 = ( n_n1440 ) | ( wire5758 ) | ( _6220 ) | ( _6221 ) ;
 assign _35468 = ( n_n2  &  wire63 ) | ( n_n2  &  wire908  &  _35033 ) ;
 assign _35470 = ( n_n268  &  wire190 ) | ( n_n268  &  wire124 ) ;
 assign _35472 = ( wire5749 ) | ( wire5778 ) | ( _35470 ) ;
 assign _35476 = ( n_n3  &  wire63 ) | ( n_n3  &  wire908  &  _35033 ) ;
 assign _35478 = ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  wire904 ) ;
 assign _35480 = ( (~ i_14_)  &  i_13_  &  (~ i_12_) ) ;
 assign _35484 = ( n_n3727 ) | ( n_n7424 ) | ( _6189 ) | ( _35476 ) ;
 assign _35485 = ( wire897  &  _35103 ) | ( wire903  &  _35109 ) ;
 assign _35487 = ( n_n256  &  wire897 ) | ( wire903  &  _35101 ) ;
 assign _35494 = ( n_n1339 ) | ( wire5734 ) | ( _6176 ) | ( _6177 ) ;
 assign _35498 = ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  wire908 ) | ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire908 ) ;
 assign _35499 = ( (~ i_14_)  &  i_13_  &  i_12_  &  wire902 ) | ( i_14_  &  (~ i_13_)  &  i_12_  &  wire902 ) | ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire902 ) | ( i_14_  &  i_13_  &  (~ i_12_)  &  wire902 ) ;
 assign _35500 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire908 ) | ( i_14_  &  i_13_  &  (~ i_12_)  &  wire908 ) ;
 assign _35502 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire903 ) | ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  wire903 ) ;
 assign _35504 = ( wire546 ) | ( wire5780 ) | ( wire19381 ) | ( _6157 ) ;
 assign _35505 = ( wire19405 ) | ( wire19413 ) | ( _35484 ) | ( _35494 ) ;
 assign _35523 = ( i_14_  &  (~ i_13_)  &  i_12_  &  (~ i_15_) ) ;
 assign _35524 = ( i_14_  &  i_13_  &  i_12_  &  i_15_ ) ;
 assign _35527 = ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  i_15_ ) ;
 assign _35528 = ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  (~ i_15_) ) ;
 assign _35529 = ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  i_15_ ) ;
 assign _35530 = ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  (~ i_15_) ) ;
 assign _35531 = ( i_14_  &  (~ i_13_)  &  i_12_  &  (~ i_15_) ) ;
 assign _35532 = ( i_14_  &  i_13_  &  i_12_  &  i_15_ ) ;
 assign _35536 = ( i_14_  &  i_13_  &  i_12_  &  (~ i_15_) ) ;
 assign _35537 = ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  i_15_ ) ;
 assign _35539 = ( i_14_  &  i_13_  &  (~ i_12_) ) ;
 assign _35544 = ( i_14_  &  (~ i_13_)  &  i_12_ ) ;
 assign _35562 = ( n_n285  &  n_n271  &  n_n230 ) ;
 assign _35563 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire908 ) | ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire908 ) ;
 assign _35565 = ( n_n57  &  n_n76 ) | ( wire56  &  _35562 ) ;
 assign _35566 = ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  wire903 ) ;
 assign _35567 = ( i_14_  &  (~ i_13_)  &  i_12_  &  wire897 ) | ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire897 ) | ( i_14_  &  i_13_  &  (~ i_12_)  &  wire897 ) ;
 assign _35572 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire900 ) | ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  wire900 ) ;
 assign _35577 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire897 ) | ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire897 ) ;
 assign _35579 = ( n_n56  &  wire19408 ) | ( n_n56  &  wire903  &  _35109 ) ;
 assign _35588 = ( wire460 ) | ( wire19539 ) | ( _6055 ) | ( _35579 ) ;
 assign _35592 = ( wire902  &  _35056 ) | ( wire904  &  _35391 ) ;
 assign _35600 = ( wire5514 ) | ( wire5515 ) | ( wire5509 ) | ( wire19559 ) ;
 assign _35601 = ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  wire900 ) ;
 assign _35603 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire900 ) | ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire900 ) ;
 assign _35613 = ( n_n4685 ) | ( n_n56  &  wire19384 ) | ( n_n56  &  _35601 ) ;
 assign _35622 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_ ) ;
 assign _35623 = ( wire80  &  n_n94 ) | ( wire902  &  n_n94  &  _35622 ) ;
 assign _35626 = ( i_14_  &  (~ i_13_)  &  (~ i_12_) ) ;
 assign _35628 = ( (~ i_14_)  &  i_13_  &  i_12_ ) ;
 assign _35629 = ( (~ i_14_)  &  i_13_  &  i_12_  &  i_15_ ) ;
 assign _35630 = ( i_14_  &  i_13_  &  (~ i_12_)  &  (~ i_15_) ) ;
 assign _35635 = ( (~ i_14_)  &  i_13_  &  i_12_  &  wire903 ) | ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire903 ) ;
 assign _35639 = ( wire459 ) | ( wire19568 ) | ( _5993 ) | ( _35623 ) ;
 assign _35640 = ( wire5510 ) | ( wire19571 ) | ( _35600 ) | ( _35639 ) ;
 assign _35644 = ( i_14_  &  (~ i_13_)  &  i_12_ ) ;
 assign _35646 = ( i_14_  &  (~ i_13_)  &  i_12_ ) ;
 assign _35648 = ( wire386 ) | ( wire372 ) ;
 assign _35651 = ( (~ i_14_)  &  i_13_  &  i_12_ ) ;
 assign _35652 = ( (~ i_14_)  &  i_13_  &  i_12_  &  wire902 ) | ( i_14_  &  i_13_  &  (~ i_12_)  &  wire902 ) ;
 assign _35661 = ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_) ) ;
 assign _35685 = ( (~ i_14_)  &  i_13_  &  i_12_ ) ;
 assign _35686 = ( n_n94  &  wire59 ) | ( wire906  &  n_n94  &  _35685 ) ;
 assign _35693 = ( i_14_  &  i_13_  &  (~ i_12_) ) ;
 assign _35695 = ( (~ i_14_)  &  i_13_  &  i_12_ ) ;
 assign _35700 = ( (~ i_14_)  &  i_13_  &  i_12_  &  wire898 ) | ( i_14_  &  i_13_  &  (~ i_12_)  &  wire898 ) ;
 assign _35702 = ( (~ i_14_)  &  i_13_  &  i_12_  &  i_15_ ) ;
 assign _35703 = ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  (~ i_15_) ) ;
 assign _35705 = ( i_14_  &  i_13_  &  (~ i_12_) ) ;
 assign _35706 = ( (~ i_14_)  &  i_13_  &  i_12_  &  wire906 ) | ( i_14_  &  i_13_  &  (~ i_12_)  &  wire906 ) ;
 assign _35709 = ( n_n3884 ) | ( _5932 ) | ( _5940 ) | ( _35686 ) ;
 assign _35711 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_ ) ;
 assign _35712 = ( (~ i_14_)  &  i_13_  &  i_12_  &  wire898 ) | ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire898 ) ;
 assign _35714 = ( n_n100  &  wire96 ) | ( wire898  &  n_n100  &  _35693 ) ;
 assign _35716 = ( i_14_  &  i_13_  &  i_12_ ) ;
 assign _35719 = ( n_n260  &  n_n285  &  n_n261 ) ;
 assign _35721 = ( wire776 ) | ( wire77  &  _35719 ) ;
 assign _35722 = ( wire5472 ) | ( _5922 ) | ( _35714 ) ;
 assign _35724 = ( wire19582 ) | ( _35709 ) | ( _35721 ) | ( _35722 ) ;
 assign _35745 = ( wire914  &  _34952 ) | ( wire905  &  _34956 ) ;
 assign _35748 = ( (~ i_14_)  &  i_13_  &  (~ i_12_) ) ;
 assign _35749 = ( (~ i_9_)  &  (~ i_10_) ) | ( wire913  &  _35748 ) ;
 assign _35750 = ( wire19601 ) | ( _5900 ) | ( _5901 ) ;
 assign _35752 = ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_) ) ;
 assign _35754 = ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_) ) ;
 assign _35763 = ( wire899  &  _35752 ) | ( wire912  &  _35754 ) ;
 assign _35769 = ( n_n127  &  wire419 ) | ( n_n127  &  wire19605 ) ;
 assign _35772 = ( i_7_  &  i_6_  &  n_n165  &  n_n284 ) | ( i_7_  &  (~ i_6_)  &  n_n165  &  n_n284 ) ;
 assign _35773 = ( wire54  &  n_n124 ) | ( wire913  &  n_n124  &  _35748 ) ;
 assign _35815 = ( wire19609 ) | ( _5889 ) | ( _35769 ) | ( _35773 ) ;
 assign _35820 = ( i_7_  &  i_6_  &  i_4_ ) ;
 assign _35831 = ( (~ i_7_)  &  i_6_  &  i_4_ ) ;
 assign _35833 = ( i_7_  &  (~ i_6_)  &  i_4_ ) ;
 assign _35835 = ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  wire914 ) ;
 assign _35836 = ( n_n165  &  wire19290  &  _35831 ) | ( n_n165  &  wire19290  &  _35833 ) ;
 assign _35837 = ( _35836 ) | ( n_n152  &  wire54 ) | ( n_n152  &  _35835 ) ;
 assign _35855 = ( n_n165  &  wire19290  &  _35831 ) | ( n_n165  &  wire19290  &  _35833 ) ;
 assign _35873 = ( i_6_  &  (~ i_7_) ) ;
 assign _35875 = ( n_n5792 ) | ( n_n165  &  wire19294  &  _35873 ) ;
 assign _35876 = ( (~ i_6_)  &  i_7_ ) ;
 assign _35878 = ( n_n5794 ) | ( n_n165  &  wire19294  &  _35876 ) ;
 assign _35880 = ( i_14_  &  (~ i_13_)  &  i_12_  &  (~ i_15_) ) ;
 assign _35881 = ( i_14_  &  i_13_  &  i_12_  &  i_15_ ) ;
 assign _35882 = ( n_n57  &  wire160 ) | ( n_n57  &  wire904  &  _35427 ) ;
 assign _35883 = ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  i_15_ ) ;
 assign _35884 = ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  (~ i_15_) ) ;
 assign _35893 = ( n_n56  &  wire246 ) | ( n_n56  &  wire19683 ) ;
 assign _35897 = ( _5807 ) | ( _5820 ) | ( _35882 ) | ( _35893 ) ;
 assign _35934 = ( n_n56  &  wire100 ) | ( n_n56  &  wire210 ) ;
 assign _35938 = ( i_14_  &  (~ i_13_)  &  (~ i_12_) ) ;
 assign _35941 = ( wire911  &  _34580 ) | ( wire913  &  _35938 ) ;
 assign _35943 = ( n_n57  &  wire247 ) | ( n_n57  &  wire210 ) ;
 assign _35946 = ( (~ i_14_)  &  i_13_  &  (~ i_12_) ) ;
 assign _35947 = ( i_14_  &  (~ i_13_)  &  i_12_  &  (~ i_15_) ) ;
 assign _35948 = ( i_14_  &  i_13_  &  i_12_  &  i_15_ ) ;
 assign _35949 = ( n_n281  &  wire907 ) | ( wire901  &  _35946 ) ;
 assign _35950 = ( i_14_  &  (~ i_13_)  &  i_12_  &  (~ i_15_) ) ;
 assign _35951 = ( i_14_  &  i_13_  &  i_12_  &  i_15_ ) ;
 assign _35953 = ( (~ i_14_)  &  i_13_  &  (~ i_12_) ) ;
 assign _35954 = ( wire118  &  n_n57 ) | ( n_n57  &  wire899  &  _35953 ) ;
 assign _35956 = ( n_n285  &  n_n266  &  n_n230 ) ;
 assign _35959 = ( wire5327 ) | ( n_n3850 ) ;
 assign _35961 = ( _5776 ) | ( _5783 ) | ( _35934 ) | ( _35943 ) ;
 assign _35962 = ( wire5343 ) | ( wire5344 ) | ( _35897 ) | ( _35961 ) ;
 assign _35964 = ( n_n285  &  n_n271  &  n_n230 ) ;
 assign _35996 = ( wire481 ) | ( wire5299 ) | ( wire165  &  _35964 ) ;
 assign _35998 = ( i_14_  &  i_13_  &  i_12_  &  (~ i_15_) ) ;
 assign _35999 = ( i_14_  &  i_13_  &  (~ i_12_)  &  (~ i_15_) ) ;
 assign _36001 = ( i_14_  &  (~ i_13_)  &  i_12_  &  i_15_ ) ;
 assign _36002 = ( i_14_  &  i_13_  &  (~ i_12_)  &  i_15_ ) ;
 assign _36030 = ( i_14_  &  (~ i_13_)  &  (~ i_12_) ) ;
 assign _36035 = ( n_n57  &  wire153 ) | ( n_n57  &  wire166 ) ;
 assign _36055 = ( wire273  &  n_n57 ) | ( n_n57  &  wire157 ) ;
 assign _36064 = ( wire704 ) | ( wire19720 ) | ( _36035 ) | ( _36055 ) ;
 assign _36066 = ( n_n4967 ) | ( wire613 ) | ( wire19730 ) | ( wire19732 ) ;
 assign _36068 = ( wire19717 ) | ( wire19718 ) | ( wire19735 ) | ( _36066 ) ;
 assign _36083 = ( wire5363 ) | ( wire5361 ) ;
 assign _36085 = ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire900 ) | ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  wire900 ) ;
 assign _36086 = ( i_14_  &  i_13_  &  i_12_  &  wire906 ) | ( (~ i_14_)  &  i_13_  &  i_12_  &  wire906 ) | ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire906 ) | ( i_14_  &  i_13_  &  (~ i_12_)  &  wire906 ) ;
 assign _36087 = ( n_n6  &  n_n42 ) | ( n_n6  &  _36085 ) | ( n_n6  &  _36086 ) ;
 assign _36090 = ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  wire904 ) | ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire904 ) ;
 assign _36091 = ( n_n5  &  n_n49 ) | ( n_n5  &  wire807 ) | ( n_n5  &  _36090 ) ;
 assign _36092 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  i_15_ ) ;
 assign _36093 = ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  (~ i_15_) ) ;
 assign _36095 = ( (~ i_14_)  &  i_13_  &  i_12_ ) ;
 assign _36096 = ( (~ i_14_)  &  i_13_  &  i_12_  &  wire912 ) | ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire912 ) ;
 assign _36098 = ( (~ i_14_)  &  i_13_  &  i_12_  &  (~ i_15_) ) ;
 assign _36099 = ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  i_15_ ) ;
 assign _36101 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire914 ) ;
 assign _36107 = ( i_14_  &  i_13_  &  (~ i_12_) ) ;
 assign _36112 = ( i_14_  &  i_13_  &  i_12_  &  (~ i_15_) ) ;
 assign _36113 = ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  i_15_ ) ;
 assign _36115 = ( i_14_  &  (~ i_13_)  &  (~ i_12_) ) ;
 assign _36116 = ( i_14_  &  i_13_  &  (~ i_12_)  &  wire907 ) | ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire907 ) ;
 assign _36121 = ( n_n1506 ) | ( _5624 ) | ( _36087 ) ;
 assign _36122 = ( n_n4330 ) | ( wire19671 ) | ( _36083 ) | ( _36121 ) ;
 assign _36137 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_ ) ;
 assign _36138 = ( (~ i_14_)  &  i_13_  &  i_12_  &  (~ i_15_) ) ;
 assign _36139 = ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  i_15_ ) ;
 assign _36140 = ( wire906  &  _35091 ) | ( wire905  &  _36137 ) ;
 assign _36143 = ( (~ i_14_)  &  i_13_  &  i_12_  &  i_15_ ) ;
 assign _36144 = ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  (~ i_15_) ) ;
 assign _36149 = ( wire5268 ) | ( wire5269 ) | ( wire5262 ) | ( _5578 ) ;
 assign _36150 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire899 ) ;
 assign _36156 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_ ) ;
 assign _36157 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire913 ) | ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire913 ) ;
 assign _36159 = ( n_n5  &  wire52 ) | ( wire911  &  n_n5  &  _34580 ) ;
 assign _36161 = ( wire911  &  _34580 ) | ( wire913  &  _35938 ) ;
 assign _36165 = ( wire699 ) | ( n_n4838 ) | ( _5559 ) | ( _36159 ) ;
 assign _36168 = ( i_14_  &  i_13_  &  i_12_ ) ;
 assign _36176 = ( wire19742 ) | ( wire19747 ) | ( _36149 ) | ( _36165 ) ;
 assign _36179 = ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  i_15_ ) ;
 assign _36180 = ( i_14_  &  (~ i_13_)  &  i_12_  &  (~ i_15_) ) ;
 assign _36184 = ( i_14_  &  i_13_  &  i_12_ ) ;
 assign _36190 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire908 ) | ( i_14_  &  i_13_  &  (~ i_12_)  &  wire908 ) ;
 assign _36192 = ( n_n5  &  wire61 ) | ( n_n5  &  wire908  &  _35212 ) ;
 assign _36193 = ( wire903  &  _35109 ) | ( wire897  &  _35124 ) ;
 assign _36195 = ( wire899  &  _34575 ) | ( wire897  &  _35103 ) ;
 assign _36198 = ( n_n4846 ) | ( n_n4842 ) | ( _5503 ) | ( _36192 ) ;
 assign _36202 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_ ) ;
 assign _36203 = ( wire912  &  _36095 ) | ( wire914  &  _36202 ) ;
 assign _36205 = ( i_14_  &  i_13_  &  (~ i_12_)  &  wire908 ) | ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire908 ) ;
 assign _36210 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_ ) ;
 assign _36212 = ( (~ i_14_)  &  i_13_  &  (~ i_12_) ) ;
 assign _36215 = ( n_n285  &  n_n230  &  n_n263 ) ;
 assign _36218 = ( n_n285  &  n_n230  &  n_n261 ) ;
 assign _36219 = ( wire55  &  _36215 ) | ( wire56  &  _36218 ) ;
 assign _36222 = ( wire5240 ) | ( wire5241 ) | ( _5480 ) | ( _5481 ) ;
 assign _36224 = ( wire912  &  _34544 ) | ( wire907  &  _36210 ) ;
 assign _36227 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire897 ) ;
 assign _36229 = ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  wire907 ) ;
 assign _36231 = ( n_n5  &  wire19407 ) | ( n_n5  &  _36227 ) | ( n_n5  &  _36229 ) ;
 assign _36234 = ( wire19659 ) | ( wire19755 ) | ( _36198 ) | ( _36222 ) ;
 assign _36235 = ( wire19677 ) | ( wire19761 ) | ( _36122 ) | ( _36176 ) ;
 assign _36238 = ( n_n3255 ) | ( wire5725 ) | ( wire5726 ) | ( _5470 ) ;
 assign _36242 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire907 ) | ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire907 ) ;
 assign _36244 = ( n_n1  &  wire89 ) | ( wire907  &  n_n1  &  _36107 ) ;
 assign _36245 = ( wire912  &  _34544 ) | ( wire907  &  _36210 ) ;
 assign _36249 = ( n_n1  &  n_n32 ) | ( n_n2  &  n_n32 ) | ( n_n1  &  wire85 ) ;
 assign _36250 = ( n_n3257 ) | ( _5462 ) | ( _36244 ) | ( _36249 ) ;
 assign _36253 = ( n_n260  &  n_n273  &  n_n285 ) ;
 assign _36255 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_ ) ;
 assign _36256 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire899 ) | ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire899 ) ;
 assign _36264 = ( n_n3523 ) | ( wire5720 ) | ( wire5721 ) | ( _5446 ) ;
 assign _36265 = ( wire905  &  _36137 ) | ( wire899  &  _36255 ) ;
 assign _36267 = ( n_n1  &  wire42 ) | ( n_n1  &  wire899  &  _34575 ) ;
 assign _36270 = ( wire911  &  _34580 ) | ( wire913  &  _35938 ) ;
 assign _36273 = ( wire468 ) | ( wire913  &  n_n220  &  n_n2 ) ;
 assign _36275 = ( wire902  &  _35056 ) | ( wire900  &  _35074 ) ;
 assign _36277 = ( n_n1  &  wire113 ) | ( n_n1  &  wire912  &  _36184 ) ;
 assign _36282 = ( wire5205 ) | ( wire19780 ) ;
 assign _36285 = ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire900 ) | ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  wire900 ) ;
 assign _36286 = ( i_14_  &  i_13_  &  i_12_  &  wire906 ) | ( (~ i_14_)  &  i_13_  &  i_12_  &  wire906 ) | ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire906 ) | ( i_14_  &  i_13_  &  (~ i_12_)  &  wire906 ) ;
 assign _36289 = ( n_n3786 ) | ( n_n3782 ) | ( wire723 ) | ( _5408 ) ;
 assign _36291 = ( wire904  &  _35153 ) | ( wire907  &  _36107 ) ;
 assign _36293 = ( n_n2  &  wire85 ) | ( n_n2  &  wire904  &  _35137 ) ;
 assign _36297 = ( n_n3260 ) | ( _5392 ) | ( _5399 ) | ( _36293 ) ;
 assign _36298 = ( n_n1  &  wire71 ) | ( n_n1  &  wire904  &  _35153 ) ;
 assign _36304 = ( wire902  &  _35056 ) | ( wire911  &  _36168 ) ;
 assign _36308 = ( wire913  &  _35004 ) | ( wire911  &  _36168 ) ;
 assign _36311 = ( wire5160 ) | ( wire5161 ) | ( _5376 ) | ( _5377 ) ;
 assign _36312 = ( n_n2579 ) | ( n_n2580 ) | ( wire19778 ) | ( wire19821 ) ;
 assign _36315 = ( wire48  &  n_n122 ) | ( wire905  &  n_n122  &  _34956 ) ;
 assign _36317 = ( _6592 ) | ( wire913  &  n_n220 ) | ( n_n220  &  wire905 ) ;
 assign _36319 = ( wire364 ) | ( _5357 ) | ( _5359 ) | ( _36315 ) ;
 assign _36324 = ( wire5442 ) | ( wire5441 ) ;
 assign _36330 = ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_) ) ;
 assign _36331 = ( wire912  &  _35754 ) | ( wire911  &  _36330 ) ;
 assign _36334 = ( wire583 ) | ( wire19825 ) | ( wire19837 ) | ( _36324 ) ;
 assign _36335 = ( wire19835 ) | ( wire19830 ) | ( _36319 ) | ( _36334 ) ;
 assign _36337 = ( i_14_  &  (~ i_13_)  &  i_12_ ) ;
 assign _36339 = ( i_14_  &  (~ i_13_)  &  i_12_ ) ;
 assign _36341 = ( i_14_  &  i_13_  &  i_12_  &  wire902 ) ;
 assign _36343 = ( i_14_  &  (~ i_13_)  &  i_12_ ) ;
 assign _36360 = ( i_14_  &  (~ i_13_)  &  i_12_ ) ;
 assign _36375 = ( wire19846 ) | ( wire19847 ) ;
 assign _36377 = ( wire911  &  _34580 ) | ( wire913  &  _35938 ) ;
 assign _36380 = ( n_n268  &  wire124 ) | ( n_n268  &  wire212 ) ;
 assign _36382 = ( i_14_  &  (~ i_13_)  &  (~ i_12_) ) ;
 assign _36383 = ( wire912  &  _34544 ) | ( wire914  &  _36382 ) ;
 assign _36392 = ( wire19854 ) | ( _5309 ) | ( _5310 ) | ( _36380 ) ;
 assign _36393 = ( n_n2550 ) | ( n_n2545 ) | ( wire19859 ) | ( _36392 ) ;
 assign _36396 = ( wire911  &  _34580 ) | ( wire913  &  _35938 ) ;
 assign _36404 = ( n_n4913 ) | ( n_n4915 ) | ( n_n4914 ) | ( _5274 ) ;
 assign _36405 = ( n_n57  &  wire140 ) | ( n_n57  &  wire165 ) ;
 assign _36410 = ( i_5_  &  i_3_  &  i_4_ ) ;
 assign _36417 = ( wire761 ) | ( wire19931 ) | ( _36405 ) ;
 assign _36421 = ( wire913  &  n_n220 ) | ( n_n220  &  wire905 ) ;
 assign _36424 = ( _5227 ) | ( wire48  &  n_n130 ) | ( n_n130  &  _5244 ) ;
 assign _36426 = ( n_n285  &  n_n271  &  n_n230 ) ;
 assign _36428 = ( n_n5796 ) | ( _5225 ) | ( wire224  &  _36426 ) ;
 assign _36430 = ( wire905  &  _34956 ) | ( wire913  &  _35748 ) ;
 assign _36442 = ( n_n5796 ) | ( wire452 ) | ( wire5812 ) ;
 assign _36443 = ( n_n5664 ) | ( n_n5679 ) | ( wire587 ) | ( wire5813 ) ;
 assign _36448 = ( n_n4489 ) | ( wire507 ) ;
 assign _36450 = ( wire19953 ) | ( wire19952 ) | ( _5218 ) | ( _5219 ) ;
 assign _36453 = ( n_n285  &  n_n271  &  n_n230 ) ;
 assign _36457 = ( n_n4955 ) | ( wire19977 ) | ( wire277  &  _36453 ) ;
 assign _36461 = ( n_n56  &  wire166 ) | ( n_n56  &  wire180 ) ;
 assign _36467 = ( wire901  &  _35946 ) | ( wire905  &  _36137 ) ;
 assign _36469 = ( n_n5  &  wire73 ) | ( n_n5  &  wire906  &  _35091 ) ;
 assign _36474 = ( wire573 ) | ( wire5076 ) | ( _5183 ) | ( _36469 ) ;
 assign _36475 = ( n_n6  &  wire19738 ) | ( wire913  &  n_n6  &  _36156 ) ;
 assign _36476 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire913 ) | ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire913 ) ;
 assign _36480 = ( wire5268 ) | ( wire5269 ) | ( _5179 ) | ( _36475 ) ;
 assign _36482 = ( i_14_  &  i_13_  &  i_12_  &  wire902 ) ;
 assign _36483 = ( n_n5  &  wire63 ) | ( n_n5  &  wire1874 ) | ( n_n5  &  _36482 ) ;
 assign _36487 = ( wire585 ) | ( wire5059 ) | ( wire5400 ) | ( _36483 ) ;
 assign _36488 = ( wire19878 ) | ( wire19882 ) | ( _36474 ) | ( _36480 ) ;
 assign _36489 = ( wire911  &  _34580 ) | ( wire908  &  _35212 ) ;
 assign _36491 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire908 ) | ( i_14_  &  i_13_  &  (~ i_12_)  &  wire908 ) ;
 assign _36495 = ( n_n4838 ) | ( n_n6  &  wire66 ) | ( n_n6  &  _36150 ) ;
 assign _36501 = ( wire5238 ) | ( wire5239 ) | ( wire5048 ) | ( _5158 ) ;
 assign _36502 = ( n_n6  &  wire53 ) | ( n_n6  &  wire897  &  _35103 ) ;
 assign _36506 = ( wire5240 ) | ( wire5241 ) | ( _5150 ) | ( _36502 ) ;
 assign _36508 = ( n_n4730 ) | ( wire19900 ) | ( wire19906 ) | ( _36501 ) ;
 assign _36510 = ( n_n206  &  n_n56 ) | ( n_n56  &  wire908  &  _35033 ) ;
 assign _36515 = ( wire5035 ) | ( wire5031 ) | ( _5145 ) | ( _36510 ) ;
 assign _36518 = ( wire905  &  _36137 ) | ( wire899  &  _36255 ) ;
 assign _36525 = ( n_n285  &  n_n266  &  n_n230 ) ;
 assign _36536 = ( n_n5  &  wire86 ) | ( wire907  &  n_n5  &  _36210 ) ;
 assign _36542 = ( wire5244 ) | ( wire5245 ) | ( _5101 ) | ( _36536 ) ;
 assign _36544 = ( n_n285  &  n_n230  &  n_n261 ) ;
 assign _36548 = ( wire632 ) | ( wire5613 ) | ( wire99  &  _36544 ) ;
 assign _36550 = ( wire674 ) | ( wire224  &  _35255 ) ;
 assign _36555 = ( wire19865 ) | ( wire19868 ) | ( _36542 ) | ( _36548 ) ;
 assign _36558 = ( wire19872 ) | ( wire19921 ) | ( wire19987 ) | ( _36555 ) ;
 assign _36563 = ( i_6_  &  i_7_ ) ;
 assign _36585 = ( (~ i_5_)  &  (~ i_3_)  &  (~ i_4_) ) ;
 assign _36611 = ( wire20002 ) | ( wire20004 ) | ( wire535 ) | ( wire20000 ) ;
 assign _36614 = ( n_n124  &  wire1686 ) | ( n_n132  &  wire1686 ) ;
 assign _36616 = ( n_n152  &  wire266 ) | ( n_n152  &  wire1705 ) ;
 assign _36619 = ( wire20007 ) | ( wire20008 ) | ( _36614 ) | ( _36616 ) ;
 assign _36620 = ( wire4905 ) | ( wire20011 ) | ( _5028 ) | ( _36619 ) ;
 assign _36682 = ( i_14_  &  (~ i_13_)  &  i_12_  &  wire912 ) ;
 assign _36683 = ( i_14_  &  i_13_  &  (~ i_12_)  &  i_15_ ) ;
 assign _36687 = ( n_n100  &  wire167 ) | ( n_n100  &  wire198 ) ;
 assign _36698 = ( n_n260  &  n_n285  &  n_n261 ) ;
 assign _36699 = ( (~ i_9_)  &  i_10_  &  (~ i_11_)  &  i_15_ ) ;
 assign _36705 = ( i_14_  &  i_13_  &  (~ i_12_) ) ;
 assign _36714 = ( wire20068 ) | ( wire1662  &  _36698 ) ;
 assign _36783 = ( i_14_  &  i_13_  &  i_12_ ) ;
 assign _36786 = ( i_14_  &  (~ i_13_)  &  i_12_ ) ;
 assign _36788 = ( i_14_  &  (~ i_13_)  &  (~ i_12_) ) ;
 assign _36790 = ( i_14_  &  i_13_  &  (~ i_12_) ) ;
 assign _36797 = ( wire877 ) | ( wire4805 ) | ( wire20081 ) | ( _4920 ) ;
 assign _36803 = ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  wire905 ) ;
 assign _36807 = ( (~ i_14_)  &  i_13_  &  i_12_ ) ;
 assign _36808 = ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire911 ) ;
 assign _36810 = ( (~ i_14_)  &  i_13_  &  i_12_ ) ;
 assign _36813 = ( n_n2713 ) | ( wire4789 ) | ( wire20100 ) | ( _4901 ) ;
 assign _36817 = ( i_14_  &  i_13_  &  i_12_ ) ;
 assign _36818 = ( n_n94  &  wire246 ) | ( wire901  &  n_n94  &  _36817 ) ;
 assign _36821 = ( wire904  &  _35427 ) | ( wire898  &  _35480 ) ;
 assign _36824 = ( n_n2724 ) | ( _4868 ) | ( _4878 ) | ( _36818 ) ;
 assign _36825 = ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  wire912 ) ;
 assign _36826 = ( wire902  &  _35056 ) | ( wire899  &  _35953 ) ;
 assign _36833 = ( i_14_  &  (~ i_13_)  &  i_12_ ) ;
 assign _36844 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_ ) ;
 assign _36856 = ( (~ i_14_)  &  i_13_  &  i_12_ ) ;
 assign _36865 = ( n_n2657 ) | ( n_n2665 ) | ( wire20073 ) | ( _36714 ) ;
 assign _36876 = ( i_14_  &  i_13_  &  (~ i_12_)  &  wire907 ) | ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire907 ) ;
 assign _36878 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire907 ) | ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire907 ) ;
 assign _36881 = ( n_n56  &  wire57 ) | ( wire912  &  n_n56  &  _34544 ) ;
 assign _36887 = ( _4792 ) | ( _6055 ) | ( _35579 ) | ( _36881 ) ;
 assign _36888 = ( _4798 ) | ( _4799 ) | ( _6077 ) | ( _35565 ) ;
 assign _36889 = ( wire4655 ) | ( wire20199 ) | ( wire20200 ) | ( _36888 ) ;
 assign _36890 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire900 ) | ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire900 ) ;
 assign _36894 = ( n_n4680 ) | ( n_n4677 ) | ( n_n4685 ) | ( _4782 ) ;
 assign _36895 = ( wire911  &  _34580 ) | ( wire913  &  _35938 ) ;
 assign _36909 = ( i_14_  &  (~ i_13_)  &  (~ i_12_) ) ;
 assign _36912 = ( n_n130  &  wire1545 ) | ( (~ i_9_)  &  (~ i_10_)  &  n_n130 ) ;
 assign _36916 = ( n_n57  &  wire96 ) | ( n_n57  &  wire904  &  _35141 ) ;
 assign _36947 = ( wire20192 ) | ( wire4636 ) | ( _36912 ) | ( _36916 ) ;
 assign _36950 = ( n_n4556 ) | ( wire20240 ) | ( wire20209 ) | ( _36889 ) ;
 assign _36951 = ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  wire913 ) ;
 assign _36952 = ( wire75  &  n_n56 ) | ( wire118  &  n_n56 ) | ( n_n56  &  _36951 ) ;
 assign _36954 = ( n_n285  &  n_n271  &  n_n230 ) ;
 assign _36957 = ( wire5033 ) | ( wire5031 ) | ( _36510 ) | ( _36952 ) ;
 assign _36958 = ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  wire914 ) ;
 assign _36959 = ( wire95  &  n_n57 ) | ( n_n57  &  wire101 ) | ( n_n57  &  _36958 ) ;
 assign _36964 = ( (~ i_14_)  &  i_13_  &  i_12_  &  wire898 ) | ( i_14_  &  i_13_  &  (~ i_12_)  &  wire898 ) ;
 assign _36967 = ( wire900  &  _35644 ) | ( wire906  &  _35685 ) ;
 assign _36969 = ( i_14_  &  i_13_  &  i_12_  &  wire906 ) | ( i_14_  &  i_13_  &  (~ i_12_)  &  wire906 ) ;
 assign _36971 = ( wire4750 ) | ( n_n6  &  _35235 ) | ( n_n6  &  _35236 ) ;
 assign _36972 = ( wire20117 ) | ( _4701 ) | ( _4702 ) | ( _4706 ) ;
 assign _36973 = ( wire20119 ) | ( _36957 ) | ( _36971 ) | ( _36972 ) ;
 assign _36974 = ( (~ i_14_)  &  i_13_  &  i_12_  &  i_15_ ) ;
 assign _36975 = ( i_14_  &  i_13_  &  (~ i_12_)  &  (~ i_15_) ) ;
 assign _36977 = ( (~ i_14_)  &  i_13_  &  i_12_ ) ;
 assign _36982 = ( (~ i_14_)  &  i_13_  &  i_12_  &  wire914 ) | ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire914 ) ;
 assign _36984 = ( wire914  &  n_n6  &  _34952 ) | ( wire914  &  n_n6  &  _36202 ) ;
 assign _36986 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_ ) ;
 assign _36988 = ( (~ i_14_)  &  i_13_  &  i_12_ ) ;
 assign _36993 = ( (~ i_14_)  &  i_13_  &  i_12_  &  wire901 ) | ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire901 ) ;
 assign _36995 = ( i_14_  &  (~ i_13_)  &  i_12_  &  wire901 ) | ( i_14_  &  i_13_  &  (~ i_12_)  &  wire901 ) ;
 assign _37000 = ( (~ i_14_)  &  i_13_  &  i_12_  &  wire901 ) | ( i_14_  &  i_13_  &  (~ i_12_)  &  wire901 ) ;
 assign _37002 = ( _4687 ) | ( _4688 ) | ( _4694 ) | ( _36984 ) ;
 assign _37003 = ( i_14_  &  (~ i_13_)  &  i_12_  &  wire902 ) | ( i_14_  &  i_13_  &  (~ i_12_)  &  wire902 ) ;
 assign _37004 = ( n_n6  &  wire86 ) | ( n_n6  &  wire901  &  _36986 ) ;
 assign _37013 = ( i_14_  &  i_13_  &  i_12_  &  (~ i_15_) ) ;
 assign _37014 = ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  i_15_ ) ;
 assign _37022 = ( i_14_  &  (~ i_13_)  &  i_12_ ) ;
 assign _37024 = ( i_14_  &  i_13_  &  i_12_  &  wire906 ) | ( i_14_  &  i_13_  &  (~ i_12_)  &  wire906 ) ;
 assign _37026 = ( n_n6  &  wire59 ) | ( n_n6  &  wire906  &  _35685 ) ;
 assign _37027 = ( (~ i_14_)  &  i_13_  &  i_12_  &  wire898 ) | ( i_14_  &  i_13_  &  (~ i_12_)  &  wire898 ) ;
 assign _37030 = ( n_n1505 ) | ( _4643 ) | ( _4653 ) | ( _37026 ) ;
 assign _37032 = ( wire902  &  n_n222 ) | ( wire911  &  _36343 ) ;
 assign _37035 = ( n_n5  &  wire20149 ) | ( n_n5  &  n_n222  &  _36699 ) ;
 assign _37037 = ( (~ i_14_)  &  i_13_  &  i_12_  &  wire902 ) | ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire902 ) ;
 assign _37042 = ( i_14_  &  i_13_  &  (~ i_12_) ) ;
 assign _37043 = ( i_14_  &  i_13_  &  i_12_  &  (~ i_15_) ) ;
 assign _37044 = ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  i_15_ ) ;
 assign _37046 = ( i_14_  &  i_13_  &  (~ i_12_) ) ;
 assign _37047 = ( wire899  &  _37042 ) | ( wire905  &  _37046 ) ;
 assign _37050 = ( wire4711 ) | ( _4631 ) | ( _4635 ) | ( _37035 ) ;
 assign _37057 = ( wire911  &  _36807 ) | ( wire913  &  _36810 ) ;
 assign _37063 = ( wire911  &  n_n258 ) | ( n_n222  &  _36699 ) ;
 assign _37064 = ( wire899  &  _37042 ) | ( wire905  &  _37046 ) ;
 assign _37066 = ( _4609 ) | ( _4610 ) | ( _4614 ) | ( _4615 ) ;
 assign _37068 = ( wire902  &  _35422 ) | ( wire903  &  _35626 ) ;
 assign _37070 = ( wire897  &  _35539 ) | ( wire903  &  _35628 ) ;
 assign _37072 = ( (~ i_14_)  &  i_13_  &  i_12_  &  wire903 ) | ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire903 ) ;
 assign _37074 = ( n_n6  &  wire40 ) | ( n_n6  &  wire897  &  _35544 ) ;
 assign _37076 = ( _4596 ) | ( _4599 ) | ( _4600 ) | ( _37074 ) ;
 assign _37077 = ( wire20153 ) | ( wire20157 ) | ( _37050 ) | ( _37066 ) ;
 assign _37084 = ( wire903  &  _35190 ) | ( wire912  &  _36184 ) ;
 assign _37086 = ( n_n5  &  wire113 ) | ( wire914  &  n_n5  &  _34565 ) ;
 assign _37087 = ( wire897  &  _35039 ) | ( wire907  &  _36833 ) ;
 assign _37089 = ( n_n6  &  wire199 ) | ( n_n6  &  wire901  &  _36817 ) ;
 assign _37091 = ( i_14_  &  i_13_  &  i_12_ ) ;
 assign _37093 = ( _4582 ) | ( _4585 ) | ( _37086 ) | ( _37089 ) ;
 assign _37095 = ( n_n6  &  wire246 ) | ( wire914  &  n_n6  &  _34565 ) ;
 assign _37097 = ( wire900  &  _35074 ) | ( wire904  &  _35391 ) ;
 assign _37099 = ( n_n5  &  wire101 ) | ( n_n5  &  wire20180 ) ;
 assign _37104 = ( n_n4605 ) | ( wire4691 ) | ( _4567 ) | ( _37099 ) ;
 assign _37105 = ( wire4694 ) | ( wire4695 ) | ( _4574 ) | ( _37095 ) ;
 assign _37106 = ( wire20176 ) | ( _37093 ) | ( _37105 ) ;
 assign _37108 = ( n_n4549 ) | ( wire20184 ) | ( _36973 ) | ( _37106 ) ;
 assign _37110 = ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  wire901 ) ;
 assign _37116 = ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  wire912 ) ;
 assign _37128 = ( (~ i_14_)  &  i_13_  &  i_12_  &  wire902 ) | ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire902 ) ;
 assign _37130 = ( wire88  &  n_n48 ) | ( wire902  &  n_n48  &  _35420 ) ;
 assign _37140 = ( wire4587 ) | ( wire20259 ) | ( _4485 ) | ( _37130 ) ;
 assign _37141 = ( wire897  &  _35539 ) | ( wire903  &  _35628 ) ;
 assign _37143 = ( n_n48  &  wire104 ) | ( n_n48  &  wire903  &  _35626 ) ;
 assign _37148 = ( wire897  &  _35539 ) | ( wire903  &  _35626 ) ;
 assign _37155 = ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  wire908 ) ;
 assign _37158 = ( i_14_  &  i_13_  &  i_12_  &  wire901 ) ;
 assign _37160 = ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  wire907 ) ;
 assign _37161 = ( i_14_  &  i_13_  &  i_12_  &  wire902 ) ;
 assign _37163 = ( i_14_  &  (~ i_13_)  &  i_12_ ) ;
 assign _37168 = ( n_n222  &  _36699 ) | ( wire911  &  _36807 ) ;
 assign _37170 = ( n_n53  &  wire62 ) | ( n_n53  &  wire20155 ) | ( n_n53  &  _4432 ) ;
 assign _37178 = ( wire904  &  _35391 ) | ( wire899  &  _37042 ) ;
 assign _37180 = ( n_n281  &  wire906 ) | ( wire899  &  _36255 ) ;
 assign _37189 = ( (~ i_14_)  &  i_13_  &  i_12_  &  wire898 ) | ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire898 ) ;
 assign _37191 = ( n_n53  &  wire96 ) | ( wire898  &  n_n53  &  _35693 ) ;
 assign _37204 = ( i_14_  &  i_13_  &  i_12_  &  wire906 ) | ( i_14_  &  i_13_  &  (~ i_12_)  &  wire906 ) ;
 assign _37208 = ( wire20300 ) | ( wire20301 ) | ( _4401 ) | ( _37191 ) ;
 assign _37209 = ( (~ i_14_)  &  i_13_  &  i_12_  &  wire914 ) | ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire914 ) ;
 assign _37211 = ( n_n53  &  wire368 ) | ( n_n53  &  n_n247  &  _36683 ) ;
 assign _37215 = ( (~ i_14_)  &  i_13_  &  i_12_  &  wire901 ) | ( i_14_  &  i_13_  &  (~ i_12_)  &  wire901 ) ;
 assign _37220 = ( n_n4174 ) | ( wire20310 ) | ( _4385 ) | ( _37211 ) ;
 assign _37222 = ( wire906  &  _35685 ) | ( wire898  &  _35693 ) ;
 assign _37224 = ( (~ i_14_)  &  i_13_  &  i_12_  &  wire898 ) | ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire898 ) ;
 assign _37226 = ( i_14_  &  i_13_  &  i_12_  &  wire906 ) | ( (~ i_14_)  &  i_13_  &  i_12_  &  wire906 ) ;
 assign _37227 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire900 ) | ( i_14_  &  i_13_  &  (~ i_12_)  &  wire900 ) | ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire900 ) | ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  wire900 ) ;
 assign _37228 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire906 ) | ( i_14_  &  i_13_  &  (~ i_12_)  &  wire906 ) | ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  wire906 ) ;
 assign _37230 = ( n_n4179 ) | ( wire809 ) | ( _4370 ) | ( _4371 ) ;
 assign _37231 = ( wire20304 ) | ( wire4530 ) | ( _37208 ) | ( _37220 ) ;
 assign _37244 = ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  wire913 ) ;
 assign _37247 = ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  wire903 ) ;
 assign _37253 = ( wire902  &  n_n53  &  _35420 ) | ( wire902  &  n_n53  &  _35422 ) ;
 assign _37256 = ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire899 ) ;
 assign _37263 = ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  wire902 ) ;
 assign _37273 = ( wire906  &  _35685 ) | ( wire901  &  _36986 ) ;
 assign _37275 = ( n_n6  &  wire51 ) | ( n_n6  &  wire912  &  _37022 ) ;
 assign _37277 = ( _4362 ) | ( _4694 ) | ( _36984 ) | ( _37275 ) ;
 assign _37280 = ( i_14_  &  (~ i_13_)  &  i_12_  &  wire902 ) | ( i_14_  &  i_13_  &  (~ i_12_)  &  wire902 ) ;
 assign _37284 = ( wire4435 ) | ( wire20437 ) | ( _4348 ) | ( _4349 ) ;
 assign _37285 = ( n_n6  &  wire71 ) | ( n_n6  &  wire898  &  _35711 ) ;
 assign _37286 = ( i_14_  &  (~ i_13_)  &  i_12_  &  wire907 ) ;
 assign _37291 = ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_) ) ;
 assign _37296 = ( wire20435 ) | ( wire20442 ) | ( _37277 ) | ( _37284 ) ;
 assign _37297 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire914 ) | ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  wire914 ) ;
 assign _37298 = ( n_n53  &  wire245 ) | ( wire912  &  n_n53  &  _36095 ) ;
 assign _37300 = ( i_14_  &  i_13_  &  (~ i_12_)  &  wire907 ) | ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire907 ) ;
 assign _37303 = ( _4324 ) | ( _4514 ) | ( _37253 ) | ( _37298 ) ;
 assign _37304 = ( wire897  &  _35039 ) | ( wire911  &  _36168 ) ;
 assign _37314 = ( wire912  &  _34544 ) | ( wire906  &  _35186 ) ;
 assign _37316 = ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire900 ) | ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  wire900 ) ;
 assign _37317 = ( i_14_  &  i_13_  &  i_12_  &  wire906 ) | ( (~ i_14_)  &  i_13_  &  i_12_  &  wire906 ) | ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire906 ) | ( i_14_  &  i_13_  &  (~ i_12_)  &  wire906 ) ;
 assign _37320 = ( wire20469 ) | ( _4310 ) | ( _4311 ) | ( _4312 ) ;
 assign _37321 = ( wire20457 ) | ( wire4409 ) | ( wire20474 ) | ( _37303 ) ;
 assign _37322 = ( wire913  &  n_n281 ) | ( wire911  &  _36168 ) ;
 assign _37323 = ( n_n53  &  wire50 ) | ( n_n53  &  wire897  &  _35039 ) ;
 assign _37326 = ( i_14_  &  (~ i_13_)  &  i_12_  &  wire905 ) ;
 assign _37333 = ( wire900  &  _35074 ) | ( wire913  &  _35748 ) ;
 assign _37335 = ( wire911  &  _34580 ) | ( wire906  &  _35091 ) ;
 assign _37340 = ( i_14_  &  i_13_  &  i_12_  &  wire901 ) ;
 assign _37341 = ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  wire905 ) ;
 assign _37346 = ( wire903  &  _35101 ) | ( wire897  &  _35103 ) ;
 assign _37348 = ( wire406 ) | ( n_n53  &  wire42 ) | ( n_n53  &  _37256 ) ;
 assign _37350 = ( wire4453 ) | ( wire20429 ) | ( wire20430 ) | ( wire20422 ) ;
 assign _37351 = ( wire4463 ) | ( wire20479 ) | ( wire20480 ) | ( _37348 ) ;
 assign _37352 = ( wire20452 ) | ( _37296 ) | ( _37320 ) | ( _37321 ) ;
 assign _37358 = ( wire899  &  _36255 ) | ( wire905  &  _37046 ) ;
 assign _37360 = ( n_n100  &  wire469 ) | ( wire899  &  n_n100  &  _37042 ) ;
 assign _37361 = ( wire911  &  _36807 ) | ( wire913  &  _36810 ) ;
 assign _37363 = ( n_n100  &  wire62 ) | ( wire898  &  n_n100  &  _35396 ) ;
 assign _37367 = ( _4249 ) | ( _4252 ) | ( _37360 ) | ( _37363 ) ;
 assign _37370 = ( wire911  &  _36168 ) | ( wire905  &  _36337 ) ;
 assign _37373 = ( i_14_  &  i_13_  &  i_12_  &  wire899 ) ;
 assign _37375 = ( i_14_  &  (~ i_13_)  &  i_12_  &  wire907 ) ;
 assign _37376 = ( n_n60  &  n_n100 ) | ( n_n100  &  _37373 ) | ( n_n100  &  _37375 ) ;
 assign _37378 = ( wire370 ) | ( wire20516 ) | ( wire20501 ) | ( wire20502 ) ;
 assign _37379 = ( wire4360 ) | ( wire20508 ) | ( _37367 ) ;
 assign _37380 = ( (~ i_14_)  &  i_13_  &  i_12_  &  wire914 ) | ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire914 ) | ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  wire914 ) ;
 assign _37381 = ( n_n100  &  wire102 ) | ( wire914  &  n_n100  &  _36382 ) ;
 assign _37382 = ( wire906  &  _35685 ) | ( wire901  &  _36986 ) ;
 assign _37390 = ( wire20532 ) | ( wire20533 ) | ( _4226 ) | ( _37381 ) ;
 assign _37396 = ( n_n177  &  n_n35 ) | ( wire913  &  n_n177  &  _35938 ) ;
 assign _37398 = ( wire20519 ) | ( wire628 ) ;
 assign _37406 = ( _4180 ) | ( wire40  &  n_n100 ) | ( n_n100  &  _4189 ) ;
 assign _37407 = ( wire20541 ) | ( wire4344 ) | ( _37390 ) ;
 assign _37409 = ( (~ i_14_)  &  i_13_  &  i_12_  &  wire912 ) | ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire912 ) ;
 assign _37411 = ( n_n57  &  wire453 ) | ( wire914  &  n_n57  &  _36202 ) ;
 assign _37415 = ( wire460 ) | ( wire4391 ) | ( wire20486 ) | ( _4170 ) ;
 assign _37416 = ( wire900  &  _35074 ) | ( wire913  &  _35748 ) ;
 assign _37422 = ( n_n4913 ) | ( n_n4914 ) | ( _4165 ) | ( _4166 ) ;
 assign _37424 = ( wire903  &  _35101 ) | ( wire897  &  _35103 ) ;
 assign _37426 = ( i_14_  &  (~ i_13_)  &  i_12_  &  wire897 ) | ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire897 ) | ( i_14_  &  i_13_  &  (~ i_12_)  &  wire897 ) ;
 assign _37428 = ( _4155 ) | ( _4156 ) | ( _4160 ) | ( _4161 ) ;
 assign _37429 = ( wire653 ) | ( wire20549 ) | ( _37415 ) | ( _37428 ) ;
 assign _37432 = ( n_n6  &  wire79 ) | ( n_n6  &  wire899  &  _36255 ) ;
 assign _37433 = ( wire898  &  _35396 ) | ( wire913  &  _36810 ) ;
 assign _37435 = ( wire904  &  _35391 ) | ( wire911  &  _36807 ) ;
 assign _37438 = ( wire411 ) | ( wire647 ) | ( _4149 ) | ( _37432 ) ;
 assign _37442 = ( i_14_  &  i_13_  &  i_12_  &  (~ i_15_) ) ;
 assign _37444 = ( (~ i_14_)  &  i_13_  &  i_12_  &  i_15_ ) ;
 assign _37445 = ( wire897  &  _35103 ) | ( wire903  &  _35628 ) ;
 assign _37448 = ( i_14_  &  (~ i_13_)  &  i_12_  &  wire905 ) ;
 assign _37463 = ( n_n2876 ) | ( n_n2875 ) | ( wire20374 ) | ( wire20381 ) ;
 assign _37464 = ( wire20382 ) | ( _4147 ) | ( _4148 ) | ( _37438 ) ;
 assign _37469 = ( i_14_  &  (~ i_13_)  &  i_12_  &  wire899 ) ;
 assign _37480 = ( i_14_  &  i_13_  &  (~ i_12_)  &  wire905 ) ;
 assign _37495 = ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  wire906 ) ;
 assign _37496 = ( n_n4  &  n_n65 ) | ( n_n4  &  wire908  &  _35046 ) ;
 assign _37497 = ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  wire905 ) ;
 assign _37499 = ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  wire900 ) ;
 assign _37508 = ( n_n3772 ) | ( wire395 ) | ( _5462 ) | ( _36244 ) ;
 assign _37509 = ( wire900  &  _35163 ) | ( wire906  &  _35186 ) ;
 assign _37511 = ( wire912  &  _34544 ) | ( wire900  &  _35167 ) ;
 assign _37516 = ( i_14_  &  (~ i_13_)  &  i_12_  &  wire897 ) | ( i_14_  &  i_13_  &  (~ i_12_)  &  wire897 ) | ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire897 ) ;
 assign _37517 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire903 ) | ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  wire903 ) ;
 assign _37520 = ( wire814 ) | ( n_n3768 ) | ( _4031 ) | ( _4032 ) ;
 assign _37521 = ( wire4319 ) | ( _4039 ) | ( _4040 ) | ( _4041 ) ;
 assign _37522 = ( n_n2860 ) | ( wire20562 ) | ( _37508 ) | ( _37520 ) ;
 assign _37523 = ( _37463 ) | ( _37464 ) | ( _37521 ) | ( _37522 ) ;
 assign _37525 = ( i_14_  &  i_13_  &  (~ i_12_)  &  wire904 ) | ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire904 ) ;
 assign _37527 = ( n_n4  &  wire71 ) | ( n_n4  &  wire904  &  _35153 ) ;
 assign _37530 = ( wire906  &  _35091 ) | ( wire913  &  _35748 ) ;
 assign _37532 = ( wire914  &  _34565 ) | ( wire912  &  _36184 ) ;
 assign _37535 = ( wire897  &  _35039 ) | ( wire911  &  _36168 ) ;
 assign _37539 = ( n_n265  &  wire200 ) | ( n_n265  &  wire112 ) | ( n_n265  &  wire277 ) ;
 assign _37544 = ( wire20608 ) | ( wire20609 ) | ( _4028 ) | ( _37527 ) ;
 assign _37546 = ( wire907  &  _36115 ) | ( wire914  &  _36202 ) ;
 assign _37548 = ( wire914  &  _34952 ) | ( wire900  &  _35167 ) ;
 assign _37550 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire907 ) | ( i_14_  &  i_13_  &  (~ i_12_)  &  wire907 ) ;
 assign _37552 = ( wire912  &  _34544 ) | ( wire906  &  _35186 ) ;
 assign _37560 = ( n_n4  &  wire52 ) | ( wire911  &  n_n4  &  _34580 ) ;
 assign _37562 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire913 ) | ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  wire913 ) ;
 assign _37565 = ( wire4302 ) | ( wire905  &  n_n4  &  n_n256 ) ;
 assign _37568 = ( i_14_  &  i_13_  &  (~ i_12_)  &  wire908 ) | ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire908 ) ;
 assign _37570 = ( n_n4  &  wire902  &  _35420 ) | ( n_n4  &  wire902  &  _35422 ) ;
 assign _37576 = ( wire640 ) | ( wire792 ) | ( _3973 ) | ( _37570 ) ;
 assign _37580 = ( i_14_  &  (~ i_13_)  &  i_12_  &  wire905 ) ;
 assign _37619 = ( i_5_  &  (~ i_3_)  &  (~ i_4_) ) ;
 assign _37630 = ( wire20633 ) | ( wire20642 ) | ( wire20643 ) | ( _3920 ) ;
 assign _37633 = ( n_n4508 ) | ( wire20648 ) | ( wire20629 ) | ( wire20630 ) ;
 assign _37639 = ( n_n4186 ) | ( wire20658 ) | ( wire559 ) | ( _3896 ) ;
 assign _37643 = ( wire20662 ) | ( wire19260 ) | ( wire19261 ) | ( wire19263 ) ;
 assign _37645 = ( wire926 ) | ( n_n116  &  n_n284  &  _36563 ) ;
 assign _37646 = ( i_7_  &  i_6_  &  n_n264  &  n_n116 ) | ( (~ i_7_)  &  i_6_  &  n_n264  &  n_n116 ) | ( i_7_  &  (~ i_6_)  &  n_n264  &  n_n116 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n264  &  n_n116 ) ;
 assign _37648 = ( wire879 ) | ( wire20665 ) | ( wire19996 ) | ( wire19997 ) ;
 assign _37657 = ( n_n5797 ) | ( wire20667 ) | ( wire20671 ) ;
 assign _37661 = ( n_n56  &  wire42 ) | ( n_n56  &  wire899  &  _34575 ) ;
 assign _37666 = ( wire705 ) | ( wire5552 ) | ( _4771 ) | ( _4775 ) ;
 assign _37673 = ( n_n57  &  wire166 ) | ( n_n56  &  wire166 ) ;
 assign _37686 = ( n_n285  &  n_n266  &  n_n230 ) ;
 assign _37688 = ( n_n285  &  n_n266  &  n_n230 ) ;
 assign _37689 = ( wire165  &  _37686 ) | ( wire198  &  _37688 ) ;
 assign _37701 = ( wire760 ) | ( wire20737 ) | ( wire20739 ) | ( _3852 ) ;
 assign _37703 = ( n_n4219 ) | ( wire20718 ) | ( wire20742 ) | ( _37701 ) ;
 assign _37710 = ( wire5099 ) | ( wire19862 ) | ( _3833 ) | ( _3834 ) ;
 assign _37712 = ( wire19753 ) | ( wire19754 ) | ( wire20689 ) | ( _37710 ) ;
 assign _37716 = ( wire19742 ) | ( wire19747 ) | ( _36149 ) | ( _36165 ) ;
 assign _37722 = ( wire5033 ) | ( wire708 ) | ( wire4196 ) | ( _36952 ) ;
 assign _37733 = ( wire19758 ) | ( wire20748 ) | ( _37712 ) | ( _37716 ) ;
 assign _37738 = ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  wire913 ) ;
 assign _37743 = ( i_14_  &  i_13_  &  i_12_ ) ;
 assign _37750 = ( wire392 ) | ( wire386 ) ;
 assign _37751 = ( wire19582 ) | ( wire20769 ) | ( _35709 ) | ( _37750 ) ;
 assign _37753 = ( wire899  &  _37042 ) | ( wire905  &  _37046 ) ;
 assign _37755 = ( wire911  &  _36807 ) | ( wire913  &  _36810 ) ;
 assign _37762 = ( wire44  &  n_n94 ) | ( wire904  &  n_n94  &  _35391 ) ;
 assign _37764 = ( n_n4682 ) | ( n_n4685 ) | ( wire20776 ) | ( _37762 ) ;
 assign _37766 = ( n_n260  &  n_n285  &  n_n263 ) ;
 assign _37772 = ( wire20775 ) | ( _3786 ) | ( _3787 ) ;
 assign _37776 = ( wire788 ) | ( n_n4680 ) | ( n_n4677 ) | ( wire20784 ) ;
 assign _37777 = ( wire19936 ) | ( wire19534 ) | ( _36404 ) | ( _37776 ) ;
 assign _37791 = ( wire662 ) | ( wire5564 ) | ( wire5565 ) | ( _6443 ) ;
 assign _37792 = ( n_n3843 ) | ( wire5569 ) | ( _35176 ) | ( _37791 ) ;
 assign _37796 = ( n_n5  &  wire123 ) | ( n_n5  &  wire227 ) ;
 assign _37825 = ( n_n4770 ) | ( n_n6  &  wire20839 ) | ( n_n6  &  wire20840 ) ;
 assign _37826 = ( wire4042 ) | ( _37796 ) | ( n_n5  &  wire1619 ) ;
 assign _37827 = ( wire20842 ) | ( _35257 ) | ( _35258 ) | ( _37825 ) ;
 assign _37828 = ( wire911  &  _34580 ) | ( wire913  &  _36156 ) ;
 assign _37830 = ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  wire913 ) | ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire913 ) ;
 assign _37833 = ( _3718 ) | ( _3719 ) | ( _3723 ) | ( _3724 ) ;
 assign _37834 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire899 ) | ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire899 ) ;
 assign _37840 = ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  wire905 ) ;
 assign _37841 = ( i_14_  &  (~ i_13_)  &  i_12_  &  wire905 ) ;
 assign _37846 = ( n_n3309 ) | ( n_n3579 ) | ( wire20824 ) | ( _3708 ) ;
 assign _37848 = ( wire20836 ) | ( _37792 ) | ( _37826 ) | ( _37827 ) ;
 assign _37849 = ( wire899  &  _34575 ) | ( wire913  &  _36156 ) ;
 assign _37852 = ( wire468 ) | ( wire913  &  n_n220  &  n_n2 ) ;
 assign _37859 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire904 ) | ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  wire904 ) ;
 assign _37860 = ( i_14_  &  (~ i_13_)  &  i_12_  &  wire899 ) | ( i_14_  &  i_13_  &  (~ i_12_)  &  wire899 ) | ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire899 ) ;
 assign _37862 = ( n_n3778 ) | ( n_n2633 ) | ( _3679 ) | ( _3680 ) ;
 assign _37876 = ( n_n4807 ) | ( n_n4808 ) | ( wire3989 ) ;
 assign _37878 = ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  wire911 ) ;
 assign _37898 = ( wire20881 ) | ( n_n3385 ) | ( wire20895 ) | ( _37876 ) ;
 assign _37899 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire899 ) | ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire899 ) ;
 assign _37901 = ( n_n3  &  wire79 ) | ( wire905  &  n_n3  &  _36137 ) ;
 assign _37905 = ( wire911  &  _34580 ) | ( wire913  &  _35748 ) ;
 assign _37907 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire913 ) | ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire913 ) ;
 assign _37910 = ( _3628 ) | ( _3629 ) | ( _3988 ) | ( _37560 ) ;
 assign _37915 = ( i_14_  &  (~ i_13_)  &  i_12_  &  wire905 ) ;
 assign _37919 = ( wire913  &  n_n281 ) | ( wire905  &  _36337 ) ;
 assign _37920 = ( wire75  &  n_n2 ) | ( wire911  &  n_n2  &  _36168 ) ;
 assign _37922 = ( wire911  &  _34580 ) | ( wire913  &  _35938 ) ;
 assign _37925 = ( wire4071 ) | ( wire20809 ) | ( _3602 ) | ( _37920 ) ;
 assign _37931 = ( n_n1440 ) | ( wire5758 ) | ( _6220 ) | ( _6221 ) ;
 assign _37932 = ( wire19383 ) | ( wire5775 ) ;
 assign _37934 = ( wire4073 ) | ( wire20814 ) | ( _37925 ) | ( _37931 ) ;
 assign _37936 = ( (~ i_14_)  &  i_13_  &  i_12_ ) ;
 assign _37951 = ( wire254  &  _35400 ) | ( wire1786  &  _35412 ) ;
 assign _37961 = ( (~ i_10_)  &  (~ i_9_) ) ;
 assign _37967 = ( wire3945 ) | ( wire20920 ) | ( wire758 ) | ( wire3946 ) ;
 assign _37968 = ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  wire907 ) ;
 assign _37969 = ( wire905  &  _34956 ) | ( wire913  &  _35748 ) ;
 assign _37976 = ( wire4745 ) | ( wire20131 ) | ( _4694 ) | ( _36984 ) ;
 assign _37977 = ( i_14_  &  i_13_  &  i_12_  &  wire912 ) ;
 assign _37989 = ( n_n4624 ) | ( wire21035 ) | ( n_n4633 ) | ( _3547 ) ;
 assign _37993 = ( wire3831 ) | ( wire3830 ) ;
 assign _37994 = ( n_n1555 ) | ( _3529 ) | ( _6461 ) | ( _35154 ) ;
 assign _38006 = ( (~ i_14_)  &  i_13_  &  i_12_  &  i_15_ ) ;
 assign _38007 = ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  (~ i_15_) ) ;
 assign _38010 = ( i_14_  &  (~ i_13_)  &  i_12_  &  wire912 ) ;
 assign _38014 = ( _4324 ) | ( _4514 ) | ( _37253 ) | ( _37298 ) ;
 assign _38018 = ( n_n264  &  n_n273  &  n_n285 ) ;
 assign _38020 = ( wire904  &  _35391 ) | ( wire905  &  _36137 ) ;
 assign _38025 = ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  wire908 ) ;
 assign _38049 = ( n_n260  &  n_n285  &  n_n261 ) ;
 assign _38050 = ( i_14_  &  i_13_  &  i_12_  &  wire912 ) ;
 assign _38057 = ( wire4117 ) | ( wire20772 ) | ( _4252 ) | ( _37360 ) ;
 assign _38062 = ( i_14_  &  i_13_  &  (~ i_12_)  &  (~ i_15_) ) ;
 assign _38063 = ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  (~ i_15_) ) ;
 assign _38067 = ( wire767 ) | ( wire21098 ) | ( _4226 ) | ( _37381 ) ;
 assign _38069 = ( wire80  &  n_n94 ) | ( wire902  &  n_n94  &  _35622 ) ;
 assign _38073 = ( wire459 ) | ( n_n1633 ) | ( _3449 ) | ( _38069 ) ;
 assign _38082 = ( wire21101 ) | ( wire21105 ) | ( _38067 ) | ( _38073 ) ;
 assign _38083 = ( n_n258  &  wire904 ) | ( wire898  &  _35396 ) ;
 assign _38087 = ( wire636 ) | ( wire21065 ) | ( _3423 ) | ( _3424 ) ;
 assign _38093 = ( _4177 ) | ( _4792 ) | ( _36881 ) | ( _37411 ) ;
 assign _38097 = ( n_n2  &  wire57 ) | ( n_n2  &  wire912  &  _34544 ) ;
 assign _38103 = ( n_n3257 ) | ( wire20959 ) | ( _3408 ) | ( _38097 ) ;
 assign _38106 = ( n_n3255 ) | ( wire814 ) | ( wire3884 ) | ( _3400 ) ;
 assign _38107 = ( wire496 ) | ( _5389 ) | ( _36298 ) ;
 assign _38108 = ( wire806 ) | ( wire20967 ) | ( _3396 ) ;
 assign _38109 = ( n_n2860 ) | ( _38106 ) | ( _38107 ) | ( _38108 ) ;
 assign _38118 = ( (~ i_14_)  &  i_13_  &  i_12_  &  wire898 ) | ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire898 ) ;
 assign _38123 = ( i_14_  &  i_13_  &  i_12_  &  wire912 ) ;
 assign _38125 = ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  wire908 ) ;
 assign _38131 = ( n_n260  &  n_n285  &  n_n263 ) ;
 assign _38132 = ( i_14_  &  (~ i_13_)  &  i_12_  &  wire914 ) ;
 assign _38136 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  i_15_ ) ;
 assign _38137 = ( i_14_  &  i_13_  &  (~ i_12_)  &  (~ i_15_) ) ;
 assign _38138 = ( wire908  &  _35120 ) | ( wire905  &  _36909 ) ;
 assign _38140 = ( i_14_  &  (~ i_13_)  &  i_12_  &  i_15_ ) ;
 assign _38141 = ( i_14_  &  i_13_  &  i_12_  &  (~ i_15_) ) ;
 assign _38142 = ( wire88  &  n_n227 ) | ( n_n227  &  wire306 ) ;
 assign _38151 = ( wire4694 ) | ( wire4695 ) | ( _4149 ) | ( _37432 ) ;
 assign _38155 = ( wire914  &  _34952 ) | ( wire908  &  _35212 ) ;
 assign _38156 = ( (~ i_14_)  &  i_13_  &  i_12_  &  wire902 ) | ( i_14_  &  (~ i_13_)  &  i_12_  &  wire902 ) | ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire902 ) | ( i_14_  &  i_13_  &  (~ i_12_)  &  wire902 ) ;
 assign _38157 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire908 ) | ( i_14_  &  i_13_  &  (~ i_12_)  &  wire908 ) ;
 assign _38161 = ( (~ i_14_)  &  i_13_  &  i_12_  &  wire912 ) ;
 assign _38164 = ( n_n111  &  n_n4 ) | ( n_n4  &  wire57 ) | ( n_n4  &  _3333 ) ;
 assign _38165 = ( wire557 ) | ( n_n4  &  wire245 ) | ( n_n4  &  _38161 ) ;
 assign _38167 = ( wire905  &  _36137 ) | ( wire899  &  _36255 ) ;
 assign _38169 = ( i_14_  &  (~ i_13_)  &  i_12_  &  wire899 ) | ( i_14_  &  i_13_  &  (~ i_12_)  &  wire899 ) | ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire899 ) ;
 assign _38171 = ( n_n208  &  n_n284  &  n_n285 ) ;
 assign _38174 = ( wire4302 ) | ( wire905  &  n_n4  &  n_n256 ) ;
 assign _38178 = ( n_n2  &  wire63 ) | ( n_n2  &  wire902  &  _35056 ) ;
 assign _38183 = ( _3311 ) | ( _5302 ) | ( _5303 ) | ( _38178 ) ;
 assign _38186 = ( wire20933 ) | ( wire20934 ) | ( _4028 ) | ( _37527 ) ;
 assign _38187 = ( wire904  &  _35391 ) | ( wire898  &  _35396 ) ;
 assign _38189 = ( wire914  &  _34565 ) | ( wire912  &  _36184 ) ;
 assign _38192 = ( wire20938 ) | ( n_n3519 ) | ( n_n3520 ) | ( _3296 ) ;
 assign _38195 = ( i_14_  &  (~ i_13_)  &  i_12_  &  wire905 ) ;
 assign _38196 = ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  wire908 ) ;
 assign _38202 = ( wire20936 ) | ( wire20942 ) | ( _38186 ) | ( _38192 ) ;
 assign _38208 = ( wire913  &  n_n220 ) | ( n_n220  &  wire914 ) ;
 assign _38211 = ( wire914  &  _34952 ) | ( wire913  &  _35748 ) ;
 assign _38238 = ( wire3726 ) | ( wire3725 ) ;
 assign _38244 = ( wire21178 ) | ( wire3720 ) | ( wire21168 ) | ( _3260 ) ;
 assign _38245 = ( wire21163 ) | ( wire21173 ) | ( _38238 ) | ( _38244 ) ;
 assign _38248 = ( n_n247  &  _36683 ) | ( n_n247  &  _37013 ) | ( n_n247  &  _37014 ) ;
 assign _38249 = ( (~ i_14_)  &  i_13_  &  i_12_  &  wire914 ) | ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire914 ) ;
 assign _38251 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire902 ) ;
 assign _38254 = ( n_n884 ) | ( n_n4  &  wire80 ) | ( n_n4  &  _38251 ) ;
 assign _38256 = ( (~ i_14_)  &  i_13_  &  i_12_  &  wire901 ) | ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire901 ) ;
 assign _38258 = ( i_14_  &  (~ i_13_)  &  i_12_  &  wire901 ) | ( i_14_  &  i_13_  &  (~ i_12_)  &  wire901 ) ;
 assign _38260 = ( (~ i_14_)  &  i_13_  &  i_12_  &  wire914 ) | ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire914 ) | ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  wire914 ) ;
 assign _38262 = ( i_14_  &  i_13_  &  (~ i_12_)  &  wire906 ) ;
 assign _38263 = ( i_14_  &  (~ i_13_)  &  i_12_  &  wire912 ) ;
 assign _38266 = ( wire914  &  _36382 ) | ( n_n247  &  _36683 ) ;
 assign _38268 = ( wire4470 ) | ( n_n4  &  wire19578 ) | ( n_n4  &  _38262 ) ;
 assign _38272 = ( n_n4  &  wire469 ) | ( n_n4  &  wire899  &  _37042 ) ;
 assign _38273 = ( i_14_  &  (~ i_13_)  &  i_12_  &  wire902 ) | ( i_14_  &  i_13_  &  (~ i_12_)  &  wire902 ) ;
 assign _38274 = ( wire897  &  _35539 ) | ( wire903  &  _35628 ) ;
 assign _38277 = ( wire902  &  _35622 ) | ( n_n222  &  _36699 ) ;
 assign _38285 = ( wire911  &  _36343 ) | ( wire913  &  _36810 ) ;
 assign _38287 = ( n_n222  &  _36699 ) | ( wire911  &  _36807 ) ;
 assign _38289 = ( wire913  &  _36810 ) | ( wire905  &  _37046 ) ;
 assign _38291 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire899 ) | ( i_14_  &  i_13_  &  (~ i_12_)  &  wire899 ) ;
 assign _38294 = ( wire519 ) | ( _3180 ) | ( _3181 ) | ( _3182 ) ;
 assign _38296 = ( i_14_  &  (~ i_13_)  &  i_12_  &  wire905 ) ;
 assign _38299 = ( i_14_  &  i_13_  &  i_12_  &  wire901 ) ;
 assign _38302 = ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  wire906 ) ;
 assign _38305 = ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  wire904 ) ;
 assign _38311 = ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  wire908 ) ;
 assign _38313 = ( i_14_  &  i_13_  &  i_12_  &  wire902 ) ;
 assign _38315 = ( n_n4  &  wire113 ) | ( wire907  &  n_n4  &  _36833 ) ;
 assign _38317 = ( n_n4005 ) | ( wire3642 ) | ( wire21238 ) | ( _38315 ) ;
 assign _38319 = ( n_n3930 ) | ( n_n3929 ) | ( n_n3406 ) | ( _38317 ) ;
 assign _38320 = ( wire21220 ) | ( wire3680 ) | ( wire3681 ) | ( _38294 ) ;
 assign _38323 = ( n_n4  &  wire42 ) | ( n_n4  &  wire899  &  _34575 ) ;
 assign _38325 = ( wire21180 ) | ( _3973 ) | ( _37570 ) | ( _38323 ) ;
 assign _38328 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire897 ) | ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire897 ) ;
 assign _38330 = ( n_n268  &  wire19408 ) | ( n_n268  &  wire903  &  _35109 ) ;
 assign _38335 = ( i_14_  &  i_13_  &  i_12_  &  wire902 ) ;
 assign _38339 = ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  wire908 ) ;
 assign _38343 = ( n_n1440 ) | ( wire5758 ) | ( _6220 ) | ( _6221 ) ;
 assign _38345 = ( wire911  &  _34580 ) | ( wire913  &  _35938 ) ;
 assign _38348 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire907 ) | ( i_14_  &  i_13_  &  (~ i_12_)  &  wire907 ) ;
 assign _38354 = ( n_n1370 ) | ( wire21281 ) | ( _3106 ) | ( _3107 ) ;
 assign _38355 = ( wire912  &  _34544 ) | ( wire911  &  _36168 ) ;
 assign _38357 = ( wire912  &  _36095 ) | ( wire914  &  _36202 ) ;
 assign _38361 = ( n_n284  &  n_n285  &  n_n266 ) ;
 assign _38365 = ( (~ i_14_)  &  i_13_  &  i_12_  &  wire898 ) | ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire898 ) ;
 assign _38367 = ( n_n4  &  wire96 ) | ( n_n4  &  wire898  &  _35693 ) ;
 assign _38368 = ( i_14_  &  i_13_  &  i_12_  &  wire906 ) | ( (~ i_14_)  &  i_13_  &  i_12_  &  wire906 ) ;
 assign _38369 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire900 ) | ( i_14_  &  i_13_  &  (~ i_12_)  &  wire900 ) | ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire900 ) | ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  wire900 ) ;
 assign _38370 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire906 ) | ( i_14_  &  i_13_  &  (~ i_12_)  &  wire906 ) | ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  wire906 ) ;
 assign _38371 = ( n_n4  &  n_n105 ) | ( n_n105  &  n_n3 ) | ( n_n4  &  wire77 ) ;
 assign _38372 = ( _3077 ) | ( _3078 ) | ( _3082 ) | ( _38367 ) ;
 assign _38374 = ( wire3626 ) | ( wire21276 ) | ( wire21288 ) | ( _38372 ) ;
 assign _38379 = ( n_n57  &  n_n99 ) | ( n_n57  &  wire19575 ) | ( n_n57  &  _3070 ) ;
 assign _38380 = ( n_n258  &  wire900 ) | ( wire906  &  _35705 ) ;
 assign _38381 = ( n_n56  &  wire19577 ) | ( n_n56  &  wire906  &  _35716 ) ;
 assign _38386 = ( wire21298 ) | ( wire21299 ) | ( _3058 ) | ( _38381 ) ;
 assign _38390 = ( (~ i_14_)  &  i_13_  &  i_12_  &  wire901 ) | ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire901 ) ;
 assign _38392 = ( i_14_  &  (~ i_13_)  &  i_12_  &  wire901 ) | ( i_14_  &  i_13_  &  (~ i_12_)  &  wire901 ) ;
 assign _38394 = ( n_n247  &  _36683 ) | ( n_n247  &  _37013 ) | ( n_n247  &  _37014 ) ;
 assign _38395 = ( (~ i_14_)  &  i_13_  &  i_12_  &  wire914 ) | ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire914 ) ;
 assign _38398 = ( wire497 ) | ( n_n1597 ) | ( _3043 ) | ( _3044 ) ;
 assign _38399 = ( wire906  &  _35685 ) | ( wire898  &  _35695 ) ;
 assign _38403 = ( i_14_  &  i_13_  &  i_12_  &  wire906 ) | ( (~ i_14_)  &  i_13_  &  i_12_  &  wire906 ) ;
 assign _38404 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire900 ) | ( i_14_  &  i_13_  &  (~ i_12_)  &  wire900 ) | ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire900 ) | ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  wire900 ) ;
 assign _38405 = ( n_n258  &  wire900 ) | ( wire906  &  _35705 ) ;
 assign _38408 = ( wire3595 ) | ( wire3588 ) | ( wire21318 ) | ( _38398 ) ;
 assign _38409 = ( wire897  &  _35539 ) | ( wire902  &  _35622 ) ;
 assign _38411 = ( wire902  &  n_n225 ) | ( wire897  &  _35544 ) ;
 assign _38413 = ( (~ i_14_)  &  i_13_  &  i_12_  &  wire903 ) | ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire903 ) ;
 assign _38418 = ( n_n247  &  _36683 ) | ( n_n247  &  _37013 ) | ( n_n247  &  _37014 ) ;
 assign _38419 = ( (~ i_14_)  &  i_13_  &  i_12_  &  wire914 ) | ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire914 ) ;
 assign _38421 = ( (~ i_14_)  &  i_13_  &  i_12_  &  wire901 ) | ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire901 ) ;
 assign _38423 = ( wire902  &  _35420 ) | ( wire901  &  _36790 ) ;
 assign _38426 = ( wire903  &  _35628 ) | ( wire899  &  _37042 ) ;
 assign _38430 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire902 ) | ( i_14_  &  i_13_  &  (~ i_12_)  &  wire902 ) ;
 assign _38432 = ( (~ i_14_)  &  i_13_  &  i_12_  &  wire902 ) | ( i_14_  &  (~ i_13_)  &  i_12_  &  wire902 ) ;
 assign _38436 = ( n_n1591 ) | ( wire3558 ) | ( _3013 ) | ( _3014 ) ;
 assign _38437 = ( wire911  &  _36807 ) | ( wire913  &  _36810 ) ;
 assign _38439 = ( wire911  &  n_n258 ) | ( n_n222  &  _36699 ) ;
 assign _38442 = ( wire589 ) | ( wire481 ) | ( _2982 ) | ( _2983 ) ;
 assign _38444 = ( n_n56  &  wire113 ) | ( wire914  &  n_n56  &  _34565 ) ;
 assign _38448 = ( wire901  &  _36817 ) | ( wire907  &  _36833 ) ;
 assign _38451 = ( wire21329 ) | ( _2965 ) | ( _2976 ) | ( _38444 ) ;
 assign _38452 = ( wire900  &  _35074 ) | ( wire899  &  _37042 ) ;
 assign _38462 = ( wire3578 ) | ( wire3551 ) | ( wire21356 ) | ( _38442 ) ;
 assign _38467 = ( wire3544 ) | ( _2946 ) | ( n_n56  &  wire955 ) ;
 assign _38468 = ( n_n2440 ) | ( n_n2439 ) | ( _38408 ) | ( _38467 ) ;
 assign _38469 = ( n_n2431 ) | ( wire21352 ) | ( _38436 ) | ( _38462 ) ;
 assign _38483 = ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  (~ i_15_) ) ;
 assign _38485 = ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  i_15_ ) ;
 assign _38513 = ( n_n56  &  wire86 ) | ( wire907  &  n_n56  &  _36210 ) ;
 assign _38522 = ( wire21467 ) | ( wire21466 ) ;
 assign _38545 = ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire898 ) ;
 assign _38550 = ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire900 ) | ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  wire900 ) ;
 assign _38551 = ( (~ i_14_)  &  i_13_  &  i_12_  &  wire906 ) | ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire906 ) | ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  wire906 ) | ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire906 ) ;
 assign _38556 = ( (~ i_9_)  &  i_10_  &  (~ i_11_)  &  (~ i_15_) ) ;
 assign _38558 = ( (~ i_9_)  &  i_10_  &  (~ i_11_)  &  i_15_ ) ;
 assign _38613 = ( n_n94  &  wire167 ) | ( n_n94  &  wire119 ) ;
 assign _38614 = ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  wire911 ) ;
 assign _38625 = ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  wire901 ) ;
 assign _38635 = ( wire21479 ) | ( _2793 ) | ( _38613 ) ;
 assign _38636 = ( n_n2097 ) | ( n_n2180 ) | ( wire3375 ) | ( wire3376 ) ;
 assign _38637 = ( wire21508 ) | ( wire21505 ) | ( wire21506 ) ;
 assign _38639 = ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  wire907 ) ;
 assign _38640 = ( wire903  &  _35190 ) | ( wire914  &  _36202 ) ;
 assign _38643 = ( wire903  &  _35109 ) | ( wire913  &  _36156 ) ;
 assign _38656 = ( wire904  &  _35139 ) | ( wire914  &  _36977 ) ;
 assign _38658 = ( n_n4  &  wire77 ) | ( n_n4  &  wire912  &  _34544 ) ;
 assign _38663 = ( wire907  &  _36115 ) | ( wire901  &  _36788 ) ;
 assign _38665 = ( n_n279  &  wire912 ) | ( wire914  &  _36977 ) ;
 assign _38666 = ( n_n279  &  wire900 ) | ( n_n279  &  wire904 ) ;
 assign _38668 = ( _2727 ) | ( _2728 ) | ( _2732 ) | ( _2733 ) ;
 assign _38670 = ( n_n2108 ) | ( _2741 ) | ( _38658 ) ;
 assign _38673 = ( n_n2  &  wire157 ) | ( n_n2  &  wire330 ) ;
 assign _38679 = ( n_n260  &  n_n285  &  n_n283 ) ;
 assign _38681 = ( n_n1  &  wire399 ) | ( n_n1  &  wire338 ) ;
 assign _38691 = ( _2711 ) | ( _38681 ) | ( wire1097  &  _38679 ) ;
 assign _38699 = ( wire911  &  _34580 ) | ( wire913  &  _36810 ) ;
 assign _38703 = ( n_n229  &  n_n284  &  n_n285 ) ;
 assign _38708 = ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  wire907 ) ;
 assign _38713 = ( wire1450  &  _38703 ) | ( wire169  &  _38708 ) ;
 assign _38722 = ( wire902  &  _35418 ) | ( wire897  &  _35661 ) ;
 assign _38723 = ( (~ i_14_)  &  i_13_  &  i_12_  &  wire903 ) | ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire903 ) | ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  wire903 ) | ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire903 ) ;
 assign _38724 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire908 ) | ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  wire908 ) | ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire908 ) ;
 assign _38725 = ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire899 ) ;
 assign _38726 = ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire897 ) | ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  wire897 ) ;
 assign _38727 = ( (~ i_14_)  &  i_13_  &  i_12_  &  wire903 ) | ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire903 ) | ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  wire903 ) | ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire903 ) ;
 assign _38729 = ( wire21614 ) | ( _2656 ) | ( _2657 ) ;
 assign _38730 = ( wire333 ) | ( wire3541 ) | ( wire3542 ) | ( wire21372 ) ;
 assign _38732 = ( n_n2099 ) | ( wire3368 ) | ( wire21525 ) | ( _2677 ) ;
 assign _38733 = ( wire21408 ) | ( wire21409 ) | ( wire21415 ) | ( _38691 ) ;
 assign _38734 = ( _38729 ) | ( _38730 ) | ( _38732 ) | ( _38733 ) ;
 assign _38740 = ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  wire908 ) ;
 assign _38741 = ( wire908  &  _35212 ) | ( wire905  &  _36909 ) ;
 assign _38748 = ( n_n260  &  n_n273  &  n_n285 ) ;
 assign _38750 = ( n_n2  &  wire241 ) | ( n_n2  &  wire242 ) ;
 assign _38769 = ( _2630 ) | ( _38750 ) | ( wire1159  &  _38748 ) ;
 assign _38770 = ( n_n2129 ) | ( wire21431 ) | ( wire21432 ) | ( _38769 ) ;
 assign _38772 = ( wire911  &  _34580 ) | ( wire913  &  _36810 ) ;
 assign _38785 = ( wire21529 ) | ( wire3354 ) ;
 assign _38788 = ( (~ i_14_)  &  i_13_  &  i_12_  &  (~ i_15_) ) ;
 assign _38789 = ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  i_15_ ) ;
 assign _38794 = ( n_n260  &  n_n285  &  n_n263 ) ;
 assign _38804 = ( wire902  &  _35418 ) | ( wire897  &  _35661 ) ;
 assign _38805 = ( (~ i_14_)  &  i_13_  &  i_12_  &  wire903 ) | ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire903 ) | ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  wire903 ) | ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire903 ) ;
 assign _38806 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire908 ) | ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  wire908 ) | ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire908 ) ;
 assign _38809 = ( _2557 ) | ( _2558 ) | ( n_n6  &  wire1486 ) ;
 assign _38844 = ( wire907  &  _36115 ) | ( wire914  &  _36977 ) ;
 assign _38846 = ( n_n5  &  wire78 ) | ( n_n5  &  wire21576 ) ;
 assign _38848 = ( wire21579 ) | ( wire3287 ) ;
 assign _38853 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire904 ) | ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  wire904 ) | ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire904 ) ;
 assign _38854 = ( n_n5  &  wire51 ) | ( n_n5  &  wire898  &  _36030 ) ;
 assign _38855 = ( wire900  &  _35167 ) | ( wire914  &  _36977 ) ;
 assign _38857 = ( n_n6  &  wire51 ) | ( n_n6  &  wire21584 ) ;
 assign _38858 = ( _2498 ) | ( _2503 ) | ( _38854 ) | ( _38857 ) ;
 assign _38860 = ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  (~ i_15_) ) ;
 assign _38862 = ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  i_15_ ) ;
 assign _38867 = ( wire907  &  _36115 ) | ( wire901  &  _36788 ) ;
 assign _38870 = ( (~ i_14_)  &  i_13_  &  i_12_  &  wire914 ) | ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire914 ) | ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  wire914 ) ;
 assign _38872 = ( _2483 ) | ( _2486 ) | ( _2487 ) ;
 assign _38874 = ( wire904  &  _35427 ) | ( wire905  &  _36909 ) ;
 assign _38877 = ( wire911  &  _34580 ) | ( wire913  &  _36810 ) ;
 assign _38880 = ( n_n53  &  n_n19 ) | ( wire899  &  n_n53  &  _35752 ) ;
 assign _38881 = ( wire456 ) | ( wire21603 ) | ( _2478 ) | ( _38880 ) ;
 assign _38882 = ( _2474 ) | ( _2475 ) | ( _2476 ) | ( _2477 ) ;
 assign _38883 = ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  (~ i_15_) ) ;
 assign _38885 = ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  i_15_ ) ;
 assign _38891 = ( n_n264  &  n_n285  &  n_n283 ) ;
 assign _38892 = ( n_n279  &  wire902 ) | ( n_n279  &  wire908 ) ;
 assign _38897 = ( n_n264  &  n_n273  &  n_n285 ) ;
 assign _38898 = ( wire69  &  _38891 ) | ( wire1528  &  _38897 ) ;
 assign _38900 = ( n_n2155 ) | ( _38872 ) | ( _38881 ) | ( _38882 ) ;
 assign _38902 = ( wire21440 ) | ( wire21612 ) | ( _38770 ) | ( _38900 ) ;
 assign _38906 = ( n_n165  &  n_n273  &  n_n284 ) ;
 assign _38907 = ( (~ i_9_)  &  (~ i_10_) ) | ( wire905  &  _34956 ) ;
 assign _38930 = ( wire21627 ) | ( wire21626 ) ;
 assign _38932 = ( n_n1670 ) | ( wire3232 ) | ( wire21628 ) | ( _38930 ) ;
 assign _38941 = ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  (~ i_15_) ) ;
 assign _38942 = ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  i_15_ ) ;
 assign _38943 = ( wire904  &  _35141 ) | ( wire898  &  _35693 ) ;
 assign _38945 = ( wire21660 ) | ( wire3198 ) ;
 assign _38957 = ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  (~ i_15_) ) ;
 assign _38958 = ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  i_15_ ) ;
 assign _38965 = ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  (~ i_15_) ) ;
 assign _38966 = ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  i_15_ ) ;
 assign _38968 = ( n_n208  &  n_n284  &  n_n285 ) ;
 assign _38969 = ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  wire904 ) ;
 assign _38971 = ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_) ) ;
 assign _38972 = ( (~ i_14_)  &  i_13_  &  i_12_  &  i_15_ ) ;
 assign _38973 = ( i_14_  &  i_13_  &  (~ i_12_)  &  (~ i_15_) ) ;
 assign _38978 = ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  (~ i_15_) ) ;
 assign _38979 = ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  i_15_ ) ;
 assign _38984 = ( wire21657 ) | ( wire21652 ) | ( _2403 ) | ( _2404 ) ;
 assign _38986 = ( wire914  &  _34952 ) | ( wire903  &  _35101 ) ;
 assign _39001 = ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  (~ i_15_) ) ;
 assign _39002 = ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  i_15_ ) ;
 assign _39005 = ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  (~ i_15_) ) ;
 assign _39006 = ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  i_15_ ) ;
 assign _39007 = ( wire903  &  _35101 ) | ( wire901  &  _36986 ) ;
 assign _39009 = ( _2337 ) | ( _2346 ) | ( _2347 ) | ( _2348 ) ;
 assign _39010 = ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  (~ i_15_) ) ;
 assign _39011 = ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  i_15_ ) ;
 assign _39044 = ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_) ) ;
 assign _39048 = ( wire900  &  _35163 ) | ( wire899  &  _37936 ) ;
 assign _39051 = ( n_n208  &  n_n284  &  n_n285 ) ;
 assign _39052 = ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  wire905 ) ;
 assign _39053 = ( i_14_  &  i_13_  &  (~ i_12_)  &  wire900 ) ;
 assign _39055 = ( wire3186 ) | ( wire3159 ) | ( n_n4  &  wire270 ) ;
 assign _39057 = ( i_14_  &  i_13_  &  (~ i_12_)  &  (~ i_15_) ) ;
 assign _39059 = ( i_14_  &  i_13_  &  (~ i_12_)  &  i_15_ ) ;
 assign _39063 = ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  wire913 ) ;
 assign _39067 = ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  wire908 ) ;
 assign _39072 = ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  (~ i_15_) ) ;
 assign _39073 = ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  i_15_ ) ;
 assign _39078 = ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  wire901 ) ;
 assign _39081 = ( i_14_  &  i_13_  &  (~ i_12_)  &  wire899 ) ;
 assign _39084 = ( (~ i_14_)  &  i_13_  &  i_12_  &  i_15_ ) ;
 assign _39085 = ( i_14_  &  i_13_  &  (~ i_12_)  &  (~ i_15_) ) ;
 assign _39091 = ( wire3120 ) | ( n_n220  &  n_n2  &  wire901 ) ;
 assign _39094 = ( n_n1697 ) | ( wire21673 ) | ( wire21648 ) | ( _38984 ) ;
 assign _39095 = ( n_n1703 ) | ( n_n1704 ) | ( wire21649 ) | ( wire21709 ) ;
 assign _39096 = ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  wire899 ) ;
 assign _39097 = ( wire904  &  _35141 ) | ( wire898  &  _35693 ) ;
 assign _39100 = ( wire900  &  _35163 ) | ( wire898  &  _35693 ) ;
 assign _39109 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire897 ) | ( i_14_  &  i_13_  &  (~ i_12_)  &  wire897 ) ;
 assign _39113 = ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  wire905 ) ;
 assign _39114 = ( (~ i_14_)  &  i_13_  &  i_12_  &  i_15_ ) ;
 assign _39115 = ( i_14_  &  i_13_  &  (~ i_12_)  &  (~ i_15_) ) ;
 assign _39118 = ( wire2961 ) | ( wire2960 ) ;
 assign _39122 = ( n_n264  &  n_n285  &  n_n283 ) ;
 assign _39131 = ( n_n264  &  n_n285  &  n_n283 ) ;
 assign _39255 = ( (~ i_9_)  &  i_10_  &  (~ i_11_)  &  (~ i_15_) ) ;
 assign _39273 = ( n_n220  &  wire898 ) | ( n_n222  &  _36699 ) ;
 assign _39274 = ( n_n53  &  wire84 ) | ( n_n222  &  n_n53  &  _39255 ) ;
 assign _39275 = ( (~ i_14_)  &  i_13_  &  i_12_  &  wire899 ) | ( i_14_  &  i_13_  &  (~ i_12_)  &  wire899 ) ;
 assign _39283 = ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  wire901 ) ;
 assign _39286 = ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  wire914 ) ;
 assign _39296 = ( wire900  &  _35163 ) | ( wire898  &  _35693 ) ;
 assign _39307 = ( n_n1774 ) | ( wire3032 ) | ( wire3033 ) | ( wire21799 ) ;
 assign _39309 = ( n_n5  &  wire195 ) | ( n_n5  &  n_n222  &  _36699 ) ;
 assign _39322 = ( (~ i_14_)  &  i_13_  &  i_12_  &  wire899 ) | ( i_14_  &  i_13_  &  (~ i_12_)  &  wire899 ) ;
 assign _39332 = ( wire21813 ) | ( wire21814 ) | ( wire2994 ) | ( _1934 ) ;
 assign _39334 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire897 ) | ( i_14_  &  i_13_  &  (~ i_12_)  &  wire897 ) ;
 assign _39337 = ( n_n5  &  wire154 ) | ( n_n5  &  n_n247  &  _36683 ) ;
 assign _39338 = ( wire908  &  _35071 ) | ( wire907  &  _36107 ) ;
 assign _39340 = ( n_n6  &  wire154 ) | ( n_n6  &  wire21821 ) ;
 assign _39341 = ( wire3005 ) | ( _1898 ) | ( _1909 ) | ( _39340 ) ;
 assign _39346 = ( n_n1689 ) | ( n_n1692 ) | ( _39094 ) | ( _39095 ) ;
 assign _39347 = ( (~ i_9_)  &  i_10_  &  (~ i_11_)  &  (~ i_15_) ) ;
 assign _39348 = ( (~ i_9_)  &  i_10_  &  (~ i_11_)  &  i_15_ ) ;
 assign _39350 = ( n_n4  &  wire143 ) | ( n_n4  &  wire899  &  _37936 ) ;
 assign _39351 = ( n_n3  &  wire195 ) | ( n_n3  &  wire230 ) ;
 assign _39356 = ( _1889 ) | ( _1892 ) | ( _39350 ) | ( _39351 ) ;
 assign _39359 = ( n_n229  &  n_n284  &  n_n285 ) ;
 assign _39360 = ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  wire901 ) ;
 assign _39363 = ( wire1668  &  _39359 ) | ( wire169  &  _39360 ) ;
 assign _39369 = ( (~ i_14_)  &  i_13_  &  i_12_  &  wire899 ) | ( i_14_  &  i_13_  &  (~ i_12_)  &  wire899 ) | ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  wire899 ) ;
 assign _39370 = ( n_n3  &  wire375 ) | ( wire902  &  n_n3  &  _35049 ) ;
 assign _39372 = ( wire21896 ) | ( n_n4  &  wire195 ) | ( n_n4  &  wire21892 ) ;
 assign _39375 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire897 ) | ( i_14_  &  i_13_  &  (~ i_12_)  &  wire897 ) ;
 assign _39379 = ( wire907  &  _36107 ) | ( wire901  &  _36790 ) ;
 assign _39382 = ( wire21635 ) | ( wire2893 ) | ( _1843 ) | ( _1853 ) ;
 assign _39384 = ( wire21904 ) | ( wire590 ) | ( wire19306 ) | ( _34942 ) ;
 assign _39387 = ( n_n268  &  wire95 ) | ( n_n268  &  wire22001 ) ;
 assign _39389 = ( wire22000 ) | ( n_n4  &  wire99 ) | ( n_n4  &  wire41 ) ;
 assign _39396 = ( wire913  &  _35938 ) | ( wire911  &  _36330 ) ;
 assign _39398 = ( wire907  &  _36783 ) | ( wire901  &  _36988 ) ;
 assign _39406 = ( n_n229  &  n_n284  &  n_n285 ) ;
 assign _39412 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire900 ) | ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  wire900 ) ;
 assign _39425 = ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  wire899 ) ;
 assign _39426 = ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  i_15_ ) ;
 assign _39427 = ( i_14_  &  (~ i_13_)  &  i_12_  &  (~ i_15_) ) ;
 assign _39432 = ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  wire898 ) ;
 assign _39441 = ( wire913  &  _35938 ) | ( wire911  &  _36330 ) ;
 assign _39449 = ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  wire908 ) ;
 assign _39450 = ( n_n3  &  _39449 ) | ( wire911  &  n_n258  &  n_n3 ) ;
 assign _39461 = ( (~ i_14_)  &  i_13_  &  i_12_  &  wire912 ) | ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  wire912 ) ;
 assign _39470 = ( i_14_  &  i_13_  &  i_12_ ) ;
 assign _39479 = ( n_n220  &  wire907 ) | ( wire901  &  _36988 ) ;
 assign _39486 = ( _1729 ) | ( _1730 ) | ( n_n4  &  wire1492 ) ;
 assign _39495 = ( n_n3731 ) | ( n_n1339 ) | ( _1718 ) | ( _1719 ) ;
 assign _39502 = ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  wire901 ) ;
 assign _39514 = ( wire907  &  _36115 ) | ( wire901  &  _37291 ) ;
 assign _39526 = ( wire914  &  _36382 ) | ( wire907  &  _36783 ) ;
 assign _39528 = ( n_n4174 ) | ( wire516 ) | ( n_n1555 ) | ( _1683 ) ;
 assign _39529 = ( i_14_  &  i_13_  &  i_12_  &  (~ i_15_) ) ;
 assign _39530 = ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  i_15_ ) ;
 assign _39534 = ( n_n53  &  wire68 ) | ( n_n53  &  wire175 ) ;
 assign _39536 = ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  i_15_ ) ;
 assign _39537 = ( i_14_  &  (~ i_13_)  &  i_12_  &  (~ i_15_) ) ;
 assign _39540 = ( wire764 ) | ( wire579 ) ;
 assign _39542 = ( wire2543 ) | ( _1673 ) | ( _39534 ) ;
 assign _39543 = ( wire2542 ) | ( wire2534 ) | ( wire22262 ) | ( _39540 ) ;
 assign _39546 = ( n_n56  &  wire60 ) | ( wire913  &  n_n56  &  _37743 ) ;
 assign _39552 = ( wire589 ) | ( wire2525 ) | ( _1652 ) | ( _39546 ) ;
 assign _39553 = ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  i_15_ ) ;
 assign _39554 = ( i_14_  &  (~ i_13_)  &  i_12_  &  (~ i_15_) ) ;
 assign _39555 = ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  i_15_ ) ;
 assign _39556 = ( i_14_  &  (~ i_13_)  &  i_12_  &  (~ i_15_) ) ;
 assign _39565 = ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  i_15_ ) ;
 assign _39566 = ( i_14_  &  (~ i_13_)  &  i_12_  &  (~ i_15_) ) ;
 assign _39571 = ( wire22270 ) | ( _39542 ) | ( _39543 ) | ( _39552 ) ;
 assign _39573 = ( i_14_  &  i_13_  &  i_12_ ) ;
 assign _39574 = ( wire898  &  _35695 ) | ( wire904  &  _39573 ) ;
 assign _39576 = ( wire166  &  n_n48 ) | ( wire180  &  n_n48 ) ;
 assign _39578 = ( n_n53  &  wire19385 ) | ( wire900  &  n_n53  &  _35163 ) ;
 assign _39580 = ( n_n4179 ) | ( n_n3843 ) | ( _1626 ) | ( _39576 ) ;
 assign _39582 = ( n_n1137 ) | ( wire2503 ) | ( wire22302 ) | ( _39528 ) ;
 assign _39584 = ( n_n6  &  wire140 ) | ( n_n6  &  wire165 ) ;
 assign _39590 = ( i_14_  &  i_13_  &  i_12_ ) ;
 assign _39594 = ( n_n4858 ) | ( n_n4864 ) | ( _1614 ) | ( _39584 ) ;
 assign _39596 = ( n_n6  &  wire102 ) | ( wire914  &  n_n6  &  _36382 ) ;
 assign _39600 = ( _1591 ) | ( _1592 ) | ( _1599 ) | ( _39596 ) ;
 assign _39601 = ( i_14_  &  i_13_  &  i_12_  &  wire903 ) | ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire903 ) ;
 assign _39632 = ( n_n264  &  n_n285  &  n_n283 ) ;
 assign _39633 = ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  wire902 ) ;
 assign _39645 = ( n_n1240 ) | ( wire22129 ) | ( wire22130 ) | ( wire22148 ) ;
 assign _39646 = ( n_n1242 ) | ( n_n1243 ) | ( wire22142 ) | ( wire22149 ) ;
 assign _39651 = ( n_n1584 ) | ( wire706 ) | ( wire2478 ) | ( wire22317 ) ;
 assign _39653 = ( wire897  &  _35124 ) | ( wire914  &  _39590 ) ;
 assign _39657 = ( wire907  &  _36115 ) | ( wire914  &  _36382 ) ;
 assign _39664 = ( wire22322 ) | ( _1526 ) | ( _1527 ) | ( _39651 ) ;
 assign _39670 = ( wire913  &  _35938 ) | ( wire902  &  _39044 ) ;
 assign _39673 = ( i_14_  &  i_13_  &  i_12_ ) ;
 assign _39674 = ( i_14_  &  i_13_  &  i_12_  &  wire905 ) | ( i_14_  &  i_13_  &  (~ i_12_)  &  wire905 ) ;
 assign _39676 = ( n_n1536 ) | ( n_n4165 ) ;
 assign _39683 = ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  i_15_ ) ;
 assign _39684 = ( i_14_  &  (~ i_13_)  &  i_12_  &  (~ i_15_) ) ;
 assign _39690 = ( i_14_  &  i_13_  &  i_12_  &  wire903 ) | ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire903 ) ;
 assign _39702 = ( (~ i_14_)  &  i_13_  &  i_12_  &  wire897 ) ;
 assign _39703 = ( i_14_  &  i_13_  &  i_12_  &  (~ i_15_) ) ;
 assign _39704 = ( i_14_  &  i_13_  &  (~ i_12_)  &  i_15_ ) ;
 assign _39707 = ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  (~ i_15_) ) ;
 assign _39708 = ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  i_15_ ) ;
 assign _39722 = ( n_n260  &  n_n285  &  n_n263 ) ;
 assign _39740 = ( wire899  &  n_n256 ) | ( wire903  &  _35101 ) ;
 assign _39743 = ( n_n1633 ) | ( wire2601 ) | ( wire140  &  _39722 ) ;
 assign _39744 = ( n_n1628 ) | ( n_n2732 ) | ( wire22185 ) | ( wire2623 ) ;
 assign _39746 = ( i_14_  &  (~ i_13_)  &  i_12_  &  wire907 ) ;
 assign _39749 = ( n_n260  &  n_n285  &  n_n263 ) ;
 assign _39750 = ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  wire912 ) ;
 assign _39753 = ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  i_15_ ) ;
 assign _39754 = ( i_14_  &  (~ i_13_)  &  i_12_  &  (~ i_15_) ) ;
 assign _39758 = ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  i_15_ ) ;
 assign _39759 = ( i_14_  &  (~ i_13_)  &  i_12_  &  (~ i_15_) ) ;
 assign _39772 = ( i_14_  &  i_13_  &  i_12_  &  wire906 ) | ( i_14_  &  i_13_  &  (~ i_12_)  &  wire906 ) ;
 assign _39785 = ( n_n1284 ) | ( wire22219 ) | ( wire22220 ) | ( wire22227 ) ;
 assign _39786 = ( n_n1286 ) | ( wire2593 ) | ( wire2594 ) | ( wire22228 ) ;
 assign _39788 = ( n_n260  &  n_n285  &  n_n263 ) ;
 assign _39793 = ( i_14_  &  (~ i_13_)  &  i_12_  &  wire901 ) ;
 assign _39796 = ( wire22236 ) | ( wire112  &  _39788 ) ;
 assign _39801 = ( n_n100  &  wire77 ) | ( wire898  &  n_n100  &  _38971 ) ;
 assign _39803 = ( n_n94  &  wire81 ) | ( wire906  &  n_n94  &  _35716 ) ;
 assign _39805 = ( _1354 ) | ( _1360 ) | ( _39801 ) | ( _39803 ) ;
 assign _39807 = ( n_n100  &  wire102 ) | ( wire914  &  n_n100  &  _36382 ) ;
 assign _39809 = ( n_n220  &  wire906 ) | ( wire904  &  _35139 ) ;
 assign _39811 = ( n_n3881 ) | ( wire784 ) | ( _1346 ) | ( _39807 ) ;
 assign _39816 = ( n_n260  &  n_n273  &  n_n285 ) ;
 assign _39817 = ( n_n2  &  _39078 ) | ( wire68  &  _39816 ) ;
 assign _39839 = ( i_14_  &  (~ i_13_)  &  i_12_  &  wire905 ) ;
 assign _39848 = ( i_14_  &  (~ i_13_)  &  i_12_  &  wire900 ) | ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  wire900 ) ;
 assign _39853 = ( i_14_  &  (~ i_13_)  &  i_12_  &  wire914 ) ;
 assign _39860 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire913 ) ;
 assign _39861 = ( wire913  &  _36339 ) | ( wire905  &  _36909 ) ;
 assign _39878 = ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  wire899 ) ;
 assign _39888 = ( n_n4624 ) | ( wire699 ) | ( _1261 ) | ( _1262 ) ;
 assign _39890 = ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  i_15_ ) ;
 assign _39891 = ( i_14_  &  (~ i_13_)  &  i_12_  &  (~ i_15_) ) ;
 assign _39892 = ( n_n5  &  wire220 ) | ( n_n5  &  wire22024 ) ;
 assign _39893 = ( wire913  &  _35938 ) | ( wire914  &  _37163 ) ;
 assign _39897 = ( n_n4828 ) | ( n_n1476 ) | ( _1251 ) | ( _39892 ) ;
 assign _39902 = ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  i_15_ ) ;
 assign _39903 = ( i_14_  &  (~ i_13_)  &  i_12_  &  (~ i_15_) ) ;
 assign _39906 = ( wire2774 ) | ( n_n6  &  wire223 ) | ( n_n6  &  wire22033 ) ;
 assign _39908 = ( wire22020 ) | ( wire2777 ) | ( _39888 ) | ( _39897 ) ;
 assign _39925 = ( i_14_  &  (~ i_13_)  &  i_12_  &  wire897 ) | ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  wire897 ) ;
 assign _39929 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire904 ) | ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  wire904 ) ;
 assign _39934 = ( i_14_  &  (~ i_13_)  &  i_12_  &  wire912 ) | ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  wire912 ) ;
 assign _39937 = ( i_14_  &  (~ i_13_)  &  i_12_  &  wire912 ) | ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  wire912 ) ;
 assign _39950 = ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  i_15_ ) ;
 assign _39951 = ( i_14_  &  (~ i_13_)  &  i_12_  &  (~ i_15_) ) ;
 assign _39957 = ( wire902  &  _35651 ) | ( wire911  &  _36330 ) ;
 assign _39959 = ( wire913  &  n_n279 ) | ( wire911  &  _36343 ) ;
 assign _39961 = ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  i_15_ ) ;
 assign _39962 = ( i_14_  &  (~ i_13_)  &  i_12_  &  (~ i_15_) ) ;
 assign _40013 = ( n_n1  &  wire41 ) | ( n_n1  &  wire898  &  _35646 ) ;
 assign _40015 = ( i_14_  &  (~ i_13_)  &  i_12_  &  i_15_ ) ;
 assign _40016 = ( i_14_  &  i_13_  &  i_12_  &  (~ i_15_) ) ;
 assign _40037 = ( wire914  &  _36382 ) | ( wire912  &  _37022 ) ;
 assign _40041 = ( n_n1  &  wire166 ) | ( n_n1  &  wire358 ) ;
 assign _40056 = ( wire2260 ) | ( _1102 ) | ( _40041 ) ;
 assign _40059 = ( wire2258 ) | ( n_n408 ) | ( wire22524 ) | ( _40013 ) ;
 assign _40065 = ( n_n268  &  wire403 ) | ( n_n268  &  wire292 ) ;
 assign _40066 = ( i_14_  &  (~ i_13_)  &  i_12_  &  i_15_ ) ;
 assign _40067 = ( i_14_  &  i_13_  &  i_12_  &  (~ i_15_) ) ;
 assign _40068 = ( i_14_  &  (~ i_13_)  &  i_12_  &  i_15_ ) ;
 assign _40069 = ( i_14_  &  i_13_  &  i_12_  &  (~ i_15_) ) ;
 assign _40070 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  i_15_ ) ;
 assign _40071 = ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  (~ i_15_) ) ;
 assign _40072 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire904 ) | ( i_14_  &  i_13_  &  (~ i_12_)  &  wire904 ) ;
 assign _40078 = ( i_14_  &  (~ i_13_)  &  i_12_  &  wire907 ) | ( i_14_  &  i_13_  &  (~ i_12_)  &  wire907 ) ;
 assign _40080 = ( _1051 ) | ( _1064 ) | ( _40065 ) ;
 assign _40086 = ( n_n2  &  wire140 ) | ( n_n2  &  wire182 ) ;
 assign _40103 = ( wire897  &  _35544 ) | ( wire911  &  _36343 ) ;
 assign _40109 = ( _1010 ) | ( n_n268  &  wire405 ) ;
 assign _40110 = ( wire22537 ) | ( wire2235 ) | ( _40086 ) ;
 assign _40111 = ( wire22533 ) | ( wire22543 ) | ( _40080 ) | ( _40109 ) ;
 assign _40115 = ( n_n94  &  wire403 ) | ( n_n94  &  wire110 ) ;
 assign _40124 = ( i_14_  &  (~ i_13_)  &  i_12_  &  i_15_ ) ;
 assign _40125 = ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  (~ i_15_) ) ;
 assign _40133 = ( i_14_  &  (~ i_13_)  &  i_12_  &  i_15_ ) ;
 assign _40134 = ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  (~ i_15_) ) ;
 assign _40140 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  (~ i_15_) ) ;
 assign _40142 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  i_15_ ) ;
 assign _40160 = ( wire2403 ) | ( wire22389 ) | ( _945 ) | ( _946 ) ;
 assign _40161 = ( wire22383 ) | ( wire22378 ) | ( wire22379 ) | ( wire22380 ) ;
 assign _40165 = ( n_n264  &  n_n285  &  n_n283 ) ;
 assign _40166 = ( i_14_  &  (~ i_13_)  &  i_12_  &  wire913 ) ;
 assign _40169 = ( wire1737  &  _40165 ) | ( wire185  &  _40166 ) ;
 assign _40173 = ( wire22409 ) | ( n_n48  &  wire187 ) | ( n_n48  &  wire22407 ) ;
 assign _40183 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire904 ) ;
 assign _40190 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_ ) ;
 assign _40195 = ( wire900  &  _35163 ) | ( wire906  &  _40190 ) ;
 assign _40198 = ( _899 ) | ( _900 ) | ( n_n6  &  _40183 ) ;
 assign _40200 = ( n_n431 ) | ( wire22412 ) | ( wire22400 ) | ( _40173 ) ;
 assign _40201 = ( n_n429 ) | ( wire22401 ) | ( wire2364 ) | ( _40198 ) ;
 assign _40205 = ( i_14_  &  (~ i_13_)  &  i_12_  &  wire899 ) ;
 assign _40208 = ( i_14_  &  (~ i_13_)  &  i_12_  &  wire902 ) ;
 assign _40217 = ( i_14_  &  (~ i_13_)  &  i_12_  &  i_15_ ) ;
 assign _40218 = ( i_14_  &  i_13_  &  i_12_  &  (~ i_15_) ) ;
 assign _40226 = ( wire900  &  _35163 ) | ( wire905  &  _36909 ) ;
 assign _40229 = ( n_n208  &  n_n284  &  n_n285 ) ;
 assign _40232 = ( i_14_  &  i_13_  &  i_12_  &  wire906 ) ;
 assign _40234 = ( wire22561 ) | ( wire22562 ) | ( wire22565 ) | ( wire2183 ) ;
 assign _40239 = ( wire913  &  _36156 ) | ( wire911  &  _36844 ) ;
 assign _40242 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire905 ) ;
 assign _40245 = ( n_n285  &  n_n230  &  n_n261 ) ;
 assign _40246 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire905 ) | ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire905 ) ;
 assign _40248 = ( n_n6  &  _40242 ) | ( wire1647  &  _40245 ) ;
 assign _40249 = ( _822 ) | ( _833 ) | ( _834 ) | ( _40248 ) ;
 assign _40250 = ( wire904  &  _35141 ) | ( wire901  &  _36986 ) ;
 assign _40252 = ( n_n5  &  wire233 ) | ( n_n5  &  wire22429 ) ;
 assign _40253 = ( i_14_  &  (~ i_13_)  &  i_12_  &  i_15_ ) ;
 assign _40254 = ( i_14_  &  i_13_  &  i_12_  &  (~ i_15_) ) ;
 assign _40255 = ( i_14_  &  i_13_  &  (~ i_12_)  &  (~ i_15_) ) ;
 assign _40258 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire914 ) ;
 assign _40259 = ( n_n247  &  _36092 ) | ( n_n247  &  _36093 ) | ( n_n247  &  _40255 ) ;
 assign _40262 = ( wire2353 ) | ( _808 ) | ( n_n6  &  _40258 ) ;
 assign _40264 = ( i_14_  &  (~ i_13_)  &  i_12_  &  i_15_ ) ;
 assign _40265 = ( i_14_  &  i_13_  &  i_12_  &  (~ i_15_) ) ;
 assign _40266 = ( wire908  &  _35079 ) | ( wire902  &  _35622 ) ;
 assign _40268 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  i_15_ ) ;
 assign _40269 = ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  (~ i_15_) ) ;
 assign _40272 = ( wire902  &  _35622 ) | ( wire903  &  _36705 ) ;
 assign _40274 = ( n_n5  &  wire276 ) | ( n_n5  &  wire22436 ) ;
 assign _40275 = ( wire2361 ) | ( _788 ) | ( _801 ) | ( _40274 ) ;
 assign _40276 = ( wire2356 ) | ( wire2344 ) | ( _40249 ) | ( _40275 ) ;
 assign _40288 = ( wire22446 ) | ( wire2336 ) | ( wire22443 ) | ( _774 ) ;
 assign _40294 = ( wire22454 ) | ( wire166  &  n_n48 ) | ( n_n48  &  wire229 ) ;
 assign _40307 = ( n_n438 ) | ( wire22463 ) | ( _40288 ) ;
 assign _40308 = ( n_n443 ) | ( wire22457 ) | ( wire22464 ) | ( _40294 ) ;
 assign _40311 = ( wire907  &  n_n258 ) | ( n_n258  &  wire899 ) ;
 assign _40313 = ( _716 ) | ( _725 ) | ( _726 ) | ( _727 ) ;
 assign _40322 = ( n_n57  &  wire42 ) | ( n_n57  &  wire899  &  _36360 ) ;
 assign _40330 = ( n_n285  &  n_n271  &  n_n230 ) ;
 assign _40336 = ( i_14_  &  (~ i_13_)  &  i_12_  &  wire897 ) ;
 assign _40337 = ( wire2306 ) | ( n_n56  &  wire53 ) | ( n_n56  &  _40336 ) ;
 assign _40338 = ( _696 ) | ( _40322 ) | ( wire1259  &  _40330 ) ;
 assign _40340 = ( wire2304 ) | ( wire2305 ) | ( _40337 ) | ( _40338 ) ;
 assign _40342 = ( wire898  &  n_n100  &  _35646 ) | ( wire898  &  n_n94  &  _35646 ) ;
 assign _40345 = ( i_15_  &  n_n256  &  n_n253 ) | ( (~ i_15_)  &  n_n256  &  n_n253 ) | ( i_15_  &  n_n256  &  n_n267 ) | ( (~ i_15_)  &  n_n256  &  n_n267 ) ;
 assign _40347 = ( wire2296 ) | ( wire22483 ) | ( wire20755 ) | ( _40342 ) ;
 assign _40371 = ( _6592 ) | ( wire913  &  n_n220 ) | ( n_n220  &  wire905 ) ;
 assign _40373 = ( (~ i_9_)  &  (~ i_10_)  &  (~ i_11_)  &  (~ i_15_) ) ;
 assign _40375 = ( (~ i_9_)  &  (~ i_10_)  &  (~ i_11_)  &  i_15_ ) ;
 assign _40381 = ( i_14_  &  (~ i_13_)  &  i_12_  &  wire902 ) ;
 assign _40385 = ( wire112  &  _39788 ) | ( n_n100  &  _40381 ) ;
 assign _40391 = ( wire22487 ) | ( wire22493 ) | ( wire22494 ) | ( _40347 ) ;
 assign _40392 = ( wire22504 ) | ( _40307 ) | ( _40308 ) | ( _40391 ) ;
 assign _40393 = ( n_n363 ) | ( n_n370 ) | ( _40276 ) | ( _40340 ) ;
 assign _40394 = ( wire22527 ) | ( _40059 ) | ( _40110 ) | ( _40111 ) ;
 assign _40395 = ( n_n346 ) | ( n_n343 ) | ( n_n341 ) | ( _40394 ) ;
 assign _40397 = ( n_n4  &  wire143 ) | ( wire905  &  n_n4  &  _36909 ) ;
 assign _40404 = ( _632 ) | ( _40397 ) | ( n_n3  &  wire1213 ) ;
 assign _40405 = ( wire900  &  _35163 ) | ( wire901  &  _36986 ) ;
 assign _40407 = ( n_n3  &  wire233 ) | ( n_n3  &  wire906  &  _40190 ) ;
 assign _40408 = ( wire900  &  _35163 ) | ( n_n247  &  _40255 ) ;
 assign _40410 = ( n_n4  &  wire351 ) | ( wire914  &  n_n4  &  _36202 ) ;
 assign _40411 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire904 ) ;
 assign _40412 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire906 ) ;
 assign _40413 = ( i_14_  &  (~ i_13_)  &  i_12_  &  wire900 ) ;
 assign _40414 = ( n_n3  &  _40411 ) | ( n_n4  &  _40412 ) ;
 assign _40416 = ( _614 ) | ( _617 ) | ( _40407 ) | ( _40410 ) ;
 assign _40418 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire903 ) | ( i_14_  &  i_13_  &  (~ i_12_)  &  wire903 ) ;
 assign _40420 = ( wire902  &  _35622 ) | ( wire901  &  _36986 ) ;
 assign _40422 = ( n_n4  &  wire233 ) | ( wire907  &  n_n4  &  _36210 ) ;
 assign _40425 = ( wire22351 ) | ( _605 ) | ( _608 ) | ( _40422 ) ;
 assign _40441 = ( wire22348 ) | ( wire22356 ) | ( _40416 ) | ( _40425 ) ;
 assign _40442 = ( wire22594 ) | ( wire590 ) | ( wire19306 ) | ( _34942 ) ;
 assign _40472 = ( (~ i_9_)  &  (~ i_10_)  &  (~ i_11_)  &  (~ i_15_) ) ;
 assign _40474 = ( (~ i_9_)  &  (~ i_10_)  &  (~ i_11_)  &  i_15_ ) ;
 assign _40517 = ( wire461 ) | ( wire2008 ) | ( wire2001 ) | ( _506 ) ;
 assign _40518 = ( wire670 ) | ( wire2002 ) | ( wire22720 ) | ( _492 ) ;
 assign _40536 = ( wire898  &  _35693 ) | ( wire901  &  _36790 ) ;
 assign _40538 = ( n_n5  &  wire134 ) | ( n_n5  &  wire901  &  _36786 ) ;
 assign _40544 = ( (~ i_14_)  &  i_13_  &  i_12_  &  (~ i_15_) ) ;
 assign _40546 = ( (~ i_14_)  &  i_13_  &  i_12_  &  i_15_ ) ;
 assign _40548 = ( i_14_  &  (~ i_13_)  &  i_12_  &  wire900 ) ;
 assign _40564 = ( i_14_  &  (~ i_13_)  &  i_12_  &  i_15_ ) ;
 assign _40565 = ( i_14_  &  i_13_  &  i_12_  &  (~ i_15_) ) ;
 assign _40568 = ( n_n100  &  n_n36 ) | ( wire901  &  n_n100  &  _36786 ) ;
 assign _40573 = ( n_n260  &  n_n285  &  n_n263 ) ;
 assign _40584 = ( i_14_  &  i_13_  &  i_12_  &  wire901 ) | ( i_14_  &  (~ i_13_)  &  i_12_  &  wire901 ) | ( i_14_  &  i_13_  &  (~ i_12_)  &  wire901 ) ;
 assign _40602 = ( n_n53  &  wire275 ) | ( n_n53  &  wire305 ) ;
 assign _40604 = ( n_n952 ) | ( wire543 ) | ( wire550 ) | ( _40602 ) ;
 assign _40607 = ( n_n2  &  wire262 ) | ( n_n2  &  wire304 ) ;
 assign _40618 = ( n_n1  &  wire224 ) | ( n_n1  &  wire335 ) ;
 assign _40620 = ( n_n2  &  wire277 ) | ( n_n2  &  wire356 ) ;
 assign _40633 = ( _367 ) | ( _370 ) | ( _40618 ) | ( _40620 ) ;
 assign _40648 = ( wire862 ) | ( wire895 ) | ( wire856 ) | ( _339 ) ;
 assign _40649 = ( wire855 ) | ( _350 ) | ( n_n268  &  wire1254 ) ;
 assign _40657 = ( n_n2  &  wire1606 ) | ( n_n2  &  wire898  &  _35396 ) ;
 assign _40658 = ( wire22778 ) | ( n_n2  &  wire227 ) | ( n_n2  &  wire305 ) ;
 assign _40660 = ( i_14_  &  (~ i_13_)  &  i_12_  &  wire901 ) ;
 assign _40671 = ( n_n4  &  wire134 ) | ( n_n4  &  wire900  &  _35644 ) ;
 assign _40672 = ( wire1976 ) | ( n_n3  &  wire134 ) | ( n_n3  &  _40660 ) ;
 assign _40675 = ( wire22763 ) | ( wire1970 ) | ( wire1971 ) | ( _40633 ) ;
 assign _40676 = ( n_n755 ) | ( n_n756 ) | ( wire22814 ) | ( _40675 ) ;
 assign _40678 = ( wire898  &  _35396 ) | ( wire899  &  _37042 ) ;
 assign _40699 = ( n_n57  &  wire224 ) | ( n_n56  &  wire224 ) ;
 assign _40701 = ( wire2138 ) | ( wire22616 ) | ( wire22618 ) | ( _40699 ) ;
 assign _40706 = ( n_n850 ) | ( wire22625 ) | ( wire22626 ) | ( _40701 ) ;
 assign _40712 = ( n_n56  &  wire275 ) | ( n_n56  &  wire305 ) | ( n_n56  &  wire348 ) ;
 assign _40713 = ( n_n57  &  wire305 ) | ( n_n57  &  wire348 ) ;
 assign _40728 = ( _231 ) | ( _235 ) | ( _40712 ) | ( _40713 ) ;
 assign _40773 = ( n_n5  &  wire114 ) | ( wire911  &  n_n5  &  _36343 ) ;
 assign _40784 = ( _140 ) | ( _40773 ) | ( n_n6  &  wire1637 ) ;
 assign _40796 = ( i_14_  &  (~ i_13_)  &  i_12_  &  wire902 ) | ( i_14_  &  i_13_  &  (~ i_12_)  &  wire902 ) ;
 assign _40807 = ( wire22678 ) | ( wire22685 ) | ( wire22686 ) | ( _40784 ) ;
 assign _40808 = ( n_n771 ) | ( n_n742 ) | ( _40706 ) ;
 assign _40811 = ( n_n741 ) | ( n_n740 ) | ( wire22822 ) | ( _40676 ) ;
 assign _40812 = ( wire902  &  _35420 ) | ( n_n222  &  _36699 ) ;
 assign _40820 = ( i_14_  &  (~ i_13_)  &  i_12_  &  wire902 ) ;
 assign _40828 = ( wire2169 ) | ( n_n3  &  wire120 ) | ( n_n3  &  _40820 ) ;
 assign _40832 = ( n_n229  &  n_n284  &  n_n285 ) ;
 assign _40833 = ( i_14_  &  i_13_  &  i_12_  &  wire911 ) ;
 assign _40836 = ( wire1777  &  _40832 ) | ( wire169  &  _40833 ) ;
 assign _40857 = ( n_n775 ) | ( wire22839 ) | ( wire22843 ) | ( _61 ) ;
 assign _40858 = ( wire2163 ) | ( wire22602 ) | ( wire22844 ) | ( _40828 ) ;
 assign _40859 = ( wire22847 ) | ( wire590 ) | ( wire19306 ) | ( _34942 ) ;


endmodule

