module seq_mapped (
	i_40_, i_30_, i_20_, i_9_, i_10_, i_7_, i_8_, i_5_, 
	i_6_, i_27_, i_14_, i_3_, i_39_, i_28_, i_13_, i_4_, i_25_, i_12_, 
	i_1_, i_26_, i_11_, i_2_, i_23_, i_18_, i_24_, i_17_, i_0_, i_21_, 
	i_16_, i_22_, i_15_, i_32_, i_31_, i_34_, i_33_, i_19_, i_36_, i_35_, 
	i_38_, i_29_, i_37_, o_1_, o_19_, o_2_, o_0_, o_29_, o_25_, o_12_, 
	o_26_, o_11_, o_27_, o_14_, o_28_, o_13_, o_34_, o_21_, o_16_, o_33_, 
	o_22_, o_15_, o_32_, o_23_, o_18_, o_31_, o_24_, o_17_, o_30_, o_20_, 
	o_10_, o_9_, o_7_, o_8_, o_5_, o_6_, o_3_, o_4_);

input i_40_, i_30_, i_20_, i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_27_, i_14_, i_3_, i_39_, i_28_, i_13_, i_4_, i_25_, i_12_, i_1_, i_26_, i_11_, i_2_, i_23_, i_18_, i_24_, i_17_, i_0_, i_21_, i_16_, i_22_, i_15_, i_32_, i_31_, i_34_, i_33_, i_19_, i_36_, i_35_, i_38_, i_29_, i_37_;

output o_1_, o_19_, o_2_, o_0_, o_29_, o_25_, o_12_, o_26_, o_11_, o_27_, o_14_, o_28_, o_13_, o_34_, o_21_, o_16_, o_33_, o_22_, o_15_, o_32_, o_23_, o_18_, o_31_, o_24_, o_17_, o_30_, o_20_, o_10_, o_9_, o_7_, o_8_, o_5_, o_6_, o_3_, o_4_;

wire wire6758, wire6759, wire1867, wire1870, wire6767, wire6770, n_n1165, wire6806, wire6807, wire6808, n_n1081, wire6914, wire6915, wire6929, wire1693, wire6933, wire6934, wire6935, n_n1581, wire6987, n_n685, wire6991, wire6994, wire6998, n_n1628, n_n1630, n_n1631, wire225, n_n1971, wire7043, n_n1011, n_n1074, n_n864, n_n1711, wire7094, wire7095, wire1505, wire7110, n_n1005, wire566, wire7118, wire7119, n_n1670, wire7190, wire7211, wire7223, n_n979, wire88, n_n1549, n_n1552, wire7270, wire7271, n_n1445, wire7301, wire570, wire7359, n_n2581, n_n1651, wire571, wire7463, wire7478, wire7508, wire1031, wire1044, wire7529, wire7530, wire7540, wire7541, wire7547, wire7548, n_n883, n_n966, n_n1012, wire7550, n_n1272, wire7615, wire7616, wire7639, n_n1330, n_n1332, n_n1187, n_n1184, wire7763, wire7764, n_n1233, wire56, wire7821, wire7822, n_n955, n_n709, wire66, wire334, wire145, wire363, n_n1014, wire45, n_n1009, wire37, wire543, n_n1055, n_n985, wire471, wire80, n_n515, n_n1008, n_n842, n_n1067, n_n982, n_n990, wire330, wire1890, wire1891, wire6772, n_n1373, wire1852, wire1853, wire1854, wire1855, n_n1164, wire1846, wire6793, wire48, n_n1061, wire241, wire6731, wire432, wire491, wire549, n_n2836, wire6818, n_n978, n_n998, n_n1021, n_n330, n_n969, n_n997, n_n793, n_n1048, n_n1047, n_n2487, n_n973, n_n158, n_n977, n_n2488, wire6831, wire6832, n_n1084, wire50, wire6920, n_n1777, wire35, n_n469, n_n1002, n_n795, n_n1993, n_n853, n_n850, wire553, n_n975, wire6938, n_n971, n_n967, wire79, wire115, wire127, wire6940, wire6941, wire6942, wire185, wire6964, wire6965, n_n1986, wire1666, wire173, n_n1607, wire1653, wire6981, n_n926, n_n970, wire318, n_n1990, n_n1072, n_n1951, wire6828, wire6897, wire555, n_n861, wire325, n_n2213, wire92, wire1626, n_n933, n_n1066, wire319, wire422, wire82, wire556, n_n761, wire87, n_n760, n_n1611, wire174, wire1610, wire7025, wire7026, wire300, wire7029, wire7030, n_n833, wire175, wire54, wire240, wire323, n_n1052, wire559, n_n968, wire59, n_n980, n_n1006, n_n989, n_n983, wire1583, wire1584, wire7048, n_n1709, n_n1716, wire1575, wire7053, wire7071, wire445, wire560, n_n865, wire1518, wire47, n_n880, n_n629, wire390, wire7115, wire411, wire436, wire526, n_n991, wire346, wire326, wire565, wire1402, wire7193, wire7194, n_n1528, wire7204, n_n976, n_n668, wire183, wire251, wire354, n_n874, n_n862, wire7237, wire46, wire810, wire7260, wire7261, wire490, n_n1453, n_n1452, wire7329, wire371, n_n837, wire245, wire364, wire348, wire44, wire492, wire7350, n_n1572, wire7384, n_n1414, n_n1412, wire7412, n_n1416, n_n1417, wire7432, wire7444, wire7445, n_n819, wire1132, wire7453, wire7454, wire99, wire365, wire572, wire1062, wire7498, n_n1489, n_n693, wire6821, wire182, n_n1023, wire301, wire574, wire474, wire7512, wire7517, wire575, n_n411, wire407, wire39, wire478, wire6798, n_n1372, wire42, wire1834, wire57, wire84, wire416, wire512, wire317, wire579, n_n949, wire7128, n_n937, wire473, wire739, n_n1374, wire120, n_n1001, n_n945, wire6789, wire7133, wire333, wire6907, wire386, n_n947, wire583, wire581, wire7531, wire146, n_n698, n_n1056, wire7626, wire131, wire402, wire495, n_n334, wire619, wire882, wire7643, wire7649, wire7650, n_n866, wire849, wire7669, wire7674, wire316, n_n848, wire587, wire94, wire106, wire7679, wire586, n_n1197, n_n1203, n_n1202, wire7737, wire7738, wire202, n_n462, wire406, n_n1237, n_n1239, n_n775, wire400, n_n785, wire129, wire7816, n_n1242, wire469, n_n528, n_n888, wire315, n_n313, wire6887, wire227, wire594, wire869, wire7654, wire68, wire504, n_n960, wire367, wire479, wire430, wire78, wire6858, wire957, wire7577, wire7578, n_n1283, wire176, wire7145, wire395, wire598, wire596, wire983, wire595, wire7559, wire7560, n_n1280, n_n1064, n_n525, wire464, wire148, wire329, wire357, wire408, wire441, n_n1073, n_n843, wire542, n_n764, wire600, wire7570, wire7571, wire7574, n_n799, wire366, wire662, wire7774, wire203, wire7784, wire7785, wire7786, n_n710, n_n715, wire602, wire7799, wire7800, n_n1235, wire420, wire160, wire7809, wire607, n_n1094, n_n2837, n_n1958, n_n1956, n_n1957, n_n964, n_n993, wire81, wire382, wire86, n_n642, n_n1015, n_n559, wire320, n_n535, wire7405, wire359, n_n952, n_n935, n_n329, n_n527, n_n688, n_n700, n_n492, wire100, n_n1065, n_n488, n_n453, wire77, wire378, n_n884, n_n928, n_n951, n_n860, n_n560, wire76, n_n484, wire60, wire401, wire465, wire103, n_n791, wire531, wire352, wire7414, wire611, wire1179, wire1181, wire1183, wire7417, wire6850, wire613, wire271, n_n777, n_n781, wire6851, wire64, wire321, wire1786, wire614, n_n1057, wire61, wire7390, n_n162, n_n801, n_n428, n_n427, wire7399, n_n907, wire6716, n_n905, wire1204, wire1205, wire1206, wire7392, wire1196, wire1197, wire1198, wire7403, wire7122, wire467, n_n164, wire1192, wire616, wire615, n_n475, wire7406, wire696, wire7427, wire113, wire617, wire506, wire433, wire7648, wire7330, n_n2439, wire624, wire421, n_n1053, wire627, wire294, wire295, wire297, wire7715, wire36, wire451, wire454, wire7692, wire633, wire446, wire7394, wire154, wire635, wire65, wire638, wire637, wire1913, wire6734, n_n1135, n_n582, n_n771, wire368, wire6859, wire369, wire7389, wire468, wire6976, wire83, wire356, wire643, wire950, wire952, wire7582, wire7583, n_n1285, wire486, wire648, wire646, n_n923, wire286, wire287, wire288, wire289, n_n1068, wire303, wire73, wire520, wire655, wire835, wire336, n_n458, n_n643, wire1681, wire1682, n_n836, wire660, wire43, wire53, wire7772, wire351, wire463, wire666, wire665, wire664, wire153, wire6773, wire184, wire6774, wire187, wire458, wire669, wire668, wire327, wire670, wire671, wire672, wire529, wire370, n_n918, n_n556, n_n798, n_n859, wire674, wire403, wire677, wire1160, wire676, wire7397, wire69, wire332, wire681, wire679, wire678, wire7227, wire7750, wire684, wire484, wire1766, wire6868, wire6869, wire6870, n_n1091, n_n1113, wire244, wire688, wire6878, wire6879, wire1751, wire6886, wire6894, wire711, n_n1108, wire689, wire6908, wire132, wire690, n_n927, n_n773, wire337, wire344, wire693, wire692, wire1173, wire1174, wire695, wire1291, wire102, wire697, wire509, wire342, wire380, wire702, wire701, wire6884, wire700, wire6968, n_n783, wire7309, n_n550, wire855, wire133, wire706, wire710, wire1749, wire1747, wire383, wire429, n_n1577, wire713, wire1099, wire7473, wire7474, wire718, wire717, wire139, wire1277, wire7311, wire488, wire723, wire7319, wire7320, wire7321, wire1269, wire724, wire727, wire7124, wire925, wire926, wire927, wire361, wire450, wire38, wire738, wire737, wire740, n_n1134, wire1901, wire1902, wire742, wire741, wire7191, wire7201, wire124, wire744, wire535, wire749, wire748, wire6974, n_n790, wire166, wire752, wire7154, wire140, wire7146, wire156, wire494, wire758, n_n765, wire761, wire763, wire762, wire767, wire1661, wire1662, wire6970, wire6971, wire101, wire772, wire373, wire7367, wire7371, n_n1575, wire775, wire7132, wire461, wire1487, wire777, wire1489, wire7129, wire7139, wire7140, wire7375, wire7200, wire779, wire782, wire67, wire7150, wire786, wire787, wire6950, wire6951, wire6952, n_n1580, wire788, wire795, wire794, wire826, wire7062, wire158, wire7176, wire6956, wire6957, wire6958, wire803, wire806, wire805, wire808, wire807, wire7258, wire811, wire7256, wire7257, wire809, wire63, wire814, wire818, wire7074, wire817, wire7452, wire822, wire825, wire1570, wire1571, wire7058, wire55, wire304, wire1795, wire1797, wire1798, wire70, wire7818, wire7819, wire104, wire121, wire830, wire829, wire831, wire837, wire375, wire482, wire7510, wire481, wire841, wire840, wire7817, wire546, wire548, wire558, wire589, wire609, wire636, wire642, wire652, wire650, wire687, wire686, wire716, wire715, wire721, wire7007, wire7008, wire729, wire1048, wire731, wire743, wire845, wire1300, wire765, wire1400, wire785, wire793, wire792, wire1563, wire797, wire801, wire7182, wire813, wire820, wire824, wire7815, wire7803, wire142, wire7805, wire143, wire7806, wire144, wire6728, wire151, wire162, wire163, wire164, wire165, wire7796, wire167, wire169, wire170, wire171, wire188, wire190, wire191, wire192, wire193, wire7777, wire198, wire199, wire7276, wire201, wire206, wire207, wire205, wire7767, wire208, wire209, wire210, wire7771, wire211, wire213, wire217, wire218, wire7760, wire229, wire231, wire232, wire234, wire235, wire7743, wire248, wire7745, wire250, wire252, wire260, wire261, wire6739, wire276, wire279, wire7717, wire7707, wire298, wire299, wire7698, wire309, wire310, wire311, wire7689, wire312, wire7694, wire7686, wire455, wire7670, wire519, wire533, wire843, wire538, wire850, wire859, wire860, wire864, wire865, wire872, wire873, wire888, wire7640, wire7627, wire890, wire7630, wire7631, wire892, wire893, wire894, wire904, wire7620, wire905, wire906, wire911, wire912, wire922, wire7610, wire913, wire930, wire932, wire928, wire929, wire934, wire7601, wire7602, wire7593, wire937, wire939, wire940, wire948, wire7586, wire942, wire967, wire7572, wire962, wire964, wire973, wire985, wire987, wire988, wire7127, wire999, wire1000, wire1008, wire1010, wire7521, wire1019, wire7522, wire1020, wire1021, wire1029, wire1022, wire1038, wire1040, wire7514, wire1046, wire7511, wire7500, wire1049, wire1050, wire1051, wire1060, wire1063, wire1075, wire1084, wire1085, wire1083, wire7479, wire1088, wire7482, wire1089, wire1090, wire1091, wire1092, wire1093, wire1112, wire1114, wire7466, wire7467, wire1113, wire1119, wire1120, wire1122, wire7435, wire1155, wire1156, wire1158, wire7347, wire1164, wire1165, wire7415, wire7121, wire1182, wire1186, wire1189, wire1199, wire1200, wire7388, wire1208, wire1219, wire7372, wire1213, wire7360, wire1222, wire1230, wire1238, wire1246, wire1247, wire1251, wire1252, wire7332, wire1253, wire7334, wire1254, wire1255, wire1256, wire1257, wire1262, wire7323, wire7324, wire1264, wire7325, wire1265, wire7314, wire1271, wire7308, wire1286, wire1294, wire1299, wire7291, wire1295, wire7275, wire1305, wire1306, wire7278, wire1307, wire1309, wire7279, wire7281, wire1316, wire1326, wire1317, wire7253, wire1328, wire1329, wire1330, wire7246, wire1340, wire1341, wire1342, wire1343, wire1344, wire7239, wire1346, wire1347, wire1348, wire7231, wire1353, wire1354, wire1362, wire7234, wire1366, wire7214, wire1381, wire1372, wire1374, wire1375, wire7205, wire1383, wire1386, wire1388, wire1389, wire1390, wire7197, wire1412, wire7181, wire1415, wire1416, wire1417, wire1428, wire1429, wire1430, wire7164, wire1442, wire1444, wire7165, wire7157, wire1452, wire1453, wire1454, wire7063, wire7148, wire1459, wire1466, wire1472, wire7142, wire1467, wire1468, wire1496, wire1499, wire1501, wire7103, wire7104, wire7105, wire7108, wire7097, wire1522, wire7089, wire7090, wire1524, wire1525, wire1539, wire1540, wire1541, wire1546, wire1547, wire1542, wire7073, wire1548, wire1550, wire1551, wire1552, wire7064, wire1555, wire1562, wire7067, wire1557, wire7055, wire1565, wire7057, wire1566, wire1568, wire1577, wire1578, wire7052, wire1592, wire1620, wire7016, wire1624, wire7011, wire1632, wire6999, wire1635, wire1657, wire6978, wire6979, wire6945, wire1700, wire1701, wire6930, wire1704, wire1705, wire1707, wire1708, wire1709, wire1730, wire1731, wire6890, wire1741, wire1742, wire6874, wire1758, wire6842, wire1780, wire6839, wire1793, wire6841, wire6824, wire1803, wire1804, wire1806, wire1807, wire1812, wire6800, wire1821, wire1822, wire1832, wire6801, wire1823, wire1839, wire1835, wire1836, wire6791, wire1845, wire1850, wire1847, wire6780, wire1860, wire1861, wire1862, wire1863, wire1878, wire1871, wire1872, wire6766, wire6749, wire1880, wire6750, wire1881, wire1882, wire1883, wire1884, wire1896, wire6736, wire1905, wire1909, wire6727, wire1910, wire6729, wire1911, wire1914, wire1926, wire1923, wire1933, wire1935, wire1936, wire6719, wire6722, wire6726, wire6746, wire6747, wire6753, wire6754, wire6757, wire6764, wire6778, wire6779, wire6786, wire6788, wire6790, wire6804, wire6844, wire6845, wire6849, wire6853, wire6854, wire6856, wire6857, wire6860, wire6861, wire6863, wire6865, wire6866, wire6873, wire6877, wire6901, wire6902, wire6904, wire6909, wire6910, wire6911, wire6924, wire6925, wire6927, wire6932, wire6948, wire6960, wire6961, wire6969, wire6975, wire6980, wire6985, wire6993, wire7001, wire7002, wire7014, wire7020, wire7033, wire7034, wire7035, wire7038, wire7044, wire7066, wire7069, wire7077, wire7079, wire7086, wire7087, wire7092, wire7100, wire7102, wire7123, wire7125, wire7130, wire7131, wire7135, wire7137, wire7143, wire7151, wire7153, wire7160, wire7161, wire7170, wire7178, wire7180, wire7184, wire7185, wire7189, wire7208, wire7218, wire7219, wire7220, wire7230, wire7233, wire7245, wire7252, wire7263, wire7265, wire7266, wire7269, wire7284, wire7285, wire7286, wire7293, wire7299, wire7304, wire7305, wire7306, wire7317, wire7333, wire7336, wire7337, wire7339, wire7341, wire7343, wire7344, wire7348, wire7349, wire7353, wire7354, wire7355, wire7356, wire7373, wire7377, wire7378, wire7411, wire7416, wire7420, wire7421, wire7423, wire7428, wire7430, wire7440, wire7441, wire7442, wire7446, wire7450, wire7456, wire7458, wire7459, wire7460, wire7476, wire7487, wire7488, wire7493, wire7494, wire7495, wire7504, wire7506, wire7518, wire7523, wire7524, wire7535, wire7538, wire7542, wire7544, wire7545, wire7554, wire7555, wire7558, wire7562, wire7563, wire7564, wire7565, wire7566, wire7568, wire7576, wire7588, wire7590, wire7591, wire7596, wire7597, wire7612, wire7614, wire7625, wire7636, wire7641, wire7645, wire7646, wire7658, wire7659, wire7661, wire7663, wire7664, wire7666, wire7667, wire7673, wire7676, wire7677, wire7680, wire7681, wire7704, wire7722, wire7728, wire7734, wire7747, wire7754, wire7755, wire7757, wire7761, wire7762, wire7791, wire7811, wire7814, _35, _38, _40, _41, _43, _44, _46, _53, _54, _56, _57, _60, _61, _63, _66, _78, _79, _86, _101, _105, _110, _111, _112, _113, _114, _115, _116, _119, _120, _122, _123, _124, _125, _129, _130, _131, _132, _145, _148, _149, _158, _159, _162, _163, _165, _172, _173, _175, _176, _177, _193, _195, _196, _207, _208, _213, _214, _218, _219, _221, _223, _224, _226, _231, _245, _250, _294, _295, _297, _320, _334, _335, _380, _381, _384, _385, _387, _406, _407, _408, _409, _410, _430, _431, _435, _440, _441, _452, _453, _456, _479, _485, _488, _494, _512, _513, _524, _525, _547, _554, _555, _567, _573, _593, _618, _619, _620, _621, _625, _626, _713, _714, _722, _725, _731, _733, _742, _743, _745, _765, _766, _768, _772, _775, _781, _782, _783, _785, _788, _789, _790, _791, _792, _805, _808, _809, _835, _836, _838, _848, _849, _856, _857, _881, _892, _893, _915, _943, _954, _959, _960, _962, _968, _970, _979, _982, _983, _984, _1021, _1045, _1046, _1052, _1053, _1063, _1065, _1075, _1076, _1080, _1081, _1171, _1174, _1178, _1204, _1213, _1215, _1216, _1217, _1218, _1219, _1226, _1227, _9032, _9036, _9039, _9041, _9052, _9057, _9080, _9083, _9086, _9110, _9111, _9118, _9119, _9131, _9170, _9179, _9188, _9216, _9236, _9262, _9283, _9284, _9291, _9302, _9303, _9305, _9306, _9322, _9369, _9411, _9416, _9420, _9425, _9430, _9433, _9445, _9451, _9473, _9479, _9483, _9498, _9527, _9531, _9533, _9535, _9543, _9547, _9549, _9552, _9553, _9554, _9555, _9558, _9580, _9598, _9615, _9621, _9636, _9680, _9690, _9694, _9700, _9705, _9715, _9718, _9721, _9723, _9724, _9728, _9732, _9735, _9737, _9741, _9747, _9752, _9755, _9756, _9762, _9769, _9770, _9774, _9785, _9794, _9797, _9801, _9806, _9811, _9823, _9825, _9831, _9879, _9883, _9886, _9905, _9907, _9914, _9917, _9921, _9935, _9966, _9971, _9977, _9980, _9982, _9983, _9987, _9989, _9990, _9999, _10009, _10010, _10011, _10028, _10068, _10069, _10072, _10073, _10082, _10085, _10089, _10093, _10114, _10120, _10125, _10131, _10136, _10141, _10142, _10143, _10151, _10152, _10173, _10177, _10178, _10179, _10180, _10181, _10182, _10186, _10187, _10194, _10207, _10212, _10213, _10233, _10277, _10285, _10296, _10305, _10311, _10330, _10339, _10358, _10361, _10362, _10388, _10392, _10403, _10409, _10411, _10421, _10434, _10435, _10436, _10437, _10483, _10507, _10519, _10525, _10530, _10535, _10542, _10545, _10546, _10547, _10549, _10552, _10554, _10561, _10584, _10586, _10588, _10607, _10613, _10615, _10617, _10634, _10636, _10643, _10651, _10653, _10657, _10668, _10677, _10678, _10691, _10693, _10696, _10699, _10704, _10705, _10712, _10718, _10723, _10724, _10772, _10803, _10804, _10809, _10810, _10818, _10830, _10837, _10867, _10875, _10886, _10890, _10896, _10897, _10899, _10903, _10904, _10925, _10927, _10931, _10933, _10935, _10941, _10943, _10946, _10973, _10982, _10987, _10989, _10991, _11002, _11007, _11009, _11018, _11020, _11022, _11043, _11046, _11057, _11058, _11060, _11064, _11066, _11073, _11074, _11076, _11079, _11080, _11089, _11092, _11094, _11095, _11099, _11107, _11109, _11112, _11116, _11119, _11124, _11128, _11145, _11153, _11155, _11161, _11170, _11184, _11201, _11220, _11232, _11234, _11241, _11244, _11249, _11256, _11261, _11278;

assign o_1_ = ( wire6758 ) | ( wire6759 ) ;
 assign o_19_ = ( wire1867 ) | ( wire1870 ) | ( wire6767 ) | ( wire6770 ) ;
 assign o_2_ = ( n_n1165 ) | ( wire6806 ) | ( wire6807 ) | ( wire6808 ) ;
 assign o_0_ = ( n_n1081 ) | ( wire6914 ) | ( wire6915 ) | ( wire6929 ) ;
 assign o_29_ = ( wire1693 ) | ( wire6933 ) | ( wire6934 ) | ( wire6935 ) ;
 assign o_25_ = ( wire185 ) | ( wire6964 ) | ( wire6965 ) | ( _9715 ) ;
 assign o_12_ = ( _982 ) | ( _983 ) ;
 assign o_26_ = ( wire1635 ) | ( wire7001 ) | ( _9732 ) | ( _9735 ) ;
 assign o_11_ = ( _954 ) | ( _9770 ) | ( wire319  &  _9756 ) ;
 assign o_27_ = ( n_n1607 ) | ( wire7038 ) | ( _9794 ) | ( _9797 ) ;
 assign o_14_ = ( wire225 ) | ( n_n1002  &  n_n975  &  _9801 ) ;
 assign o_28_ = ( n_n1971 ) | ( wire7043 ) | ( _915 ) ;
 assign o_13_ = ( wire225 ) | ( n_n1011  &  n_n1074  &  n_n864 ) ;
 assign o_34_ = ( n_n1711 ) | ( wire7094 ) | ( wire7095 ) ;
 assign o_21_ = ( wire1505 ) | ( _835 ) | ( _836 ) | ( _9921 ) ;
 assign o_16_ = ( wire7118 ) | ( wire7119 ) | ( n_n1005  &  wire566 ) ;
 assign o_33_ = ( n_n1670 ) | ( wire7185 ) | ( _10068 ) | ( _10073 ) ;
 assign o_22_ = ( wire7223 ) | ( wire7204 ) | ( _731 ) | ( _10136 ) ;
 assign o_15_ = ( i_7_  &  i_33_ ) ;
 assign o_32_ = ( n_n1005  &  n_n979  &  wire88 ) ;
 assign o_23_ = ( n_n1549 ) | ( n_n1552 ) | ( wire7270 ) | ( wire7271 ) ;
 assign o_18_ = ( n_n1445 ) | ( wire7344 ) | ( _10361 ) | ( _10362 ) ;
 assign o_31_ = ( wire7359 ) | ( i_22_  &  wire570 ) ;
 assign o_24_ = ( n_n1572 ) | ( wire7384 ) | ( _10409 ) | ( _10411 ) ;
 assign o_17_ = ( n_n1416 ) | ( n_n1417 ) | ( wire7432 ) | ( _10547 ) ;
 assign o_30_ = ( n_n1651 ) | ( wire7463 ) | ( i_24_  &  wire571 ) ;
 assign o_20_ = ( wire7478 ) | ( wire7508 ) | ( _453 ) | ( _10586 ) ;
 assign o_10_ = ( wire1031 ) | ( _380 ) | ( _381 ) | ( _10705 ) ;
 assign o_9_ = ( wire7529 ) | ( wire7530 ) ;
 assign o_7_ = ( wire7540 ) | ( wire7541 ) | ( wire7547 ) | ( wire7548 ) ;
 assign o_8_ = ( wire7550 ) | ( n_n883  &  n_n966  &  n_n1012 ) ;
 assign o_5_ = ( n_n1272 ) | ( wire7615 ) | ( wire7616 ) | ( wire7639 ) ;
 assign o_6_ = ( wire7669 ) | ( wire7674 ) | ( _10973 ) | ( _11009 ) ;
 assign o_3_ = ( n_n1187 ) | ( n_n1184 ) | ( wire7763 ) | ( wire7764 ) ;
 assign o_4_ = ( n_n1233 ) | ( wire56 ) | ( wire7821 ) | ( wire7822 ) ;
 assign wire6758 = ( wire1883 ) | ( wire1923 ) | ( wire6726 ) | ( wire6754 ) ;
 assign wire6759 = ( n_n1135 ) | ( n_n1134 ) | ( wire6747 ) | ( wire6757 ) ;
 assign wire1867 = ( _1178 ) | ( n_n842  &  n_n1067  &  wire1878 ) ;
 assign wire1870 = ( _1174 ) | ( wire546  &  _9188 ) ;
 assign wire6767 = ( _1171 ) | ( n_n979  &  wire88  &  n_n982 ) ;
 assign wire6770 = ( wire1871 ) | ( wire1872 ) | ( n_n515  &  wire6764 ) ;
 assign n_n1165 = ( wire1846 ) | ( wire6793 ) | ( _9236 ) ;
 assign wire6806 = ( n_n1164 ) | ( wire6778 ) | ( wire6779 ) ;
 assign wire6807 = ( n_n1373 ) | ( wire1821 ) | ( wire6804 ) ;
 assign wire6808 = ( n_n1372 ) | ( wire1823 ) | ( wire1835 ) | ( wire1836 ) ;
 assign n_n1081 = ( n_n1091 ) | ( wire6878 ) | ( wire6879 ) ;
 assign wire6914 = ( wire6909 ) | ( wire6910 ) | ( wire6911 ) | ( _9430 ) ;
 assign wire6915 = ( n_n1094 ) | ( wire6904 ) | ( _9531 ) ;
 assign wire6929 = ( wire6818 ) | ( n_n1084 ) | ( wire6927 ) | ( _9554 ) ;
 assign wire1693 = ( wire48  &  wire35  &  wire1700 ) | ( wire48  &  wire35  &  wire1701 ) ;
 assign wire6933 = ( n_n1993 ) | ( n_n1012  &  n_n799  &  wire529 ) ;
 assign wire6934 = ( wire529  &  wire509 ) | ( wire366  &  wire535 ) ;
 assign wire6935 = ( wire509  &  wire535 ) | ( wire553  &  wire6932 ) ;
 assign n_n1581 = ( wire127 ) | ( wire6940 ) | ( wire6941 ) | ( wire6942 ) ;
 assign wire6987 = ( n_n2581 ) | ( wire173 ) | ( wire6985 ) | ( _984 ) ;
 assign n_n685 = ( (~ i_7_)  &  i_5_  &  (~ i_0_) ) ;
 assign wire6991 = ( (~ i_40_)  &  i_8_ ) ;
 assign wire6994 = ( _979 ) | ( i_0_  &  wire79  &  wire6993 ) ;
 assign wire6998 = ( n_n2837 ) | ( n_n1958 ) | ( _9728 ) ;
 assign n_n1628 = ( n_n2487 ) | ( n_n2488 ) | ( wire173 ) | ( n_n1611 ) ;
 assign n_n1630 = ( wire174 ) | ( wire1610 ) | ( wire7025 ) | ( wire7026 ) ;
 assign n_n1631 = ( wire127 ) | ( wire300 ) | ( wire7029 ) | ( wire7030 ) ;
 assign wire225 = ( o_15_ ) | ( n_n1074  &  n_n968  &  wire59 ) ;
 assign n_n1971 = ( n_n971  &  n_n967  &  wire79  &  (~ wire115) ) ;
 assign wire7043 = ( (~ i_40_)  &  (~ i_38_)  &  wire542 ) | ( (~ i_39_)  &  (~ i_38_)  &  wire542 ) ;
 assign n_n1011 = ( (~ i_39_)  &  (~ i_38_) ) ;
 assign n_n1074 = ( (~ i_32_)  &  (~ i_34_)  &  i_33_ ) ;
 assign n_n864 = ( i_36_  &  i_35_  &  (~ i_37_) ) ;
 assign n_n1711 = ( n_n1716 ) | ( wire1575 ) | ( wire7053 ) | ( wire7071 ) ;
 assign wire7094 = ( wire1524 ) | ( wire7077 ) | ( n_n1074  &  wire817 ) ;
 assign wire7095 = ( n_n1709 ) | ( wire7086 ) | ( wire7087 ) | ( wire7092 ) ;
 assign wire1505 = ( wire7103  &  wire7105 ) | ( wire7104  &  wire7105 ) ;
 assign wire7110 = ( (~ i_33_) ) | ( n_n978  &  n_n865  &  wire7100 ) ;
 assign n_n1005 = ( (~ i_39_)  &  i_38_  &  i_37_ ) ;
 assign wire566 = ( i_40_  &  n_n979  &  n_n861 ) | ( (~ i_40_)  &  n_n861  &  n_n991 ) ;
 assign wire7118 = ( wire1499 ) | ( wire526  &  wire565 ) ;
 assign wire7119 = ( wire1496 ) | ( wire1501 ) | ( wire411  &  wire436 ) ;
 assign n_n1670 = ( wire7176 ) | ( wire1429 ) | ( _10010 ) | ( _10028 ) ;
 assign wire7190 = ( wire7189 ) | ( _10072 ) ;
 assign wire7211 = ( wire1383 ) | ( wire1386 ) | ( _722 ) ;
 assign wire7223 = ( n_n1528 ) | ( wire7218 ) | ( wire7219 ) | ( wire7220 ) ;
 assign n_n979 = ( (~ i_34_)  &  (~ i_36_)  &  i_35_ ) ;
 assign wire88 = ( (~ i_40_)  &  (~ i_7_)  &  (~ i_32_)  &  i_33_ ) ;
 assign n_n1549 = ( wire7237 ) | ( _10152 ) ;
 assign n_n1552 = ( wire7260 ) | ( wire7261 ) | ( wire46  &  wire810 ) ;
 assign wire7270 = ( wire7230 ) | ( wire7245 ) | ( _10194 ) ;
 assign wire7271 = ( wire1343 ) | ( wire1344 ) | ( wire7252 ) | ( wire7269 ) ;
 assign n_n1445 = ( n_n1453 ) | ( n_n1452 ) | ( wire7329 ) ;
 assign wire7301 = ( wire7284 ) | ( wire7285 ) | ( wire7286 ) | ( wire7299 ) ;
 assign wire570 = ( wire348  &  wire7350 ) | ( wire348  &  wire44  &  wire492 ) ;
 assign wire7359 = ( wire7353 ) | ( wire7354 ) | ( wire7355 ) | ( wire7356 ) ;
 assign n_n2581 = ( wire88  &  n_n975  &  wire6938 ) ;
 assign n_n1651 = ( wire1132 ) | ( wire7453 ) | ( wire7454 ) ;
 assign wire571 = ( wire348  &  wire7350 ) | ( wire348  &  wire44  &  wire492 ) ;
 assign wire7463 = ( wire1122 ) | ( wire7458 ) | ( wire7459 ) | ( wire7460 ) ;
 assign wire7478 = ( wire251 ) | ( wire1093 ) | ( wire718  &  wire7476 ) ;
 assign wire7508 = ( n_n1489 ) | ( wire7494 ) | ( wire7495 ) | ( wire7506 ) ;
 assign wire1031 = ( _387 ) | ( i_20_  &  i_21_  &  wire1038 ) ;
 assign wire1044 = ( wire35  &  wire7512  &  _10699 ) ;
 assign wire7529 = ( n_n1373 ) | ( n_n1372 ) | ( wire1021 ) | ( wire1022 ) ;
 assign wire7530 = ( wire1019 ) | ( wire1020 ) | ( wire7523 ) | ( wire7524 ) ;
 assign wire7540 = ( wire140 ) | ( _10724 ) | ( wire7123  &  _10723 ) ;
 assign wire7541 = ( wire1412 ) | ( wire7189 ) | ( wire7535 ) | ( wire7538 ) ;
 assign wire7547 = ( n_n1372 ) | ( wire999 ) | ( wire1835 ) | ( wire1836 ) ;
 assign wire7548 = ( n_n1373 ) | ( wire1000 ) | ( wire7544 ) | ( wire7545 ) ;
 assign n_n883 = ( i_40_  &  (~ i_39_)  &  i_38_ ) ;
 assign n_n966 = ( (~ i_32_)  &  i_34_  &  i_33_ ) ;
 assign n_n1012 = ( (~ i_36_)  &  (~ i_35_)  &  i_37_ ) ;
 assign wire7550 = ( o_15_ ) | ( wire45  &  n_n693  &  wire7531 ) ;
 assign n_n1272 = ( n_n1280 ) | ( wire7570 ) | ( wire7571 ) | ( wire7574 ) ;
 assign wire7615 = ( wire927 ) | ( wire912 ) | ( wire913 ) | ( _10809 ) ;
 assign wire7616 = ( n_n1283 ) | ( n_n1285 ) | ( wire7591 ) | ( wire7614 ) ;
 assign wire7639 = ( wire892 ) | ( wire7636 ) | ( _10903 ) | ( _10904 ) ;
 assign n_n1330 = ( wire882 ) | ( wire7643 ) | ( n_n334  &  wire619 ) ;
 assign n_n1332 = ( wire7650 ) | ( _226 ) ;
 assign n_n1187 = ( n_n1197 ) | ( _158 ) | ( _159 ) | ( _11058 ) ;
 assign n_n1184 = ( n_n1203 ) | ( n_n1202 ) | ( wire7737 ) | ( wire7738 ) ;
 assign wire7763 = ( wire7747 ) | ( wire7761 ) | ( _11099 ) ;
 assign wire7764 = ( wire311 ) | ( wire7704 ) | ( wire7762 ) | ( _11161 ) ;
 assign n_n1233 = ( n_n1237 ) | ( n_n1239 ) | ( wire7791 ) | ( _11220 ) ;
 assign wire56 = ( _63 ) | ( _11232 ) ;
 assign wire7821 = ( _60 ) | ( _61 ) | ( n_n427  &  _11234 ) ;
 assign wire7822 = ( n_n1242 ) | ( n_n1235 ) | ( wire7814 ) ;
 assign n_n955 = ( i_9_  &  (~ i_5_)  &  i_11_ ) ;
 assign n_n709 = ( (~ i_38_)  &  (~ i_37_) ) ;
 assign wire66 = ( i_40_  &  i_39_ ) | ( i_39_  &  (~ i_38_) ) ;
 assign wire334 = ( i_35_  &  (~ i_37_) ) ;
 assign wire145 = ( o_15_ ) | ( n_n1074  &  n_n883  &  wire334 ) ;
 assign wire363 = ( (~ i_39_)  &  (~ i_38_)  &  n_n1074  &  n_n1012 ) ;
 assign n_n1014 = ( i_40_  &  i_39_ ) ;
 assign wire45 = ( (~ i_32_)  &  (~ i_34_)  &  i_33_  &  (~ i_35_) ) ;
 assign n_n1009 = ( (~ i_36_)  &  i_38_  &  (~ i_37_) ) ;
 assign wire37 = ( i_17_ ) | ( i_16_ ) ;
 assign wire543 = ( (~ i_40_)  &  i_39_ ) | ( i_39_  &  (~ i_38_) ) ;
 assign n_n1055 = ( (~ i_39_)  &  (~ i_38_)  &  i_37_ ) ;
 assign n_n985 = ( (~ i_36_)  &  (~ i_38_)  &  i_37_ ) ;
 assign wire471 = ( (~ i_3_)  &  (~ i_4_)  &  (~ i_1_)  &  (~ i_2_) ) ;
 assign wire80 = ( (~ i_32_)  &  i_34_  &  i_33_  &  (~ i_35_) ) ;
 assign n_n515 = ( (~ i_7_)  &  wire471  &  wire80 ) ;
 assign n_n1008 = ( (~ i_40_)  &  (~ i_39_) ) ;
 assign n_n842 = ( (~ i_7_)  &  (~ i_3_)  &  i_4_ ) ;
 assign n_n1067 = ( (~ i_1_)  &  (~ i_2_)  &  i_0_ ) ;
 assign n_n982 = ( (~ i_39_)  &  i_38_  &  (~ i_37_) ) ;
 assign n_n990 = ( i_39_  &  (~ i_38_)  &  (~ i_37_) ) ;
 assign wire330 = ( i_40_  &  i_39_  &  (~ i_38_)  &  i_37_ ) ;
 assign wire1890 = ( i_9_  &  (~ i_5_)  &  (~ i_11_)  &  _9039 ) ;
 assign wire1891 = ( i_9_  &  (~ i_5_)  &  i_11_  &  _9036 ) ;
 assign wire6772 = ( n_n1048  &  n_n1047  &  wire400 ) ;
 assign n_n1373 = ( wire1891  &  wire6772 ) | ( wire6772  &  n_n928  &  _9039 ) ;
 assign wire1852 = ( n_n1012  &  n_n799  &  wire668  &  wire6780 ) ;
 assign wire1853 = ( n_n1048  &  n_n1047  &  wire458  &  wire669 ) ;
 assign wire1854 = ( n_n1074  &  n_n968  &  n_n1064  &  n_n884 ) ;
 assign wire1855 = ( wire471  &  n_n998  &  wire46  &  n_n1001 ) ;
 assign n_n1164 = ( wire1852 ) | ( wire1853 ) | ( wire1854 ) | ( wire1855 ) ;
 assign wire1846 = ( n_n528  &  n_n905 ) | ( n_n528  &  wire1850 ) ;
 assign wire6793 = ( (~ i_12_)  &  i_11_  &  wire407  &  wire84 ) | ( i_12_  &  (~ i_11_)  &  wire407  &  wire84 ) ;
 assign wire48 = ( (~ i_21_)  &  i_15_ ) ;
 assign n_n1061 = ( i_36_  &  i_38_  &  (~ i_37_) ) ;
 assign wire241 = ( i_40_  &  (~ i_39_)  &  n_n1074  &  n_n1061 ) ;
 assign wire6731 = ( (~ i_36_)  &  i_35_  &  i_37_ ) ;
 assign wire432 = ( (~ i_39_)  &  (~ i_38_)  &  n_n1074  &  wire6731 ) ;
 assign wire491 = ( i_23_  &  i_24_  &  i_22_  &  i_19_ ) ;
 assign wire549 = ( i_40_  &  (~ i_38_) ) | ( i_39_  &  (~ i_38_) ) ;
 assign n_n2836 = ( (~ i_7_)  &  i_1_  &  wire80  &  n_n926 ) ;
 assign wire6818 = ( n_n2837 ) | ( n_n1958 ) | ( _9552 ) ;
 assign n_n978 = ( i_40_  &  (~ i_39_)  &  (~ i_38_) ) ;
 assign n_n998 = ( i_34_  &  (~ i_36_)  &  (~ i_35_) ) ;
 assign n_n1021 = ( (~ i_40_)  &  i_39_ ) ;
 assign n_n330 = ( (~ i_7_)  &  (~ i_5_)  &  i_13_ ) ;
 assign n_n969 = ( (~ i_40_)  &  (~ i_39_)  &  (~ i_38_) ) ;
 assign n_n997 = ( i_39_  &  i_38_  &  i_37_ ) ;
 assign n_n793 = ( (~ i_9_)  &  (~ i_7_)  &  (~ i_5_) ) ;
 assign n_n1048 = ( (~ i_32_)  &  (~ i_31_)  &  i_33_ ) ;
 assign n_n1047 = ( (~ i_34_)  &  (~ i_36_)  &  (~ i_35_) ) ;
 assign n_n2487 = ( n_n997  &  n_n793  &  n_n1048  &  n_n1047 ) ;
 assign n_n973 = ( i_40_  &  i_39_  &  (~ i_38_) ) ;
 assign n_n158 = ( i_15_  &  (~ i_32_)  &  i_33_ ) ;
 assign n_n977 = ( (~ i_40_)  &  i_39_  &  i_38_ ) ;
 assign n_n2488 = ( n_n793  &  n_n1048  &  n_n1047  &  n_n977 ) ;
 assign wire6831 = ( wire182 ) | ( wire1803 ) | ( wire1807 ) ;
 assign wire6832 = ( wire1804 ) | ( wire1806 ) | ( i_2_  &  wire835 ) ;
 assign n_n1084 = ( wire6831 ) | ( wire6832 ) | ( _1052 ) | ( _1053 ) ;
 assign wire50 = ( (~ i_32_)  &  (~ i_34_)  &  i_33_  &  i_35_ ) ;
 assign wire6920 = ( i_0_  &  (~ i_36_)  &  i_38_  &  i_37_ ) ;
 assign n_n1777 = ( (~ i_7_)  &  wire50  &  wire6920 ) ;
 assign wire35 = ( (~ i_7_)  &  (~ i_5_)  &  i_12_ ) | ( (~ i_7_)  &  (~ i_5_)  &  i_11_ ) ;
 assign n_n469 = ( (~ i_40_)  &  i_39_  &  i_38_  &  (~ i_37_) ) ;
 assign n_n1002 = ( (~ i_34_)  &  i_36_  &  i_35_ ) ;
 assign n_n795 = ( i_39_  &  (~ i_38_)  &  i_37_ ) ;
 assign n_n1993 = ( wire88  &  n_n1002  &  n_n795 ) ;
 assign n_n853 = ( (~ i_7_)  &  (~ i_5_)  &  i_11_ ) ;
 assign n_n850 = ( (~ i_7_)  &  (~ i_5_)  &  i_12_ ) ;
 assign wire553 = ( (~ i_21_)  &  i_15_  &  n_n853 ) | ( (~ i_21_)  &  i_15_  &  n_n850 ) ;
 assign n_n975 = ( (~ i_39_)  &  (~ i_38_)  &  (~ i_37_) ) ;
 assign wire6938 = ( i_34_  &  i_36_  &  (~ i_35_) ) ;
 assign n_n971 = ( i_36_  &  (~ i_35_)  &  (~ i_37_) ) ;
 assign n_n967 = ( (~ i_40_)  &  (~ i_39_)  &  i_38_ ) ;
 assign wire79 = ( (~ i_7_)  &  (~ i_32_)  &  (~ i_34_)  &  i_33_ ) ;
 assign wire115 = ( (~ i_10_) ) | ( (~ i_27_) ) ;
 assign wire127 = ( wire348  &  wire329 ) | ( n_n775  &  n_n781 ) ;
 assign wire6940 = ( n_n1012  &  n_n799  &  wire529 ) | ( n_n1012  &  n_n799  &  wire535 ) ;
 assign wire6941 = ( wire479  &  wire368 ) | ( n_n765  &  wire101 ) ;
 assign wire6942 = ( wire430  &  wire772 ) | ( i_39_  &  (~ i_37_)  &  wire430 ) ;
 assign wire185 = ( wire6956 ) | ( wire6957 ) | ( wire6958 ) ;
 assign wire6964 = ( wire175 ) | ( wire240 ) | ( wire6960 ) | ( wire6961 ) ;
 assign wire6965 = ( n_n1611 ) | ( wire6950 ) | ( wire6951 ) | ( wire6952 ) ;
 assign n_n1986 = ( (~ i_24_)  &  wire50  &  wire87  &  wire371 ) ;
 assign wire1666 = ( (~ i_24_)  &  wire50  &  wire87  &  n_n833 ) ;
 assign wire173 = ( n_n1993 ) | ( n_n1986 ) | ( wire1666 ) ;
 assign n_n1607 = ( wire1661 ) | ( wire1662 ) | ( wire6970 ) | ( wire6971 ) ;
 assign wire1653 = ( wire1657  &  wire6979 ) | ( wire6978  &  wire6979 ) ;
 assign wire6981 = ( n_n783  &  wire6975 ) | ( n_n790  &  wire6975 ) | ( n_n790  &  wire6980 ) ;
 assign n_n926 = ( (~ i_39_)  &  (~ i_36_)  &  (~ i_38_)  &  i_37_ ) ;
 assign n_n970 = ( i_36_  &  (~ i_35_)  &  i_37_ ) ;
 assign wire318 = ( i_1_  &  i_0_ ) ;
 assign n_n1990 = ( n_n883  &  wire79  &  n_n970  &  wire318 ) ;
 assign n_n1072 = ( i_40_  &  i_39_  &  i_38_ ) ;
 assign n_n1951 = ( n_n971  &  wire79  &  wire318  &  n_n1072 ) ;
 assign wire6828 = ( (~ i_7_)  &  i_3_  &  i_0_ ) ;
 assign wire6897 = ( (~ i_7_)  &  i_2_  &  i_0_ ) ;
 assign wire555 = ( n_n1074  &  wire6828 ) | ( n_n1074  &  wire6897 ) ;
 assign n_n861 = ( (~ i_7_)  &  (~ i_32_)  &  i_33_ ) ;
 assign wire325 = ( i_40_  &  i_39_  &  (~ i_38_)  &  (~ i_37_) ) ;
 assign n_n2213 = ( n_n998  &  n_n861  &  wire325 ) ;
 assign wire92 = ( i_40_  &  i_39_  &  n_n1009 ) ;
 assign wire1626 = ( wire48  &  n_n428  &  n_n427  &  wire727 ) ;
 assign n_n933 = ( i_17_  &  (~ i_32_)  &  (~ i_31_) ) ;
 assign n_n1066 = ( (~ i_34_)  &  i_33_  &  (~ i_35_) ) ;
 assign wire319 = ( (~ i_34_)  &  i_33_  &  (~ i_35_)  &  _9747 ) ;
 assign wire422 = ( (~ i_32_)  &  (~ i_31_)  &  i_33_  &  (~ i_35_) ) ;
 assign wire82 = ( (~ i_7_)  &  (~ i_5_)  &  i_11_  &  i_15_ ) ;
 assign wire556 = ( i_40_  &  (~ i_39_)  &  i_38_ ) | ( (~ i_39_)  &  i_38_  &  (~ i_37_) ) ;
 assign n_n761 = ( (~ i_21_)  &  i_15_  &  wire50  &  n_n850 ) ;
 assign wire87 = ( (~ i_7_)  &  (~ i_5_)  &  i_12_  &  i_15_ ) ;
 assign n_n760 = ( (~ i_22_)  &  wire50  &  wire87 ) ;
 assign n_n1611 = ( wire176 ) | ( wire1681 ) | ( wire1682 ) ;
 assign wire174 = ( wire504  &  n_n960 ) | ( wire367  &  wire479 ) ;
 assign wire1610 = ( wire68  &  wire504 ) ;
 assign wire7025 = ( _943 ) | ( (~ i_22_)  &  wire82  &  wire337 ) ;
 assign wire7026 = ( n_n764  &  wire359 ) | ( n_n761  &  wire101 ) | ( n_n764  &  wire101 ) ;
 assign wire300 = ( i_39_  &  i_38_  &  wire430 ) | ( i_40_  &  (~ i_38_)  &  wire430 ) ;
 assign wire7029 = ( wire479  &  wire368 ) | ( wire365  &  wire337 ) ;
 assign wire7030 = ( n_n765  &  wire825 ) | ( wire430  &  wire6863 ) ;
 assign n_n833 = ( i_39_  &  (~ i_36_)  &  i_38_  &  (~ i_37_) ) ;
 assign wire175 = ( (~ i_22_)  &  wire50  &  wire82  &  n_n833 ) ;
 assign wire54 = ( i_39_  &  (~ i_36_)  &  i_38_  &  (~ i_37_) ) | ( (~ i_39_)  &  (~ i_36_)  &  (~ i_38_)  &  (~ i_37_) ) ;
 assign wire240 = ( (~ i_24_)  &  wire50  &  wire82  &  wire54 ) ;
 assign wire323 = ( (~ i_40_)  &  i_39_  &  n_n1009 ) ;
 assign n_n1052 = ( (~ i_36_)  &  (~ i_38_)  &  (~ i_37_) ) ;
 assign wire559 = ( i_40_  &  (~ i_39_)  &  n_n985 ) | ( (~ i_40_)  &  (~ i_39_)  &  n_n1052 ) ;
 assign n_n968 = ( (~ i_36_)  &  i_35_  &  (~ i_37_) ) ;
 assign wire59 = ( (~ i_40_)  &  (~ i_39_)  &  i_38_ ) | ( i_40_  &  i_39_  &  (~ i_38_) ) ;
 assign n_n980 = ( i_5_  &  (~ i_32_)  &  i_33_ ) ;
 assign n_n1006 = ( i_5_  &  (~ i_0_)  &  (~ i_32_) ) ;
 assign n_n989 = ( (~ i_15_)  &  (~ i_32_)  &  (~ i_31_) ) ;
 assign n_n983 = ( (~ i_34_)  &  i_33_  &  (~ i_36_) ) ;
 assign wire1583 = ( i_5_  &  (~ i_36_)  &  wire45  &  wire795 ) ;
 assign wire1584 = ( n_n1047  &  n_n980  &  wire794 ) ;
 assign wire7048 = ( o_15_ ) | ( n_n980  &  wire65  &  wire7044 ) ;
 assign n_n1709 = ( wire1583 ) | ( wire1584 ) | ( wire7048 ) ;
 assign n_n1716 = ( wire7062 ) | ( wire76  &  wire826 ) ;
 assign wire1575 = ( i_17_  &  wire1577 ) | ( i_16_  &  wire1577 ) | ( i_17_  &  wire1578 ) | ( i_16_  &  wire1578 ) ;
 assign wire7053 = ( wire84  &  _892 ) | ( wire84  &  _893 ) | ( wire84  &  _9831 ) ;
 assign wire7071 = ( wire1557 ) | ( wire7069 ) | ( _881 ) ;
 assign wire445 = ( (~ i_40_)  &  (~ i_39_)  &  i_38_  &  (~ i_37_) ) ;
 assign wire560 = ( n_n979  &  n_n978 ) | ( n_n1012  &  n_n973 ) ;
 assign n_n865 = ( i_36_  &  i_35_  &  i_37_ ) ;
 assign wire1518 = ( n_n864  &  n_n1072  &  wire7097 ) ;
 assign wire47 = ( (~ i_7_)  &  (~ i_5_) ) ;
 assign n_n880 = ( i_40_  &  (~ i_38_) ) ;
 assign n_n629 = ( (~ i_7_)  &  (~ i_12_)  &  (~ i_11_) ) ;
 assign wire390 = ( (~ i_7_)  &  (~ i_12_)  &  (~ i_11_)  &  _10657 ) ;
 assign wire7115 = ( i_1_  &  (~ i_2_)  &  i_0_ ) ;
 assign wire411 = ( n_n1074  &  n_n842  &  wire7115 ) ;
 assign wire436 = ( i_36_  &  i_35_  &  i_37_  &  _9935 ) ;
 assign wire526 = ( (~ i_3_)  &  (~ i_4_)  &  n_n1067  &  wire79 ) ;
 assign n_n991 = ( (~ i_34_)  &  i_36_  &  (~ i_35_) ) ;
 assign wire346 = ( (~ i_39_)  &  i_38_ ) ;
 assign wire326 = ( i_36_  &  (~ i_35_) ) ;
 assign wire565 = ( (~ i_37_)  &  n_n1072  &  wire326 ) | ( i_37_  &  wire346  &  wire326 ) ;
 assign wire1402 = ( n_n1066  &  wire166  &  wire7197 ) ;
 assign wire7193 = ( (~ i_17_)  &  (~ i_16_) ) | ( i_38_  &  i_37_ ) ;
 assign wire7194 = ( (~ i_40_)  &  i_38_ ) | ( (~ i_39_)  &  i_38_ ) | ( i_39_  &  (~ i_38_) ) | ( (~ i_38_)  &  (~ i_37_) ) ;
 assign n_n1528 = ( wire1402 ) | ( _713 ) | ( _714 ) ;
 assign wire7204 = ( wire301 ) | ( wire1390 ) | ( _733 ) ;
 assign n_n976 = ( i_33_  &  (~ i_36_)  &  (~ i_35_) ) ;
 assign n_n668 = ( (~ i_7_)  &  i_5_  &  (~ i_32_) ) ;
 assign wire183 = ( wire330  &  n_n976  &  n_n668 ) ;
 assign wire251 = ( n_n975  &  n_n983  &  n_n668 ) ;
 assign wire354 = ( (~ i_34_)  &  (~ i_36_)  &  (~ i_35_)  &  _10089 ) ;
 assign n_n874 = ( (~ i_32_)  &  i_33_  &  (~ i_35_) ) ;
 assign n_n862 = ( (~ i_36_)  &  (~ i_35_)  &  i_38_ ) ;
 assign wire7237 = ( wire1353 ) | ( wire1354 ) | ( n_n880  &  wire803 ) ;
 assign wire46 = ( (~ i_32_)  &  i_33_ ) ;
 assign wire810 = ( wire464  &  wire7256 ) | ( n_n1047  &  wire7257 ) ;
 assign wire7260 = ( wire1328 ) | ( n_n710  &  wire811 ) ;
 assign wire7261 = ( wire1329 ) | ( wire1330 ) | ( wire77  &  wire809 ) ;
 assign wire490 = ( (~ i_34_)  &  (~ i_35_) ) ;
 assign n_n1453 = ( wire1277 ) | ( wire7311 ) | ( n_n559  &  wire139 ) ;
 assign n_n1452 = ( wire7319 ) | ( wire7320 ) | ( wire7321 ) ;
 assign wire7329 = ( wire1264 ) | ( wire1265 ) | ( wire526  &  wire724 ) ;
 assign wire371 = ( i_40_  &  (~ i_39_)  &  (~ i_36_)  &  (~ i_38_) ) ;
 assign n_n837 = ( (~ i_24_)  &  wire50  &  wire82 ) ;
 assign wire245 = ( (~ i_24_)  &  wire50  &  wire87  &  wire54 ) ;
 assign wire364 = ( i_21_  &  i_22_  &  i_15_  &  wire35 ) ;
 assign wire348 = ( wire6731  &  n_n978  &  _9621 ) ;
 assign wire44 = ( wire469 ) | ( i_18_  &  wire35 ) ;
 assign wire492 = ( (~ i_21_)  &  i_15_  &  i_19_ ) ;
 assign wire7350 = ( n_n859  &  wire7349 ) | ( wire1797  &  wire7349 ) | ( wire1798  &  wire7349 ) ;
 assign n_n1572 = ( n_n1577 ) | ( n_n1575 ) | ( wire7375 ) ;
 assign wire7384 = ( n_n1581 ) | ( n_n1113 ) | ( n_n1580 ) | ( wire7377 ) ;
 assign n_n1414 = ( wire1204 ) | ( wire1205 ) | ( wire1206 ) | ( wire7392 ) ;
 assign n_n1412 = ( wire1196 ) | ( wire1197 ) | ( wire1198 ) | ( wire7403 ) ;
 assign wire7412 = ( wire7411 ) | ( n_n1001  &  wire616 ) ;
 assign n_n1416 = ( wire1179 ) | ( wire1181 ) | ( wire1183 ) | ( wire7417 ) ;
 assign n_n1417 = ( wire7427 ) | ( n_n1011  &  n_n1012  &  wire696 ) ;
 assign wire7432 = ( wire7430 ) | ( _10519 ) ;
 assign wire7444 = ( wire332  &  wire678 ) | ( wire679  &  wire7441 ) ;
 assign wire7445 = ( _494 ) | ( n_n1065  &  wire69  &  _10530 ) ;
 assign n_n819 = ( i_24_  &  (~ i_22_)  &  n_n1074  &  wire82 ) ;
 assign wire1132 = ( _485 ) | ( wire824  &  _10549 ) ;
 assign wire7453 = ( n_n819  &  wire386 ) | ( wire99  &  wire7450 ) ;
 assign wire7454 = ( _479 ) | ( n_n968  &  wire132  &  _10561 ) ;
 assign wire99 = ( (~ i_36_)  &  i_35_  &  (~ i_37_)  &  _10554 ) ;
 assign wire365 = ( (~ i_21_)  &  i_15_  &  n_n853 ) ;
 assign wire572 = ( (~ i_40_)  &  i_39_  &  i_38_ ) | ( (~ i_40_)  &  (~ i_39_)  &  (~ i_38_) ) ;
 assign wire1062 = ( _435 ) | ( (~ i_15_)  &  wire79  &  wire793 ) ;
 assign wire7498 = ( wire183 ) | ( wire1060 ) | ( wire1063 ) ;
 assign n_n1489 = ( wire1062 ) | ( wire7498 ) | ( _440 ) | ( _441 ) ;
 assign n_n693 = ( i_36_  &  (~ i_38_)  &  (~ i_37_) ) ;
 assign wire6821 = ( i_40_  &  i_39_  &  i_11_ ) ;
 assign wire182 = ( (~ i_7_)  &  wire45  &  n_n693  &  wire6821 ) ;
 assign n_n1023 = ( (~ i_34_)  &  i_33_  &  i_35_ ) ;
 assign wire301 = ( n_n833  &  n_n668  &  n_n1023 ) | ( n_n668  &  wire371  &  n_n1023 ) ;
 assign wire574 = ( (~ i_9_)  &  (~ i_17_) ) | ( (~ i_9_)  &  (~ i_16_) ) | ( (~ i_17_)  &  (~ i_16_) ) ;
 assign wire474 = ( n_n968  &  wire7510  &  _10693 ) ;
 assign wire7512 = ( (~ i_32_)  &  i_33_  &  n_n998  &  n_n973 ) ;
 assign wire7517 = ( i_21_  &  i_22_  &  i_15_  &  _10704 ) ;
 assign wire575 = ( wire364  &  wire7512 ) | ( wire474  &  wire7517 ) ;
 assign n_n411 = ( i_23_  &  i_24_  &  i_22_ ) ;
 assign wire407 = ( (~ i_5_)  &  i_17_  &  i_16_  &  i_15_ ) ;
 assign wire39 = ( (~ i_12_)  &  i_11_ ) | ( i_12_  &  (~ i_11_) ) ;
 assign wire478 = ( i_9_  &  (~ i_5_)  &  i_11_  &  _9041 ) ;
 assign wire6798 = ( n_n1048  &  n_n1047  &  wire400 ) ;
 assign n_n1372 = ( wire6798  &  _9291 ) | ( n_n955  &  wire6798  &  _9041 ) ;
 assign wire42 = ( i_9_  &  (~ i_5_)  &  i_12_ ) | ( i_9_  &  (~ i_5_)  &  i_11_ ) ;
 assign wire1834 = ( i_9_  &  (~ i_5_)  &  i_11_  &  i_19_ ) ;
 assign wire57 = ( wire1834 ) | ( i_18_  &  wire42 ) ;
 assign wire84 = ( n_n1055  &  n_n1048  &  n_n1047 ) ;
 assign wire416 = ( n_n1048  &  n_n1047  &  _9306 ) ;
 assign wire512 = ( n_n1074  &  wire48  &  wire6731  &  n_n978 ) ;
 assign wire317 = ( i_9_  &  (~ i_5_) ) ;
 assign wire579 = ( (~ i_12_)  &  i_11_  &  i_15_  &  wire317 ) | ( i_12_  &  (~ i_11_)  &  i_15_  &  wire317 ) ;
 assign n_n949 = ( (~ i_5_)  &  i_11_  &  i_15_ ) ;
 assign wire7128 = ( i_24_  &  i_21_  &  i_22_ ) ;
 assign n_n937 = ( n_n1074  &  n_n949  &  wire7128 ) ;
 assign wire473 = ( n_n985  &  n_n1023  &  n_n1064  &  wire7124 ) ;
 assign wire739 = ( wire484 ) | ( i_18_  &  wire36 ) ;
 assign n_n1374 = ( i_19_  &  wire473  &  wire739 ) ;
 assign wire120 = ( i_40_  &  i_39_  &  i_38_ ) | ( (~ i_40_)  &  (~ i_39_)  &  (~ i_38_) ) ;
 assign n_n1001 = ( i_39_  &  i_38_  &  (~ i_37_) ) ;
 assign n_n945 = ( i_24_  &  (~ i_32_)  &  i_33_ ) ;
 assign wire6789 = ( i_22_  &  (~ i_34_)  &  (~ i_36_)  &  i_35_ ) ;
 assign wire7133 = ( i_23_  &  i_21_ ) ;
 assign wire333 = ( n_n1001  &  n_n945  &  wire6789  &  wire7133 ) ;
 assign wire6907 = ( (~ i_36_)  &  i_35_  &  i_37_ ) ;
 assign wire386 = ( (~ i_36_)  &  i_35_  &  i_37_  &  _9425 ) ;
 assign n_n947 = ( (~ i_5_)  &  i_12_  &  i_15_ ) ;
 assign wire583 = ( n_n1074  &  n_n949  &  wire7128 ) | ( n_n1074  &  wire7128  &  n_n947 ) ;
 assign wire581 = ( (~ i_5_)  &  i_12_  &  i_15_ ) | ( (~ i_5_)  &  i_11_  &  i_15_ ) ;
 assign wire7531 = ( i_40_  &  i_39_  &  i_12_  &  (~ i_11_) ) ;
 assign wire146 = ( wire45  &  n_n693  &  wire7531 ) ;
 assign n_n698 = ( i_35_  &  (~ i_38_)  &  i_37_ ) ;
 assign n_n1056 = ( (~ i_34_)  &  i_33_  &  i_36_ ) ;
 assign wire7626 = ( (~ i_7_)  &  i_11_  &  (~ i_32_) ) ;
 assign wire131 = ( wire325  &  n_n1056  &  wire7626 ) ;
 assign wire402 = ( i_40_  &  i_36_  &  (~ i_35_)  &  i_38_ ) ;
 assign wire495 = ( i_40_  &  i_39_  &  (~ i_37_) ) ;
 assign n_n334 = ( i_13_  &  wire315  &  wire76 ) ;
 assign wire619 = ( i_40_  &  i_39_  &  n_n1073 ) | ( i_39_  &  (~ i_38_)  &  n_n1073 ) | ( (~ i_40_)  &  (~ i_39_)  &  i_38_  &  n_n1073 ) ;
 assign wire882 = ( wire888  &  wire7640 ) | ( n_n1066  &  n_n989  &  wire7640 ) ;
 assign wire7643 = ( wire321  &  wire506 ) | ( wire106  &  wire7641 ) ;
 assign wire7649 = ( i_40_  &  (~ i_38_)  &  n_n1074  &  wire6731 ) ;
 assign wire7650 = ( wire7304  &  wire7305 ) | ( wire433  &  wire7646 ) ;
 assign n_n866 = ( i_40_  &  (~ i_38_)  &  i_37_ ) ;
 assign wire849 = ( wire855  &  _10946 ) | ( _218  &  _10946 ) | ( _219  &  _10946 ) ;
 assign wire7669 = ( wire7666 ) | ( wire7667 ) | ( n_n515  &  wire92 ) ;
 assign wire7674 = ( wire7663 ) | ( wire7664 ) | ( wire7673 ) ;
 assign wire316 = ( i_38_  &  (~ i_37_) ) ;
 assign n_n848 = ( i_21_  &  i_22_  &  i_15_ ) ;
 assign wire587 = ( n_n853  &  n_n945  &  n_n848 ) | ( n_n850  &  n_n945  &  n_n848 ) ;
 assign wire94 = ( i_40_  &  (~ i_34_)  &  (~ i_36_)  &  i_35_ ) ;
 assign wire106 = ( n_n853  &  n_n945  &  n_n848 ) | ( n_n850  &  n_n945  &  n_n848 ) ;
 assign wire7679 = ( i_40_  &  i_15_  &  n_n945  &  wire6789 ) ;
 assign wire586 = ( wire94  &  wire106 ) | ( wire44  &  wire7679 ) ;
 assign n_n1197 = ( wire294 ) | ( wire295 ) | ( wire297 ) | ( wire7715 ) ;
 assign n_n1203 = ( _148 ) | ( _149 ) | ( wire6739  &  _11060 ) ;
 assign n_n1202 = ( wire271 ) | ( _145 ) | ( wire6739  &  _11064 ) ;
 assign wire7737 = ( wire7734 ) | ( n_n1055  &  n_n998  &  _11066 ) ;
 assign wire7738 = ( wire260 ) | ( wire261 ) | ( _11076 ) ;
 assign wire202 = ( i_28_ ) | ( i_29_ ) ;
 assign n_n462 = ( i_40_  &  (~ i_39_)  &  (~ i_36_)  &  i_38_ ) ;
 assign wire406 = ( (~ i_5_)  &  n_n462 ) ;
 assign n_n1237 = ( wire7774 ) | ( wire211 ) | ( wire213 ) | ( _86 ) ;
 assign n_n1239 = ( wire203 ) | ( wire7784 ) | ( wire7785 ) | ( wire7786 ) ;
 assign n_n775 = ( (~ i_34_)  &  (~ i_36_)  &  (~ i_35_)  &  _9420 ) ;
 assign wire400 = ( i_40_  &  i_39_  &  i_38_  &  (~ i_37_) ) ;
 assign n_n785 = ( (~ i_34_)  &  (~ i_36_)  &  (~ i_35_)  &  wire400 ) ;
 assign wire129 = ( wire48  &  n_n428  &  n_n427  &  wire706 ) ;
 assign wire7816 = ( i_40_  &  i_23_  &  (~ i_38_)  &  i_37_ ) ;
 assign n_n1242 = ( wire129 ) | ( _53 ) | ( _54 ) ;
 assign wire469 = ( i_9_  &  (~ i_7_)  &  (~ i_5_)  &  i_12_ ) ;
 assign n_n528 = ( i_40_  &  (~ i_39_)  &  (~ i_37_) ) ;
 assign n_n888 = ( (~ i_34_)  &  i_35_  &  (~ i_37_) ) ;
 assign wire315 = ( (~ i_7_)  &  (~ i_5_)  &  (~ i_12_)  &  (~ i_11_) ) ;
 assign n_n313 = ( i_13_  &  wire50  &  wire315 ) ;
 assign wire6887 = ( i_40_  &  (~ i_36_)  &  (~ i_38_) ) ;
 assign wire227 = ( n_n330  &  n_n1066  &  n_n989  &  wire6887 ) ;
 assign wire594 = ( i_40_  &  (~ i_38_)  &  i_37_ ) | ( i_39_  &  i_38_  &  (~ i_37_) ) ;
 assign wire869 = ( n_n979  &  wire594  &  n_n700  &  wire7276 ) ;
 assign wire7654 = ( wire873 ) | ( _195 ) | ( _196 ) ;
 assign wire68 = ( i_40_  &  (~ i_38_) ) | ( i_39_  &  (~ i_37_) ) ;
 assign wire504 = ( n_n793  &  n_n1047  &  wire78  &  wire6858 ) ;
 assign n_n960 = ( i_39_  &  i_38_ ) ;
 assign wire367 = ( i_12_  &  i_15_  &  n_n793 ) ;
 assign wire479 = ( n_n1048  &  n_n1047  &  wire6859 ) ;
 assign wire430 = ( n_n793  &  n_n1047  &  wire86  &  wire6850 ) ;
 assign wire78 = ( i_12_  &  i_15_ ) ;
 assign wire6858 = ( (~ i_16_)  &  (~ i_32_)  &  (~ i_31_)  &  i_33_ ) ;
 assign wire957 = ( wire68  &  wire504 ) ;
 assign wire7577 = ( wire479  &  wire368 ) | ( wire432  &  wire7576 ) ;
 assign wire7578 = ( wire430  &  wire837 ) | ( i_39_  &  (~ i_37_)  &  wire430 ) ;
 assign n_n1283 = ( wire174 ) | ( wire957 ) | ( wire7577 ) | ( wire7578 ) ;
 assign wire176 = ( (~ i_22_)  &  wire50  &  wire87  &  n_n833 ) ;
 assign wire7145 = ( i_40_  &  i_39_  &  (~ i_36_)  &  (~ i_38_) ) ;
 assign wire395 = ( wire80  &  wire7145 ) ;
 assign wire598 = ( wire50  &  wire82 ) | ( wire50  &  wire87 ) ;
 assign wire596 = ( (~ i_24_)  &  wire50  &  wire82 ) | ( (~ i_24_)  &  wire50  &  wire87 ) ;
 assign wire983 = ( (~ i_40_)  &  (~ i_39_)  &  (~ i_36_)  &  (~ i_38_) ) ;
 assign wire595 = ( n_n926 ) | ( wire983 ) ;
 assign wire7559 = ( wire176 ) | ( _334 ) | ( _335 ) ;
 assign wire7560 = ( n_n760  &  wire595 ) | ( wire598  &  wire7558 ) ;
 assign n_n1280 = ( wire7559 ) | ( wire7560 ) | ( n_n833  &  wire596 ) ;
 assign n_n1064 = ( i_40_  &  (~ i_39_) ) ;
 assign n_n525 = ( (~ i_13_)  &  wire50  &  wire315 ) ;
 assign wire464 = ( (~ i_3_)  &  (~ i_1_)  &  i_2_  &  i_0_ ) ;
 assign wire148 = ( (~ i_7_)  &  wire80  &  n_n1052  &  wire464 ) ;
 assign wire329 = ( (~ i_21_)  &  i_15_  &  n_n850 ) ;
 assign wire357 = ( (~ i_40_)  &  (~ i_39_)  &  n_n1009 ) ;
 assign wire408 = ( i_13_  &  wire315 ) ;
 assign wire441 = ( i_40_  &  (~ i_39_)  &  i_38_  &  i_37_ ) ;
 assign n_n1073 = ( (~ i_36_)  &  (~ i_35_)  &  (~ i_37_) ) ;
 assign n_n843 = ( (~ i_1_)  &  i_2_  &  i_0_ ) ;
 assign wire542 = ( n_n966  &  n_n842  &  n_n1073  &  n_n843 ) ;
 assign n_n764 = ( (~ i_22_)  &  wire50  &  wire82 ) ;
 assign wire600 = ( (~ i_21_)  &  i_15_  &  n_n853 ) | ( (~ i_21_)  &  i_15_  &  n_n850 ) ;
 assign wire7570 = ( wire973 ) | ( wire7566 ) | ( (~ i_38_)  &  wire542 ) ;
 assign wire7571 = ( wire7565 ) | ( wire7568 ) | ( i_40_  &  wire148 ) ;
 assign wire7574 = ( wire962 ) | ( wire964 ) | ( wire395  &  wire600 ) ;
 assign n_n799 = ( (~ i_40_)  &  i_39_  &  (~ i_38_) ) ;
 assign wire366 = ( (~ i_36_)  &  (~ i_35_)  &  i_37_  &  _9322 ) ;
 assign wire662 = ( wire46  &  wire43 ) | ( wire53  &  wire7772 ) ;
 assign wire7774 = ( wire208 ) | ( wire209 ) | ( wire210 ) ;
 assign wire203 = ( i_40_  &  wire206 ) | ( i_40_  &  wire207 ) ;
 assign wire7784 = ( wire198 ) | ( wire199 ) ;
 assign wire7785 = ( wire201 ) | ( (~ i_13_)  &  wire45  &  wire506 ) ;
 assign wire7786 = ( wire205 ) | ( n_n1055  &  n_n1047  &  wire463 ) ;
 assign n_n710 = ( (~ i_4_)  &  (~ i_1_)  &  i_0_ ) ;
 assign n_n715 = ( (~ i_34_)  &  i_35_  &  i_37_ ) ;
 assign wire602 = ( i_40_  &  (~ i_38_)  &  i_37_ ) | ( i_39_  &  i_38_  &  (~ i_37_) ) | ( (~ i_39_)  &  (~ i_38_)  &  (~ i_37_) ) ;
 assign wire7799 = ( n_n2581 ) | ( wire167 ) | ( wire170 ) ;
 assign wire7800 = ( wire165 ) | ( wire169 ) | ( wire171 ) ;
 assign n_n1235 = ( wire7799 ) | ( wire7800 ) | ( _46 ) ;
 assign wire420 = ( (~ i_7_)  &  (~ i_5_)  &  (~ i_15_) ) ;
 assign wire160 = ( wire45  &  _11278 ) ;
 assign wire7809 = ( (~ i_32_)  &  i_31_  &  (~ i_34_)  &  i_33_ ) ;
 assign wire607 = ( i_12_  &  (~ i_18_) ) | ( i_11_  &  (~ i_18_) ) | ( i_11_  &  (~ i_19_) ) ;
 assign n_n1094 = ( _1075 ) | ( _1076 ) | ( wire512  &  _9433 ) ;
 assign n_n2837 = ( (~ i_7_)  &  i_3_  &  wire80  &  n_n926 ) ;
 assign n_n1958 = ( (~ i_7_)  &  i_4_  &  wire80  &  n_n833 ) ;
 assign n_n1956 = ( (~ i_7_)  &  i_3_  &  wire80  &  n_n833 ) ;
 assign n_n1957 = ( (~ i_7_)  &  i_1_  &  wire80  &  n_n833 ) ;
 assign n_n964 = ( (~ i_36_)  &  (~ i_35_) ) ;
 assign n_n993 = ( (~ i_36_)  &  (~ i_35_)  &  (~ i_38_) ) ;
 assign wire81 = ( (~ i_38_)  &  i_37_ ) ;
 assign wire382 = ( (~ i_32_)  &  (~ i_31_) ) ;
 assign wire86 = ( i_11_  &  i_15_ ) ;
 assign n_n642 = ( i_17_  &  (~ i_32_)  &  i_33_ ) ;
 assign n_n1015 = ( i_39_  &  (~ i_38_) ) ;
 assign n_n559 = ( n_n853  &  n_n945  &  n_n848 ) ;
 assign wire320 = ( (~ i_31_)  &  (~ i_34_)  &  i_33_  &  (~ i_35_) ) ;
 assign n_n535 = ( i_16_  &  wire87  &  wire320 ) ;
 assign wire7405 = ( (~ i_24_)  &  (~ i_32_)  &  i_33_ ) ;
 assign wire359 = ( i_40_  &  (~ i_39_)  &  n_n985 ) ;
 assign n_n952 = ( i_40_  &  (~ i_39_)  &  n_n985  &  n_n1023 ) ;
 assign n_n935 = ( n_n1074  &  wire7128  &  n_n947 ) ;
 assign n_n329 = ( n_n330  &  n_n1066  &  n_n989 ) ;
 assign n_n527 = ( (~ i_7_)  &  (~ i_5_)  &  (~ i_11_) ) ;
 assign n_n688 = ( (~ i_39_)  &  (~ i_36_)  &  i_38_ ) ;
 assign n_n700 = ( (~ i_15_)  &  (~ i_32_)  &  i_33_ ) ;
 assign n_n492 = ( (~ i_9_)  &  (~ i_5_)  &  i_11_ ) ;
 assign wire100 = ( i_38_  &  i_37_ ) ;
 assign n_n1065 = ( i_36_  &  i_38_  &  i_37_ ) ;
 assign n_n488 = ( (~ i_9_)  &  (~ i_5_)  &  i_12_ ) ;
 assign n_n453 = ( i_3_  &  i_0_  &  (~ i_32_) ) ;
 assign wire77 = ( (~ i_32_)  &  i_33_  &  n_n998 ) ;
 assign wire378 = ( (~ i_5_)  &  (~ i_15_) ) ;
 assign n_n884 = ( (~ i_5_)  &  (~ i_13_)  &  (~ i_15_) ) ;
 assign n_n928 = ( i_9_  &  (~ i_5_)  &  (~ i_11_) ) ;
 assign n_n951 = ( i_9_  &  (~ i_5_)  &  i_12_ ) ;
 assign n_n860 = ( i_9_  &  (~ i_7_)  &  (~ i_5_) ) ;
 assign n_n560 = ( (~ i_39_)  &  (~ i_38_)  &  n_n1012 ) ;
 assign wire76 = ( (~ i_32_)  &  (~ i_31_)  &  (~ i_34_)  &  i_33_ ) ;
 assign n_n484 = ( (~ i_16_)  &  i_15_  &  n_n492  &  wire76 ) ;
 assign wire60 = ( i_40_  &  (~ i_39_)  &  (~ i_38_)  &  i_37_ ) | ( (~ i_40_)  &  (~ i_39_)  &  (~ i_38_)  &  (~ i_37_) ) ;
 assign wire401 = ( i_40_  &  (~ i_36_)  &  (~ i_35_)  &  (~ i_38_) ) ;
 assign wire465 = ( i_39_  &  (~ i_36_)  &  (~ i_35_)  &  (~ i_37_) ) ;
 assign wire103 = ( wire401 ) | ( wire465 ) ;
 assign n_n791 = ( (~ i_21_)  &  (~ i_32_)  &  i_33_ ) ;
 assign wire531 = ( n_n979  &  n_n949  &  n_n791 ) ;
 assign wire352 = ( (~ i_16_)  &  i_15_ ) ;
 assign wire7414 = ( (~ i_17_)  &  i_15_ ) ;
 assign wire611 = ( n_n492  &  wire76  &  wire352 ) | ( n_n492  &  wire76  &  wire7414 ) ;
 assign wire1179 = ( wire611  &  wire7415 ) ;
 assign wire1181 = ( n_n985  &  wire467  &  wire7121 ) | ( n_n985  &  wire468  &  wire7121 ) ;
 assign wire1183 = ( _524 ) | ( _525 ) ;
 assign wire7417 = ( wire1182 ) | ( (~ wire37)  &  n_n947  &  wire7416 ) ;
 assign wire6850 = ( (~ i_16_)  &  (~ i_32_)  &  (~ i_31_)  &  i_33_ ) ;
 assign wire613 = ( i_40_  &  (~ i_34_)  &  (~ i_36_)  &  i_35_ ) | ( i_40_  &  (~ i_34_)  &  i_36_  &  (~ i_35_) ) ;
 assign wire271 = ( i_40_  &  (~ i_38_)  &  n_n1074  &  n_n970 ) ;
 assign n_n777 = ( i_11_  &  i_15_  &  n_n793  &  wire6850 ) ;
 assign n_n781 = ( (~ i_17_)  &  (~ i_16_)  &  n_n1048  &  wire87 ) ;
 assign wire6851 = ( (~ i_40_)  &  i_38_  &  (~ i_37_) ) ;
 assign wire64 = ( n_n1055  &  n_n1047 ) | ( n_n1047  &  wire6851 ) ;
 assign wire321 = ( (~ i_31_)  &  wire45 ) ;
 assign wire1786 = ( (~ i_9_)  &  (~ i_7_)  &  (~ i_5_)  &  i_12_ ) ;
 assign wire614 = ( wire1786 ) | ( (~ i_18_)  &  wire35 ) ;
 assign n_n1057 = ( (~ i_3_)  &  i_4_  &  (~ i_32_) ) ;
 assign wire61 = ( i_12_ ) | ( i_11_ ) ;
 assign wire7390 = ( (~ i_22_)  &  (~ i_32_)  &  i_33_ ) ;
 assign n_n162 = ( n_n979  &  n_n947  &  wire7390 ) ;
 assign n_n801 = ( (~ i_7_)  &  (~ i_5_)  &  (~ i_28_) ) ;
 assign n_n428 = ( i_24_  &  i_22_  &  (~ i_32_) ) ;
 assign n_n427 = ( i_40_  &  i_39_  &  n_n1009  &  n_n1023 ) ;
 assign wire7399 = ( (~ i_24_)  &  (~ i_32_)  &  i_33_ ) ;
 assign n_n907 = ( (~ i_5_)  &  (~ i_12_)  &  (~ i_11_) ) ;
 assign wire6716 = ( (~ i_13_)  &  (~ i_32_)  &  i_33_ ) ;
 assign n_n905 = ( n_n979  &  n_n907  &  wire6716 ) ;
 assign wire1204 = ( n_n1052  &  n_n1057  &  n_n1053  &  wire7388 ) ;
 assign wire1205 = ( _547 ) | ( n_n947  &  n_n791  &  wire642 ) ;
 assign wire1206 = ( n_n979  &  n_n469  &  n_n947  &  wire7347 ) ;
 assign wire7392 = ( wire1208 ) | ( (~ i_5_)  &  n_n462  &  wire468 ) ;
 assign wire1196 = ( n_n1061  &  wire69  &  _10434 ) | ( n_n1061  &  _10434  &  _10435 ) ;
 assign wire1197 = ( n_n979  &  n_n947  &  wire7399  &  wire660 ) ;
 assign wire1198 = ( n_n843  &  n_n1057  &  n_n1053  &  n_n836 ) ;
 assign wire7403 = ( wire154 ) | ( wire1199 ) | ( wire1200 ) ;
 assign wire7122 = ( (~ i_30_)  &  (~ i_32_)  &  (~ i_31_) ) ;
 assign wire467 = ( i_28_  &  (~ i_29_)  &  n_n1066  &  wire7122 ) ;
 assign n_n164 = ( n_n979  &  n_n949  &  wire7406 ) ;
 assign wire1192 = ( n_n979  &  n_n947  &  n_n791 ) ;
 assign wire616 = ( wire531 ) | ( n_n162 ) | ( n_n164 ) | ( wire1192 ) ;
 assign wire615 = ( i_40_  &  (~ i_39_)  &  (~ i_38_) ) | ( i_39_  &  i_38_  &  (~ i_37_) ) | ( (~ i_39_)  &  (~ i_38_)  &  (~ i_37_) ) ;
 assign n_n475 = ( (~ i_16_)  &  i_15_  &  n_n488  &  wire76 ) ;
 assign wire7406 = ( (~ i_22_)  &  (~ i_32_)  &  i_33_ ) ;
 assign wire696 = ( n_n484 ) | ( wire113 ) | ( wire1173 ) | ( wire1174 ) ;
 assign wire7427 = ( wire7420  &  wire7421 ) | ( wire695  &  wire7423 ) ;
 assign wire113 = ( n_n488  &  wire76  &  wire352 ) | ( n_n488  &  wire76  &  wire7414 ) ;
 assign wire617 = ( wire401 ) | ( wire465 ) ;
 assign wire506 = ( i_40_  &  i_39_  &  n_n1052  &  wire315 ) ;
 assign wire433 = ( n_n945  &  wire6789  &  n_n860 ) ;
 assign wire7648 = ( i_15_  &  wire491 ) ;
 assign wire7330 = ( (~ i_40_)  &  i_39_  &  (~ i_37_) ) ;
 assign n_n2439 = ( n_n1002  &  n_n861  &  wire7330 ) ;
 assign wire624 = ( (~ i_34_)  &  i_36_  &  i_37_ ) | ( (~ i_34_)  &  i_35_  &  i_37_ ) ;
 assign wire421 = ( (~ i_32_)  &  i_33_  &  (~ i_36_)  &  (~ i_35_) ) ;
 assign n_n1053 = ( i_34_  &  i_33_  &  (~ i_35_) ) ;
 assign wire627 = ( (~ i_9_)  &  (~ i_5_)  &  i_12_ ) | ( (~ i_9_)  &  (~ i_5_)  &  i_11_ ) ;
 assign wire294 = ( (~ i_36_)  &  wire45  &  wire627  &  wire7707 ) ;
 assign wire295 = ( (~ wire37)  &  n_n947  &  wire400  &  wire421 ) ;
 assign wire297 = ( _175 ) | ( _176 ) | ( _177 ) ;
 assign wire7715 = ( wire298 ) | ( _172 ) | ( _173 ) ;
 assign wire36 = ( (~ i_5_)  &  i_12_  &  i_15_ ) | ( (~ i_5_)  &  i_11_  &  i_15_ ) ;
 assign wire451 = ( n_n1009  &  n_n1021  &  n_n874  &  wire7686 ) ;
 assign wire454 = ( n_n979  &  wire81  &  n_n791  &  wire36 ) ;
 assign wire7692 = ( wire455 ) | ( _119 ) | ( _120 ) ;
 assign wire633 = ( (~ i_5_)  &  i_12_  &  i_15_ ) | ( (~ i_5_)  &  i_11_  &  i_15_ ) ;
 assign wire446 = ( _110 ) | ( _111 ) | ( _112 ) ;
 assign wire7394 = ( (~ i_40_)  &  i_10_  &  i_27_  &  (~ i_39_) ) ;
 assign wire154 = ( wire45  &  n_n1061  &  wire7394 ) ;
 assign wire635 = ( (~ i_9_)  &  (~ i_5_)  &  i_12_ ) | ( (~ i_9_)  &  (~ i_5_)  &  (~ i_15_) ) ;
 assign wire65 = ( i_39_  &  i_38_  &  (~ i_37_) ) | ( (~ i_39_)  &  (~ i_38_)  &  (~ i_37_) ) ;
 assign wire638 = ( i_40_  &  i_39_  &  (~ i_37_) ) | ( i_40_  &  (~ i_38_)  &  (~ i_37_) ) | ( i_39_  &  (~ i_38_)  &  (~ i_37_) ) ;
 assign wire637 = ( n_n1055  &  n_n1047 ) | ( n_n1047  &  wire638 ) ;
 assign wire1913 = ( _1215 ) | ( _1216 ) | ( _1217 ) ;
 assign wire6734 = ( wire1910 ) | ( wire1911 ) | ( wire1914 ) ;
 assign n_n1135 = ( wire1913 ) | ( wire6734 ) | ( _1218 ) | ( _1219 ) ;
 assign n_n582 = ( (~ i_36_)  &  i_38_  &  i_37_ ) ;
 assign n_n771 = ( i_12_  &  i_15_  &  n_n793  &  wire6858 ) ;
 assign wire368 = ( i_11_  &  i_15_  &  n_n793 ) ;
 assign wire6859 = ( i_39_  &  (~ i_17_)  &  i_38_ ) ;
 assign wire369 = ( wire50  &  wire82 ) ;
 assign wire7389 = ( i_30_  &  (~ i_28_)  &  i_29_ ) ;
 assign wire468 = ( (~ i_31_)  &  wire45  &  wire7389 ) ;
 assign wire6976 = ( (~ i_39_)  &  (~ i_19_)  &  (~ i_38_)  &  i_37_ ) ;
 assign wire83 = ( n_n979  &  n_n791  &  wire6976 ) ;
 assign wire356 = ( (~ i_40_)  &  (~ i_39_)  &  i_38_  &  _10830 ) ;
 assign wire643 = ( i_12_  &  i_15_  &  n_n793 ) | ( i_11_  &  i_15_  &  n_n793 ) ;
 assign wire950 = ( n_n979  &  n_n1055  &  n_n783 ) | ( n_n979  &  n_n1055  &  n_n790 ) ;
 assign wire952 = ( n_n1055  &  n_n1047  &  n_n777 ) | ( n_n1055  &  n_n1047  &  n_n771 ) ;
 assign wire7582 = ( n_n793  &  wire84  &  _9411 ) | ( n_n793  &  wire84  &  _9416 ) ;
 assign wire7583 = ( n_n777  &  wire356 ) | ( wire83  &  wire643 ) ;
 assign n_n1285 = ( wire950 ) | ( wire952 ) | ( wire7582 ) | ( wire7583 ) ;
 assign wire486 = ( i_15_  &  wire35 ) ;
 assign wire648 = ( (~ wire37)  &  n_n1048  &  wire82 ) | ( (~ wire37)  &  n_n1048  &  wire87 ) ;
 assign wire646 = ( n_n1055  &  n_n1047 ) | ( n_n1072  &  n_n1073 ) ;
 assign n_n923 = ( i_39_  &  (~ i_36_)  &  i_38_ ) ;
 assign wire286 = ( wire45  &  n_n488  &  n_n923  &  wire7717 ) ;
 assign wire287 = ( _165 ) | ( n_n791  &  wire652  &  wire650 ) ;
 assign wire288 = ( n_n979  &  n_n969  &  n_n949  &  n_n791 ) ;
 assign wire289 = ( n_n979  &  n_n949  &  n_n1001  &  wire7406 ) ;
 assign n_n1068 = ( i_17_  &  i_16_  &  i_15_ ) ;
 assign wire303 = ( i_39_  &  i_38_  &  n_n1074  &  n_n968 ) ;
 assign wire73 = ( (~ i_14_) ) | ( (~ i_12_) ) | ( (~ i_11_) ) ;
 assign wire520 = ( n_n1014  &  n_n1009  &  n_n874  &  (~ wire73) ) ;
 assign wire655 = ( (~ i_9_)  &  (~ i_5_)  &  i_12_ ) | ( (~ i_9_)  &  (~ i_5_)  &  i_11_ ) ;
 assign wire835 = ( (~ i_7_)  &  wire80  &  n_n926 ) | ( (~ i_7_)  &  wire80  &  n_n833 ) ;
 assign wire336 = ( i_40_  &  i_39_  &  n_n966  &  n_n993 ) ;
 assign n_n458 = ( i_2_  &  i_0_  &  (~ i_32_) ) ;
 assign n_n643 = ( i_16_  &  (~ i_32_)  &  i_33_ ) ;
 assign wire1681 = ( (~ i_24_)  &  wire50  &  wire87  &  wire6945 ) ;
 assign wire1682 = ( (~ i_24_)  &  wire50  &  wire82  &  wire371 ) ;
 assign n_n836 = ( (~ i_39_)  &  (~ i_36_)  &  (~ i_38_) ) ;
 assign wire660 = ( i_40_  &  (~ i_39_)  &  (~ i_38_) ) | ( i_39_  &  i_38_  &  (~ i_37_) ) ;
 assign wire43 = ( (~ i_7_)  &  (~ i_5_)  &  i_28_  &  i_29_ ) | ( (~ i_7_)  &  (~ i_5_)  &  (~ i_28_)  &  (~ i_29_) ) ;
 assign wire53 = ( (~ i_30_)  &  i_29_ ) | ( i_30_  &  (~ i_29_) ) ;
 assign wire7772 = ( (~ i_7_)  &  (~ i_5_)  &  (~ i_32_)  &  i_33_ ) ;
 assign wire351 = ( i_17_  &  i_16_  &  (~ i_32_)  &  i_33_ ) ;
 assign wire463 = ( (~ i_14_)  &  wire87  &  wire351 ) ;
 assign wire666 = ( (~ i_40_)  &  i_38_ ) | ( i_39_  &  i_38_ ) ;
 assign wire665 = ( (~ i_40_)  &  (~ i_38_) ) | ( i_39_  &  (~ i_38_) ) ;
 assign wire664 = ( (~ i_5_)  &  (~ i_38_)  &  i_37_ ) | ( i_35_  &  (~ i_38_)  &  i_37_ ) ;
 assign wire153 = ( n_n1074  &  n_n864  &  n_n977 ) ;
 assign wire6773 = ( (~ i_10_)  &  (~ i_39_)  &  i_38_  &  (~ i_37_) ) ;
 assign wire184 = ( (~ i_32_)  &  i_33_  &  n_n991  &  wire6773 ) ;
 assign wire6774 = ( (~ i_27_)  &  (~ i_39_)  &  i_38_  &  (~ i_37_) ) ;
 assign wire187 = ( (~ i_32_)  &  i_33_  &  n_n991  &  wire6774 ) ;
 assign wire458 = ( i_40_  &  (~ i_5_)  &  (~ i_39_)  &  i_38_ ) ;
 assign wire669 = ( (~ i_30_)  &  i_29_ ) | ( i_28_  &  i_29_ ) | ( i_30_  &  (~ i_29_) ) ;
 assign wire668 = ( (~ i_30_)  &  i_29_ ) | ( i_28_  &  i_29_ ) | ( i_30_  &  (~ i_29_) ) | ( (~ i_28_)  &  (~ i_29_) ) ;
 assign wire327 = ( (~ i_36_)  &  (~ i_35_)  &  (~ i_37_)  &  _10233 ) ;
 assign wire670 = ( i_9_  &  i_17_  &  i_15_ ) | ( i_9_  &  i_16_  &  i_15_ ) | ( i_17_  &  i_16_  &  i_15_ ) ;
 assign wire671 = ( i_39_  &  i_38_ ) | ( i_40_  &  (~ i_38_) ) | ( i_39_  &  (~ i_37_) ) ;
 assign wire672 = ( wire54 ) | ( wire371 ) ;
 assign wire529 = ( i_30_  &  i_29_  &  wire76  &  n_n801 ) ;
 assign wire370 = ( wire50  &  wire87 ) ;
 assign n_n918 = ( i_39_  &  (~ i_36_)  &  (~ i_38_) ) ;
 assign n_n556 = ( n_n850  &  n_n945  &  n_n848 ) ;
 assign n_n798 = ( (~ i_7_)  &  (~ i_5_)  &  i_28_ ) ;
 assign n_n859 = ( i_11_  &  i_18_  &  i_15_ ) ;
 assign wire674 = ( (~ i_9_)  &  (~ i_17_) ) | ( (~ i_9_)  &  (~ i_16_) ) | ( (~ i_17_)  &  (~ i_16_) ) ;
 assign wire403 = ( (~ i_40_)  &  (~ i_38_)  &  i_37_ ) ;
 assign wire677 = ( i_3_ ) | ( i_4_ ) | ( i_1_ ) | ( i_2_ ) ;
 assign wire1160 = ( (~ i_39_)  &  i_2_  &  (~ i_38_)  &  i_37_ ) ;
 assign wire676 = ( wire1160 ) | ( n_n1001  &  wire677 ) ;
 assign wire7397 = ( i_3_  &  i_0_ ) ;
 assign wire69 = ( n_n1066  &  _10436 ) | ( n_n1066  &  _10437 ) ;
 assign wire332 = ( i_4_  &  i_0_  &  wire45 ) ;
 assign wire681 = ( i_3_  &  i_0_  &  (~ i_32_) ) | ( i_2_  &  i_0_  &  (~ i_32_) ) ;
 assign wire679 = ( n_n1021  &  n_n862 ) | ( n_n1012  &  n_n960 ) ;
 assign wire678 = ( i_40_  &  i_39_  &  n_n1061 ) | ( i_40_  &  (~ i_39_)  &  n_n1065 ) ;
 assign wire7227 = ( i_0_  &  (~ i_32_)  &  i_33_  &  i_37_ ) ;
 assign wire7750 = ( (~ i_4_)  &  i_0_ ) | ( (~ i_1_)  &  i_0_ ) ;
 assign wire684 = ( (~ i_32_)  &  n_n1023  &  wire7397 ) | ( (~ i_32_)  &  n_n1023  &  wire7750 ) ;
 assign wire484 = ( i_9_  &  (~ i_5_)  &  i_12_  &  i_15_ ) ;
 assign wire1766 = ( (~ i_40_)  &  i_38_  &  n_n334  &  n_n1073 ) ;
 assign wire6868 = ( wire479  &  wire368 ) | ( wire366  &  wire535 ) ;
 assign wire6869 = ( wire430  &  wire6863 ) | ( wire303  &  wire6866 ) ;
 assign wire6870 = ( n_n334  &  n_n560 ) | ( wire430  &  wire837 ) ;
 assign n_n1091 = ( wire1766 ) | ( wire6868 ) | ( wire6869 ) | ( wire6870 ) ;
 assign n_n1113 = ( _554 ) | ( _555 ) ;
 assign wire244 = ( n_n330  &  n_n926  &  n_n1066  &  n_n989 ) ;
 assign wire688 = ( wire50  &  wire82 ) | ( wire50  &  wire87 ) ;
 assign wire6878 = ( wire175 ) | ( wire176 ) | ( wire244 ) | ( wire1758 ) ;
 assign wire6879 = ( wire6860 ) | ( wire6861 ) | ( wire6877 ) ;
 assign wire1751 = ( n_n979  &  n_n158  &  wire702  &  wire701 ) ;
 assign wire6886 = ( wire245 ) | ( n_n469  &  wire700 ) ;
 assign wire6894 = ( n_n1990 ) | ( wire227 ) | ( wire1741 ) | ( wire1742 ) ;
 assign wire711 = ( i_37_  &  n_n883  &  wire326 ) | ( (~ i_37_)  &  n_n1072  &  wire326 ) ;
 assign n_n1108 = ( n_n1971 ) | ( n_n1074  &  wire6897  &  wire711 ) ;
 assign wire689 = ( i_30_  &  (~ i_28_)  &  i_29_  &  wire47 ) | ( (~ i_30_)  &  i_28_  &  (~ i_29_)  &  wire47 ) ;
 assign wire6908 = ( i_24_  &  (~ i_22_) ) ;
 assign wire132 = ( n_n1074  &  wire82  &  wire6908 ) | ( n_n1074  &  wire87  &  wire6908 ) ;
 assign wire690 = ( (~ wire37)  &  n_n1048  &  wire82 ) | ( (~ wire37)  &  n_n1048  &  wire87 ) ;
 assign n_n927 = ( i_16_  &  (~ i_32_)  &  (~ i_31_) ) ;
 assign n_n773 = ( (~ i_17_)  &  (~ i_16_)  &  n_n1048  &  wire82 ) ;
 assign wire337 = ( i_40_  &  i_39_  &  n_n985  &  wire80 ) ;
 assign wire344 = ( i_9_  &  (~ i_7_) ) ;
 assign wire693 = ( (~ i_14_) ) | ( (~ i_11_) ) ;
 assign wire692 = ( (~ i_12_)  &  n_n642 ) | ( (~ i_12_)  &  n_n643 ) | ( n_n642  &  wire693 ) | ( n_n643  &  wire693 ) ;
 assign wire1173 = ( (~ i_17_)  &  (~ i_16_)  &  n_n949  &  wire76 ) ;
 assign wire1174 = ( (~ i_17_)  &  i_15_  &  n_n492  &  wire76 ) ;
 assign wire695 = ( n_n492  &  wire76  &  wire352 ) | ( n_n488  &  wire76  &  wire352 ) ;
 assign wire1291 = ( i_30_  &  (~ i_7_)  &  (~ i_5_)  &  (~ i_29_) ) ;
 assign wire102 = ( wire43 ) | ( wire1291 ) ;
 assign wire697 = ( i_40_  &  (~ i_39_)  &  (~ i_38_)  &  i_37_ ) | ( i_40_  &  i_39_  &  (~ i_38_)  &  (~ i_37_) ) ;
 assign wire509 = ( i_40_  &  (~ i_39_)  &  n_n862 ) ;
 assign wire342 = ( i_40_  &  (~ i_39_)  &  (~ i_38_)  &  i_37_ ) ;
 assign wire380 = ( i_18_  &  wire36 ) ;
 assign wire702 = ( (~ i_40_)  &  i_39_  &  i_38_  &  (~ i_37_) ) | ( (~ i_40_)  &  (~ i_39_)  &  (~ i_38_)  &  (~ i_37_) ) ;
 assign wire701 = ( (~ i_7_)  &  (~ i_5_)  &  i_12_ ) | ( (~ i_7_)  &  (~ i_5_)  &  i_11_ ) ;
 assign wire6884 = ( (~ i_7_)  &  (~ i_5_)  &  (~ i_12_) ) ;
 assign wire700 = ( n_n1048  &  n_n1047  &  n_n527 ) | ( n_n1048  &  n_n1047  &  wire6884 ) ;
 assign wire6968 = ( (~ i_18_)  &  (~ i_21_)  &  (~ i_32_)  &  i_33_ ) ;
 assign n_n783 = ( i_12_  &  i_15_  &  n_n793  &  wire6968 ) ;
 assign wire7309 = ( (~ i_7_)  &  (~ i_34_)  &  i_33_ ) ;
 assign n_n550 = ( n_n1068  &  (~ wire73)  &  wire7309 ) ;
 assign wire855 = ( i_40_  &  (~ i_13_)  &  wire50  &  wire315 ) ;
 assign wire133 = ( i_9_  &  (~ i_7_)  &  (~ i_5_)  &  i_11_ ) ;
 assign wire706 = ( wire133 ) | ( i_18_  &  wire35 ) ;
 assign wire710 = ( wire54 ) | ( wire371 ) ;
 assign wire1749 = ( n_n1074  &  n_n883  &  n_n970  &  wire6828 ) ;
 assign wire1747 = ( n_n1074  &  n_n971  &  n_n1072  &  wire6828 ) ;
 assign wire383 = ( (~ i_36_)  &  (~ i_37_) ) ;
 assign wire429 = ( (~ i_7_)  &  i_2_  &  i_0_  &  _9527 ) ;
 assign n_n1577 = ( n_n1951 ) | ( n_n1108 ) | ( _567 ) | ( _10388 ) ;
 assign wire713 = ( (~ i_39_)  &  (~ i_36_)  &  i_38_ ) | ( i_39_  &  (~ i_36_)  &  (~ i_38_) ) | ( (~ i_36_)  &  i_38_  &  i_37_ ) | ( (~ i_36_)  &  (~ i_38_)  &  (~ i_37_) ) ;
 assign wire1099 = ( (~ i_40_)  &  (~ i_36_)  &  i_38_ ) ;
 assign wire7473 = ( (~ i_39_)  &  (~ i_36_)  &  i_38_ ) | ( (~ i_36_)  &  (~ i_38_)  &  (~ i_37_) ) ;
 assign wire7474 = ( i_39_  &  (~ i_36_)  &  (~ i_38_) ) | ( (~ i_36_)  &  i_38_  &  i_37_ ) ;
 assign wire718 = ( wire1099 ) | ( wire7473 ) | ( wire7474 ) ;
 assign wire717 = ( (~ i_9_)  &  (~ i_17_) ) | ( (~ i_9_)  &  (~ i_16_) ) | ( (~ i_17_)  &  (~ i_16_) ) ;
 assign wire139 = ( i_40_  &  i_38_  &  n_n979 ) | ( (~ i_38_)  &  i_37_  &  n_n979 ) ;
 assign wire1277 = ( i_17_  &  wire721  &  wire7308 ) | ( i_16_  &  wire721  &  wire7308 ) ;
 assign wire7311 = ( wire327  &  n_n550 ) | ( wire7304  &  wire7305 ) ;
 assign wire488 = ( (~ i_31_)  &  i_33_ ) ;
 assign wire723 = ( i_16_  &  wire82  &  wire320 ) | ( i_16_  &  wire87  &  wire320 ) ;
 assign wire7319 = ( wire1271 ) | ( n_n1008  &  wire411  &  n_n698 ) ;
 assign wire7320 = ( wire364  &  wire336 ) | ( n_n560  &  n_n550 ) ;
 assign wire7321 = ( n_n556  &  wire139 ) | ( n_n559  &  wire7317 ) | ( n_n556  &  wire7317 ) ;
 assign wire1269 = ( i_40_  &  (~ i_39_)  &  i_36_  &  (~ i_35_) ) ;
 assign wire724 = ( wire402 ) | ( wire1269 ) ;
 assign wire727 = ( i_18_  &  wire35 ) | ( n_n860  &  wire61 ) ;
 assign wire7124 = ( i_23_  &  i_24_  &  i_22_  &  (~ i_32_) ) ;
 assign wire925 = ( n_n1048  &  n_n973  &  n_n1073  &  wire420 ) ;
 assign wire926 = ( n_n1074  &  wire6897  &  wire402 ) | ( n_n1074  &  wire6897  &  wire930 ) ;
 assign wire927 = ( _297 ) | ( (~ i_40_)  &  i_39_  &  wire932 ) ;
 assign wire361 = ( (~ i_30_)  &  (~ i_32_)  &  (~ i_31_)  &  _9966 ) ;
 assign wire450 = ( i_9_  &  (~ i_14_) ) ;
 assign wire38 = ( i_17_  &  (~ i_32_)  &  i_33_ ) | ( i_16_  &  (~ i_32_)  &  i_33_ ) ;
 assign wire738 = ( (~ i_14_) ) | ( (~ i_12_) ) | ( (~ i_11_) ) ;
 assign wire737 = ( wire450  &  wire38 ) | ( wire351  &  wire738 ) ;
 assign wire740 = ( i_39_  &  i_38_  &  i_37_ ) | ( (~ i_39_)  &  (~ i_38_)  &  i_37_ ) | ( (~ i_39_)  &  i_38_  &  (~ i_37_) ) ;
 assign n_n1134 = ( wire1909 ) | ( _9119 ) | ( n_n967  &  wire758 ) ;
 assign wire1901 = ( n_n1074  &  n_n1073  &  wire743 ) ;
 assign wire1902 = ( (~ i_39_)  &  (~ i_38_)  &  n_n1074  &  n_n968 ) ;
 assign wire742 = ( wire363 ) | ( wire303 ) | ( wire1901 ) | ( wire1902 ) ;
 assign wire741 = ( i_37_  &  n_n973  &  n_n964 ) | ( (~ i_37_)  &  n_n967  &  n_n964 ) ;
 assign wire7191 = ( (~ i_7_)  &  i_33_ ) ;
 assign wire7201 = ( i_12_  &  i_16_  &  i_15_ ) ;
 assign wire124 = ( i_40_  &  (~ i_38_)  &  (~ i_37_) ) | ( i_39_  &  (~ i_38_)  &  (~ i_37_) ) ;
 assign wire744 = ( (~ i_24_)  &  wire50  &  wire82 ) | ( (~ i_24_)  &  wire50  &  wire87 ) ;
 assign wire535 = ( (~ i_30_)  &  (~ i_29_)  &  wire76  &  n_n798 ) ;
 assign wire749 = ( i_40_  &  (~ i_39_)  &  (~ i_37_) ) | ( (~ i_39_)  &  (~ i_38_)  &  (~ i_37_) ) ;
 assign wire748 = ( (~ n_n1014)  &  n_n985 ) | ( i_35_  &  wire749 ) ;
 assign wire6974 = ( (~ i_18_)  &  (~ i_21_)  &  (~ i_32_)  &  i_33_ ) ;
 assign n_n790 = ( i_11_  &  i_15_  &  n_n793  &  wire6974 ) ;
 assign wire166 = ( (~ i_12_) ) | ( (~ i_11_) ) | ( (~ i_15_) ) ;
 assign wire752 = ( n_n979  &  n_n861 ) | ( (~ i_40_)  &  n_n861  &  n_n991 ) ;
 assign wire7154 = ( (~ i_30_)  &  (~ i_28_)  &  (~ i_29_) ) ;
 assign wire140 = ( n_n976  &  wire382  &  wire458  &  wire7154 ) ;
 assign wire7146 = ( i_21_  &  i_22_ ) ;
 assign wire156 = ( wire80  &  wire7145  &  wire36  &  wire7146 ) ;
 assign wire494 = ( (~ i_7_)  &  (~ i_5_)  &  i_29_ ) ;
 assign wire758 = ( (~ i_34_)  &  wire6731  &  wire46 ) | ( i_34_  &  wire46  &  n_n1073 ) ;
 assign n_n765 = ( (~ i_21_)  &  i_15_  &  wire50  &  n_n853 ) ;
 assign wire761 = ( (~ i_36_)  &  i_38_  &  i_37_  &  n_n1008 ) | ( (~ i_36_)  &  (~ i_38_)  &  (~ i_37_)  &  n_n1008 ) ;
 assign wire763 = ( i_40_  &  (~ i_39_)  &  (~ i_36_)  &  i_37_ ) | ( i_40_  &  i_39_  &  (~ i_36_)  &  (~ i_37_) ) ;
 assign wire762 = ( wire78  &  wire320  &  n_n860 ) | ( wire86  &  wire320  &  n_n860 ) ;
 assign wire767 = ( i_40_  &  (~ i_39_)  &  (~ i_38_) ) | ( i_40_  &  (~ i_39_)  &  (~ i_37_) ) ;
 assign wire1661 = ( n_n777  &  wire64 ) | ( wire64  &  n_n771 ) ;
 assign wire1662 = ( (~ i_21_)  &  i_15_  &  n_n853  &  wire348 ) ;
 assign wire6970 = ( n_n793  &  wire84  &  _9411 ) | ( n_n793  &  wire84  &  _9416 ) ;
 assign wire6971 = ( n_n775  &  n_n773 ) | ( n_n783  &  wire6969 ) ;
 assign wire101 = ( (~ i_40_)  &  (~ i_39_)  &  n_n1052 ) ;
 assign wire772 = ( i_39_  &  i_38_ ) | ( i_40_  &  (~ i_38_) ) ;
 assign wire373 = ( (~ i_40_)  &  (~ i_38_) ) ;
 assign wire7367 = ( o_32_ ) | ( n_n2836 ) | ( n_n1993 ) ;
 assign wire7371 = ( n_n2837 ) | ( n_n1958 ) | ( _10392 ) ;
 assign n_n1575 = ( wire7367 ) | ( wire7371 ) | ( i_2_  &  wire835 ) ;
 assign wire775 = ( wire334  &  n_n969 ) | ( (~ i_36_)  &  wire334  &  n_n1014 ) ;
 assign wire7132 = ( (~ i_5_)  &  (~ i_14_) ) | ( (~ i_5_)  &  (~ i_12_) ) | ( (~ i_5_)  &  (~ i_11_) ) ;
 assign wire461 = ( n_n1066  &  wire7132  &  _9971 ) ;
 assign wire1487 = ( i_40_  &  i_39_  &  (~ i_36_)  &  i_38_ ) ;
 assign wire777 = ( n_n926 ) | ( wire1487 ) ;
 assign wire1489 = ( n_n1014  &  wire380  &  wire482 ) | ( n_n1014  &  wire482  &  wire7127 ) ;
 assign wire7129 = ( wire386  &  n_n935 ) | ( n_n937  &  wire775 ) | ( n_n935  &  wire775 ) ;
 assign wire7139 = ( n_n1374 ) | ( _805 ) | ( _808 ) | ( _809 ) ;
 assign wire7140 = ( wire7135 ) | ( wire7137 ) | ( wire473  &  wire7125 ) ;
 assign wire7375 = ( wire1749 ) | ( wire1213 ) | ( wire7373 ) | ( _1065 ) ;
 assign wire7200 = ( i_9_  &  i_11_  &  i_15_ ) ;
 assign wire779 = ( (~ i_40_)  &  i_39_  &  i_35_  &  i_38_ ) | ( i_40_  &  (~ i_39_)  &  (~ i_35_)  &  i_38_ ) ;
 assign wire782 = ( n_n998  &  n_n973 ) | ( n_n969  &  n_n888 ) ;
 assign wire67 = ( (~ i_14_) ) | ( (~ i_12_) ) ;
 assign wire7150 = ( i_40_  &  (~ i_14_) ) ;
 assign wire786 = ( n_n926  &  wire67 ) | ( n_n923  &  wire7150 ) ;
 assign wire787 = ( i_40_  &  (~ i_39_)  &  n_n985 ) | ( (~ i_40_)  &  (~ i_39_)  &  n_n1052 ) ;
 assign wire6950 = ( wire365  &  wire337 ) | ( (~ i_22_)  &  wire82  &  wire337 ) ;
 assign wire6951 = ( wire323  &  n_n765 ) | ( (~ i_23_)  &  wire323  &  wire369 ) ;
 assign wire6952 = ( wire504  &  wire671 ) | ( n_n764  &  wire787 ) ;
 assign n_n1580 = ( wire6950 ) | ( wire6951 ) | ( wire6952 ) ;
 assign wire788 = ( (~ i_40_)  &  (~ i_39_)  &  i_38_ ) | ( i_40_  &  i_39_  &  (~ i_38_) ) ;
 assign wire795 = ( (~ i_14_) ) | ( (~ i_12_) ) | ( (~ i_11_) ) | ( (~ i_15_) ) ;
 assign wire794 = ( i_39_ ) | ( i_38_ ) | ( (~ i_37_) ) ;
 assign wire826 = ( wire1570 ) | ( (~ wire61)  &  wire1571 ) | ( (~ wire61)  &  wire7058 ) ;
 assign wire7062 = ( wire1565 ) | ( wire1566 ) | ( wire1568 ) ;
 assign wire158 = ( wire325  &  n_n991  &  _9886 ) ;
 assign wire7176 = ( wire1430 ) | ( wire1452 ) | ( wire7160 ) | ( wire7161 ) ;
 assign wire6956 = ( wire329  &  wire337 ) | ( (~ i_22_)  &  wire87  &  wire337 ) ;
 assign wire6957 = ( _1021 ) | ( n_n793  &  wire479  &  _9369 ) ;
 assign wire6958 = ( n_n761  &  wire830 ) | ( n_n760  &  wire829 ) ;
 assign wire803 = ( n_n1074  &  wire326 ) | ( wire490  &  n_n700 ) ;
 assign wire806 = ( (~ i_12_)  &  (~ i_11_) ) | ( (~ i_9_)  &  (~ i_16_) ) ;
 assign wire805 = ( wire45  &  n_n880 ) | ( wire316  &  wire421 ) ;
 assign wire808 = ( i_3_ ) | ( i_4_ ) | ( i_1_ ) ;
 assign wire807 = ( i_40_  &  (~ i_38_) ) | ( i_39_  &  (~ i_38_) ) ;
 assign wire7258 = ( i_35_  &  i_38_  &  i_37_ ) ;
 assign wire811 = ( i_34_  &  wire46  &  n_n1073 ) | ( (~ i_34_)  &  wire46  &  wire7258 ) ;
 assign wire7256 = ( (~ i_34_)  &  i_35_  &  i_38_  &  i_37_ ) ;
 assign wire7257 = ( (~ i_9_)  &  i_39_  &  i_38_ ) ;
 assign wire809 = ( (~ i_38_)  &  wire464 ) | ( i_2_  &  (~ i_38_)  &  i_37_ ) ;
 assign wire63 = ( i_9_  &  (~ i_5_)  &  (~ i_12_) ) | ( i_9_  &  (~ i_5_)  &  (~ i_11_) ) ;
 assign wire814 = ( wire63 ) | ( i_9_  &  (~ i_5_)  &  (~ i_15_) ) ;
 assign wire818 = ( (~ i_9_)  &  (~ i_17_) ) | ( (~ i_9_)  &  (~ i_16_) ) | ( (~ i_17_)  &  (~ i_16_) ) ;
 assign wire7074 = ( i_5_  &  (~ i_36_)  &  (~ i_35_) ) ;
 assign wire817 = ( n_n977  &  n_n971 ) | ( wire818  &  wire7074 ) ;
 assign wire7452 = ( (~ i_40_)  &  i_39_  &  (~ i_23_)  &  i_38_ ) ;
 assign wire822 = ( (~ i_40_)  &  i_39_  &  i_38_ ) | ( (~ i_40_)  &  (~ i_39_)  &  (~ i_38_) ) ;
 assign wire825 = ( (~ i_40_)  &  i_39_  &  n_n1009 ) | ( (~ i_40_)  &  (~ i_39_)  &  n_n1052 ) ;
 assign wire1570 = ( i_17_  &  i_16_  &  n_n1072  &  n_n1073 ) ;
 assign wire1571 = ( i_40_  &  i_39_  &  _9823 ) | ( i_39_  &  (~ i_38_)  &  _9823 ) ;
 assign wire7058 = ( n_n1011  &  n_n1012 ) | ( n_n1009  &  n_n1008 ) ;
 assign wire55 = ( (~ i_9_)  &  (~ i_17_) ) | ( (~ i_17_)  &  (~ i_16_) ) ;
 assign wire304 = ( (~ i_40_)  &  (~ i_39_)  &  (~ i_38_)  &  (~ i_37_) ) ;
 assign wire1795 = ( i_12_  &  (~ i_21_)  &  i_15_  &  i_19_ ) ;
 assign wire1797 = ( i_11_  &  i_15_  &  i_19_ ) ;
 assign wire1798 = ( i_12_  &  i_18_  &  i_15_ ) ;
 assign wire70 = ( wire1795 ) | ( _1080 ) | ( _1081 ) ;
 assign wire7818 = ( (~ i_12_)  &  i_11_  &  i_15_ ) ;
 assign wire7819 = ( (~ i_14_)  &  i_12_  &  i_15_ ) ;
 assign wire104 = ( n_n642  &  wire7818 ) | ( n_n643  &  wire7818 ) | ( n_n643  &  wire7819 ) ;
 assign wire121 = ( (~ i_40_)  &  (~ i_38_)  &  (~ i_37_) ) | ( (~ i_39_)  &  (~ i_38_)  &  (~ i_37_) ) ;
 assign wire830 = ( (~ i_40_)  &  i_39_  &  n_n1009 ) | ( (~ i_40_)  &  (~ i_39_)  &  n_n1052 ) ;
 assign wire829 = ( i_40_  &  (~ i_39_)  &  n_n985 ) | ( (~ i_40_)  &  (~ i_39_)  &  n_n1052 ) ;
 assign wire831 = ( (~ wire37)  &  n_n1048  &  wire82 ) | ( (~ wire37)  &  n_n1048  &  wire87 ) ;
 assign wire837 = ( i_39_  &  i_38_ ) | ( i_40_  &  (~ i_38_) ) ;
 assign wire375 = ( (~ i_30_)  &  (~ i_29_) ) ;
 assign wire482 = ( i_24_  &  i_22_  &  n_n1074  &  n_n968 ) ;
 assign wire7510 = ( i_39_  &  i_23_  &  i_38_ ) ;
 assign wire481 = ( i_16_  &  wire82  &  wire320 ) ;
 assign wire841 = ( (~ i_7_)  &  (~ i_5_)  &  (~ i_12_)  &  i_11_ ) | ( (~ i_7_)  &  (~ i_5_)  &  i_12_  &  (~ i_11_) ) ;
 assign wire840 = ( (~ i_14_)  &  wire469 ) | ( i_16_  &  wire841 ) ;
 assign wire7817 = ( i_17_  &  i_15_  &  (~ i_32_)  &  i_33_ ) ;
 assign wire546 = ( n_n1061  &  wire50 ) | ( wire80  &  n_n582 ) ;
 assign wire548 = ( (~ i_40_)  &  (~ i_38_) ) | ( (~ i_39_)  &  (~ i_38_) ) ;
 assign wire558 = ( n_n933  &  n_n1066 ) | ( n_n1066  &  n_n927 ) ;
 assign wire589 = ( (~ i_40_)  &  i_39_  &  n_n1009 ) | ( i_40_  &  (~ i_39_)  &  n_n985 ) ;
 assign wire609 = ( i_12_  &  i_18_  &  i_15_ ) | ( i_11_  &  i_18_  &  i_15_ ) ;
 assign wire636 = ( (~ i_34_)  &  n_n865  &  wire46 ) | ( i_34_  &  wire46  &  n_n1073 ) ;
 assign wire642 = ( wire330  &  n_n998 ) | ( n_n979  &  wire60 ) ;
 assign wire652 = ( n_n998  &  n_n866 ) | ( n_n977  &  n_n888 ) ;
 assign wire650 = ( (~ i_5_)  &  i_12_  &  i_15_ ) | ( (~ i_5_)  &  i_11_  &  i_15_ ) ;
 assign wire687 = ( i_17_ ) | ( i_16_ ) ;
 assign wire686 = ( i_12_  &  wire407 ) | ( wire484  &  wire687 ) ;
 assign wire716 = ( (~ i_39_)  &  (~ i_38_)  &  i_37_ ) | ( i_39_  &  i_38_  &  (~ i_37_) ) ;
 assign wire715 = ( n_n795  &  n_n976 ) | ( n_n983  &  wire716 ) ;
 assign wire721 = ( i_37_  &  n_n1011  &  n_n964 ) | ( (~ i_37_)  &  n_n1072  &  n_n964 ) ;
 assign wire7007 = ( (~ i_12_)  &  i_11_  &  i_15_ ) ;
 assign wire7008 = ( i_17_  &  i_15_  &  (~ i_32_)  &  (~ i_31_) ) ;
 assign wire729 = ( n_n927  &  wire7007 ) | ( wire39  &  wire7008 ) ;
 assign wire1048 = ( (~ i_40_)  &  (~ i_39_)  &  wire50  &  n_n1052 ) ;
 assign wire731 = ( (~ i_7_)  &  (~ i_5_)  &  i_12_ ) | ( (~ i_7_)  &  (~ i_5_)  &  i_11_ ) ;
 assign wire743 = ( i_40_  &  i_39_ ) | ( i_40_  &  (~ i_38_) ) | ( i_39_  &  (~ i_38_) ) ;
 assign wire845 = ( (~ i_31_)  &  wire45  &  wire43 ) ;
 assign wire1300 = ( (~ i_30_)  &  (~ i_7_)  &  (~ i_5_)  &  i_29_ ) | ( i_30_  &  (~ i_7_)  &  (~ i_5_)  &  (~ i_29_) ) ;
 assign wire765 = ( wire43 ) | ( wire1300 ) ;
 assign wire1400 = ( i_9_  &  i_12_  &  i_15_ ) ;
 assign wire785 = ( i_40_  &  i_39_  &  (~ i_37_) ) | ( i_39_  &  (~ i_38_)  &  (~ i_37_) ) ;
 assign wire793 = ( i_9_  &  n_n833 ) | ( i_13_  &  wire371 ) ;
 assign wire792 = ( (~ i_39_)  &  (~ i_36_)  &  (~ i_38_)  &  i_37_ ) | ( i_39_  &  (~ i_36_)  &  (~ i_38_)  &  (~ i_37_) ) ;
 assign wire1563 = ( i_39_  &  i_36_  &  i_38_  &  (~ i_37_) ) ;
 assign wire797 = ( wire1563 ) | ( i_40_  &  (~ i_39_)  &  n_n1065 ) ;
 assign wire801 = ( i_37_  &  n_n1011  &  n_n964 ) | ( (~ i_37_)  &  wire66  &  n_n964 ) ;
 assign wire7182 = ( i_9_  &  (~ i_5_)  &  (~ i_12_) ) ;
 assign wire813 = ( n_n933  &  wire63 ) | ( n_n927  &  wire7182 ) ;
 assign wire820 = ( (~ i_39_)  &  (~ i_38_)  &  i_37_ ) | ( i_39_  &  i_38_  &  (~ i_37_) ) ;
 assign wire824 = ( n_n969  &  n_n968 ) | ( n_n978  &  wire6907 ) ;
 assign wire7815 = ( i_9_  &  (~ i_7_)  &  (~ i_5_)  &  (~ i_21_) ) ;
 assign wire7803 = ( (~ i_34_)  &  i_36_  &  (~ i_37_) ) ;
 assign wire142 = ( n_n883  &  n_n861  &  wire7803 ) ;
 assign wire7805 = ( (~ i_40_)  &  (~ i_39_)  &  i_37_ ) ;
 assign wire143 = ( n_n979  &  n_n861  &  wire7805 ) ;
 assign wire7806 = ( (~ i_9_)  &  (~ i_7_)  &  (~ i_5_)  &  (~ i_17_) ) ;
 assign wire144 = ( i_31_  &  (~ i_36_)  &  wire45  &  wire7806 ) ;
 assign wire6728 = ( (~ i_32_)  &  i_31_  &  i_33_ ) ;
 assign wire151 = ( n_n1047  &  wire420  &  wire6728 ) ;
 assign wire162 = ( (~ i_36_)  &  (~ i_35_)  &  i_38_  &  i_37_ ) ;
 assign wire163 = ( i_39_  &  (~ i_36_)  &  (~ i_35_)  &  (~ i_38_) ) ;
 assign wire164 = ( (~ i_36_)  &  (~ i_35_)  &  (~ i_38_)  &  (~ i_37_) ) ;
 assign wire165 = ( wire50  &  n_n693  &  _11256 ) ;
 assign wire7796 = ( (~ i_7_)  &  (~ i_5_)  &  (~ i_12_) ) ;
 assign wire167 = ( n_n1047  &  wire6728  &  wire7796 ) ;
 assign wire169 = ( wire88  &  n_n982  &  n_n998 ) ;
 assign wire170 = ( wire88  &  n_n997  &  n_n991 ) ;
 assign wire171 = ( n_n469  &  n_n1002  &  n_n861 ) ;
 assign wire188 = ( n_n979  &  n_n330  &  wire602  &  n_n700 ) ;
 assign wire190 = ( wire45  &  n_n462  &  n_n801  &  wire375 ) ;
 assign wire191 = ( n_n977  &  n_n861  &  n_n710  &  n_n715 ) ;
 assign wire192 = ( n_n998  &  n_n861  &  n_n799  &  n_n710 ) ;
 assign wire193 = ( n_n883  &  n_n1002  &  n_n861  &  n_n710 ) ;
 assign wire7777 = ( i_39_  &  (~ i_36_)  &  (~ i_38_)  &  i_37_ ) ;
 assign wire198 = ( i_13_  &  wire80  &  wire315  &  wire7777 ) ;
 assign wire199 = ( n_n975  &  wire46  &  wire94  &  wire315 ) ;
 assign wire7276 = ( (~ i_7_)  &  (~ i_5_)  &  (~ i_13_) ) ;
 assign wire201 = ( n_n1047  &  wire325  &  n_n700  &  wire7276 ) ;
 assign wire206 = ( wire50  &  wire315  &  _11184 ) ;
 assign wire207 = ( n_n998  &  n_n975  &  n_n861  &  n_n710 ) ;
 assign wire205 = ( i_13_  &  wire50  &  wire54  &  wire315 ) ;
 assign wire7767 = ( i_12_  &  (~ i_11_)  &  i_36_  &  (~ i_35_) ) ;
 assign wire208 = ( n_n973  &  wire79  &  wire7767 ) ;
 assign wire209 = ( n_n998  &  n_n330  &  n_n795  &  n_n700 ) ;
 assign wire210 = ( wire50  &  n_n693  &  _11170 ) ;
 assign wire7771 = ( (~ i_9_)  &  (~ i_7_)  &  (~ i_5_)  &  (~ i_16_) ) ;
 assign wire211 = ( i_31_  &  (~ i_36_)  &  wire45  &  wire7771 ) ;
 assign wire213 = ( (~ i_40_)  &  (~ i_7_)  &  wire50  &  wire6920 ) ;
 assign wire217 = ( wire45  &  n_n462  &  _11092 ) ;
 assign wire218 = ( _101 ) | ( n_n874  &  n_n884  &  wire589 ) ;
 assign wire7760 = ( (~ i_5_)  &  (~ i_13_)  &  (~ i_12_) ) ;
 assign wire229 = ( (~ i_9_)  &  (~ i_5_)  &  wire45  &  n_n997 ) ;
 assign wire231 = ( n_n1002  &  n_n975  &  _11153 ) ;
 assign wire232 = ( n_n1074  &  n_n864  &  n_n883 ) ;
 assign wire234 = ( n_n1055  &  n_n998  &  _11155 ) ;
 assign wire235 = ( n_n966  &  n_n1012  &  n_n978 ) ;
 assign wire7743 = ( i_40_  &  i_36_  &  i_37_ ) ;
 assign wire248 = ( n_n1023  &  n_n458  &  wire403 ) ;
 assign wire7745 = ( i_12_  &  (~ i_11_)  &  i_36_ ) ;
 assign wire250 = ( (~ i_40_)  &  i_39_  &  n_n979  &  wire7227 ) ;
 assign wire252 = ( n_n1055  &  n_n998  &  _11089 ) ;
 assign wire260 = ( n_n1074  &  wire6731  &  wire665 ) ;
 assign wire261 = ( n_n966  &  n_n1073  &  wire666 ) ;
 assign wire6739 = ( (~ i_5_)  &  i_31_  &  (~ i_36_)  &  (~ i_35_) ) ;
 assign wire276 = ( wire45  &  (~ wire37)  &  n_n926  &  n_n947 ) ;
 assign wire279 = ( wire445  &  n_n492  &  wire352  &  wire421 ) ;
 assign wire7717 = ( i_14_  &  i_15_ ) | ( (~ i_17_)  &  i_15_ ) ;
 assign wire7707 = ( i_40_  &  (~ i_16_)  &  i_15_  &  (~ i_38_) ) ;
 assign wire298 = ( n_n1023  &  n_n843  &  n_n1065  &  n_n1057 ) ;
 assign wire299 = ( (~ i_40_)  &  (~ i_36_)  &  (~ i_37_) ) ;
 assign wire7698 = ( i_39_  &  (~ i_16_)  &  i_15_ ) ;
 assign wire309 = ( (~ i_36_)  &  wire45  &  n_n488  &  wire7698 ) ;
 assign wire310 = ( n_n1074  &  n_n1021  &  n_n862  &  wire635 ) ;
 assign wire311 = ( _105 ) | ( n_n1008  &  n_n710  &  wire636 ) ;
 assign wire7689 = ( (~ i_5_)  &  i_15_  &  (~ i_32_)  &  i_33_ ) ;
 assign wire312 = ( n_n1055  &  n_n1047  &  wire39  &  wire7689 ) ;
 assign wire7694 = ( (~ i_23_)  &  (~ i_32_)  &  i_33_ ) ;
 assign wire7686 = ( (~ i_5_)  &  (~ i_12_)  &  i_15_ ) ;
 assign wire455 = ( n_n1073  &  wire7689  &  _11112 ) ;
 assign wire7670 = ( i_40_  &  (~ i_39_)  &  i_24_  &  (~ i_37_) ) ;
 assign wire519 = ( wire50  &  wire82  &  wire7670 ) | ( wire50  &  wire87  &  wire7670 ) ;
 assign wire533 = ( n_n1066  &  n_n462  &  wire7122  &  wire494 ) ;
 assign wire843 = ( n_n1002  &  n_n861  &  n_n710  &  wire100 ) ;
 assign wire538 = ( n_n883  &  n_n1002  &  n_n861  &  n_n710 ) ;
 assign wire850 = ( i_13_  &  wire315  &  wire76  &  wire401 ) ;
 assign wire859 = ( n_n1048  &  n_n1047  &  wire420  &  wire697 ) ;
 assign wire860 = ( wire330  &  n_n998  &  n_n700  &  wire7276 ) ;
 assign wire864 = ( n_n998  &  n_n861  &  wire441 ) ;
 assign wire865 = ( (~ i_38_)  &  (~ i_37_)  &  n_n1002  &  n_n861 ) ;
 assign wire872 = ( i_13_  &  wire50  &  n_n528  &  wire315 ) ;
 assign wire873 = ( n_n977  &  n_n1002  &  n_n861  &  n_n710 ) ;
 assign wire888 = ( (~ i_12_)  &  (~ i_31_)  &  wire45 ) | ( (~ i_11_)  &  (~ i_31_)  &  wire45 ) ;
 assign wire7640 = ( (~ i_40_)  &  i_39_  &  n_n1009  &  n_n860 ) ;
 assign wire7627 = ( (~ i_40_)  &  i_39_  &  i_0_ ) ;
 assign wire890 = ( wire50  &  wire7627  &  _10886 ) ;
 assign wire7630 = ( (~ i_40_)  &  i_35_  &  (~ i_38_)  &  i_37_ ) ;
 assign wire7631 = ( i_4_  &  i_0_ ) ;
 assign wire892 = ( _245 ) | ( wire79  &  wire402  &  wire7631 ) ;
 assign wire893 = ( n_n998  &  n_n861  &  wire495 ) ;
 assign wire894 = ( (~ i_7_)  &  i_2_  &  wire80  &  n_n926 ) ;
 assign wire904 = ( n_n991  &  wire740  &  _10867 ) ;
 assign wire7620 = ( (~ i_7_)  &  i_12_  &  (~ i_32_) ) ;
 assign wire905 = ( wire325  &  n_n1056  &  wire7620 ) ;
 assign wire906 = ( wire88  &  n_n982  &  n_n998 ) ;
 assign wire911 = ( n_n975  &  wire94  &  n_n700  &  wire7276 ) ;
 assign wire912 = ( _294 ) | ( _295 ) ;
 assign wire922 = ( n_n1048  &  n_n1047  &  n_n527 ) ;
 assign wire7610 = ( n_n1048  &  n_n1047  &  wire420 ) | ( n_n1048  &  n_n1047  &  wire6884 ) ;
 assign wire913 = ( n_n469  &  wire922 ) | ( n_n469  &  wire7610 ) ;
 assign wire930 = ( (~ i_40_)  &  i_35_  &  (~ i_38_)  &  i_37_ ) ;
 assign wire932 = ( n_n1048  &  wire934  &  wire7602 ) | ( n_n1048  &  wire7601  &  wire7602 ) ;
 assign wire928 = ( n_n971  &  wire79  &  _10804 ) ;
 assign wire929 = ( (~ i_7_)  &  i_2_  &  wire80  &  n_n833 ) ;
 assign wire934 = ( i_30_  &  (~ i_7_)  &  (~ i_5_) ) ;
 assign wire7601 = ( (~ i_7_)  &  (~ i_5_)  &  i_28_ ) | ( (~ i_7_)  &  (~ i_5_)  &  i_29_ ) ;
 assign wire7602 = ( (~ i_34_)  &  (~ i_38_)  &  i_37_ ) ;
 assign wire7593 = ( (~ i_7_)  &  (~ i_5_)  &  (~ i_29_) ) ;
 assign wire937 = ( n_n1066  &  n_n462  &  wire7122  &  wire7593 ) ;
 assign wire939 = ( (~ i_39_)  &  (~ i_36_)  &  (~ i_38_)  &  wire744 ) ;
 assign wire940 = ( n_n998  &  n_n861  &  n_n710  &  wire124 ) ;
 assign wire948 = ( n_n1048  &  n_n1072  &  n_n1073 ) ;
 assign wire7586 = ( (~ i_14_)  &  i_12_  &  i_15_ ) ;
 assign wire942 = ( n_n853  &  wire84  &  wire7586 ) | ( n_n853  &  wire948  &  wire7586 ) ;
 assign wire967 = ( (~ i_40_)  &  (~ i_39_)  &  (~ i_36_)  &  (~ i_38_) ) ;
 assign wire7572 = ( wire48  &  wire50  &  n_n853 ) | ( wire48  &  wire50  &  n_n850 ) ;
 assign wire962 = ( n_n833  &  n_n764 ) | ( n_n764  &  wire967 ) | ( n_n833  &  wire7572 ) | ( wire967  &  wire7572 ) ;
 assign wire964 = ( (~ i_22_)  &  wire50  &  n_n926  &  wire82 ) ;
 assign wire973 = ( n_n1002  &  n_n861  &  wire441  &  n_n710 ) ;
 assign wire985 = ( n_n861  &  n_n799  &  wire624 ) ;
 assign wire987 = ( (~ i_38_)  &  i_37_  &  n_n979  &  wire88 ) ;
 assign wire988 = ( n_n990  &  n_n1002  &  n_n861 ) ;
 assign wire7127 = ( i_15_  &  wire42 ) ;
 assign wire999 = ( n_n1072  &  wire380  &  wire482 ) | ( n_n1072  &  wire482  &  wire7127 ) ;
 assign wire1000 = ( n_n978  &  n_n937  &  wire6907 ) ;
 assign wire1008 = ( n_n1074  &  n_n864  &  n_n883 ) ;
 assign wire1010 = ( n_n966  &  n_n973  &  n_n1073 ) ;
 assign wire7521 = ( n_n411  &  wire1834 ) | ( i_18_  &  n_n411  &  wire42 ) ;
 assign wire1019 = ( wire512  &  wire7521 ) ;
 assign wire7522 = ( n_n1074  &  wire6731  &  wire491  &  n_n978 ) ;
 assign wire1020 = ( wire7522  &  _10718 ) | ( wire36  &  wire7522  &  _9284 ) ;
 assign wire1021 = ( n_n1048  &  n_n1047  &  wire579  &  _9306 ) ;
 assign wire1029 = ( i_9_  &  (~ i_5_)  &  (~ i_11_)  &  _10712 ) ;
 assign wire1022 = ( wire84  &  wire1029 ) | ( n_n955  &  wire84  &  _9041 ) ;
 assign wire1038 = ( n_n952  &  wire7514 ) | ( n_n427  &  wire7514 ) | ( wire1040  &  wire7514 ) ;
 assign wire1040 = ( (~ i_40_)  &  (~ i_39_)  &  n_n1052  &  n_n1023 ) ;
 assign wire7514 = ( wire82  &  n_n428 ) | ( wire87  &  n_n428 ) ;
 assign wire1046 = ( n_n968  &  wire7510  &  _10693  &  _10696 ) ;
 assign wire7511 = ( i_25_  &  i_21_  &  i_22_  &  i_15_ ) ;
 assign wire7500 = ( (~ i_7_)  &  (~ i_38_) ) ;
 assign wire1049 = ( n_n1047  &  n_n980  &  wire574  &  wire7500 ) ;
 assign wire1050 = ( _409 ) | ( _410 ) ;
 assign wire1051 = ( n_n1074  &  n_n865  &  _10668 ) ;
 assign wire1060 = ( n_n469  &  n_n983  &  n_n668 ) ;
 assign wire1063 = ( n_n1052  &  n_n874  &  _10607 ) ;
 assign wire1075 = ( n_n685  &  n_n1074  &  n_n971  &  n_n1072 ) ;
 assign wire1084 = ( n_n1047  &  n_n1001  &  wire344  &  wire38 ) ;
 assign wire1085 = ( wire79  &  n_n1073  &  _10636 ) ;
 assign wire1083 = ( (~ i_12_)  &  wire1084 ) | ( (~ i_12_)  &  wire1085 ) ;
 assign wire7479 = ( (~ i_7_)  &  (~ i_34_)  &  (~ i_36_) ) ;
 assign wire1088 = ( n_n980  &  n_n1001  &  wire674  &  wire7479 ) ;
 assign wire7482 = ( (~ i_7_)  &  (~ i_14_) ) | ( (~ i_7_)  &  (~ i_12_) ) | ( (~ i_7_)  &  (~ i_11_) ) ;
 assign wire1089 = ( n_n1055  &  n_n1047  &  wire351  &  wire7482 ) ;
 assign wire1090 = ( n_n1074  &  n_n969  &  n_n968  &  n_n629 ) ;
 assign wire1091 = ( n_n685  &  n_n1074  &  n_n1064  &  n_n1065 ) ;
 assign wire1092 = ( n_n1074  &  n_n967  &  n_n629  &  n_n1073 ) ;
 assign wire1093 = ( wire717  &  wire6728  &  _10588 ) ;
 assign wire1112 = ( _406 ) | ( _407 ) | ( _408 ) ;
 assign wire1114 = ( (~ i_36_)  &  wire1119 ) | ( (~ i_36_)  &  wire1120 ) ;
 assign wire7466 = ( i_40_  &  i_39_  &  n_n1009 ) | ( i_40_  &  (~ i_39_)  &  n_n985 ) ;
 assign wire7467 = ( n_n1064  &  n_n993 ) | ( n_n1073  &  n_n1015 ) ;
 assign wire1113 = ( wire390  &  wire1114 ) | ( wire390  &  wire7466 ) | ( wire390  &  wire7467 ) ;
 assign wire1119 = ( i_40_  &  (~ i_39_)  &  i_13_  &  (~ i_38_) ) ;
 assign wire1120 = ( i_9_  &  i_39_  &  i_38_  &  (~ i_37_) ) ;
 assign wire1122 = ( n_n969  &  n_n968  &  n_n819 ) ;
 assign wire7435 = ( (~ i_4_)  &  i_0_  &  i_36_ ) ;
 assign wire1155 = ( wire50  &  wire403  &  wire7435 ) ;
 assign wire1156 = ( n_n1055  &  n_n998  &  _10535 ) ;
 assign wire1158 = ( n_n1074  &  n_n865  &  n_n799 ) ;
 assign wire7347 = ( (~ i_23_)  &  (~ i_32_)  &  i_33_ ) ;
 assign wire1164 = ( n_n979  &  n_n469  &  n_n949  &  wire7347 ) ;
 assign wire1165 = ( n_n979  &  n_n949  &  wire60  &  wire7406 ) ;
 assign wire7415 = ( i_39_  &  (~ i_36_)  &  (~ i_35_)  &  i_38_ ) ;
 assign wire7121 = ( (~ i_40_)  &  (~ i_5_)  &  i_39_ ) ;
 assign wire1182 = ( n_n979  &  n_n949  &  wire60  &  n_n791 ) ;
 assign wire1186 = ( n_n979  &  n_n949  &  wire7405  &  wire615 ) ;
 assign wire1189 = ( n_n979  &  n_n975  &  n_n947  &  wire7399 ) ;
 assign wire1199 = ( n_n1023  &  n_n843  &  n_n1065  &  n_n1057 ) ;
 assign wire1200 = ( n_n1066  &  n_n1064  &  n_n1065  &  n_n458 ) ;
 assign wire7388 = ( (~ i_40_)  &  (~ i_1_)  &  i_2_  &  i_0_ ) ;
 assign wire1208 = ( n_n979  &  n_n947  &  wire60  &  wire7390 ) ;
 assign wire1219 = ( (~ i_4_)  &  i_0_  &  wire79 ) | ( (~ i_1_)  &  i_0_  &  wire79 ) ;
 assign wire7372 = ( n_n1074  &  wire6828 ) | ( n_n1074  &  wire6897 ) ;
 assign wire1213 = ( n_n865  &  wire373  &  wire1219 ) | ( n_n865  &  wire373  &  wire7372 ) ;
 assign wire7360 = ( (~ i_39_)  &  (~ i_32_)  &  i_34_  &  i_33_ ) ;
 assign wire1222 = ( n_n842  &  n_n843  &  n_n993  &  wire7360 ) ;
 assign wire1230 = ( (~ i_24_)  &  wire50  &  wire82  &  wire371 ) ;
 assign wire1238 = ( (~ i_39_)  &  i_38_  &  n_n998  &  n_n861 ) ;
 assign wire1246 = ( n_n979  &  n_n795  &  n_n861 ) ;
 assign wire1247 = ( n_n977  &  n_n861  &  n_n991 ) ;
 assign wire1251 = ( (~ i_40_)  &  (~ i_10_)  &  i_38_ ) | ( (~ i_40_)  &  (~ i_27_)  &  i_38_ ) ;
 assign wire1252 = ( i_40_  &  (~ i_11_)  &  (~ i_38_) ) ;
 assign wire7332 = ( (~ i_40_)  &  i_39_  &  i_37_ ) ;
 assign wire1253 = ( n_n998  &  n_n861  &  wire7332 ) ;
 assign wire7334 = ( n_n709  &  n_n1002 ) | ( n_n991  &  wire7333 ) ;
 assign wire1254 = ( n_n861  &  wire7334 ) | ( n_n969  &  n_n971  &  n_n861 ) ;
 assign wire1255 = ( i_38_  &  i_37_  &  n_n861  &  wire94 ) ;
 assign wire1256 = ( (~ i_38_)  &  i_37_  &  n_n979  &  wire88 ) ;
 assign wire1257 = ( n_n1005  &  n_n979  &  n_n861 ) ;
 assign wire1262 = ( n_n883  &  n_n861  &  n_n888 ) ;
 assign wire7323 = ( wire78  &  wire320  &  n_n860 ) | ( wire86  &  wire320  &  n_n860 ) ;
 assign wire7324 = ( i_40_  &  i_39_  &  (~ i_36_)  &  (~ i_38_) ) ;
 assign wire1264 = ( n_n535  &  wire7324 ) | ( wire481  &  wire7324 ) | ( wire7323  &  wire7324 ) ;
 assign wire7325 = ( (~ i_40_)  &  (~ i_39_)  &  (~ i_36_)  &  i_38_ ) ;
 assign wire1265 = ( wire481  &  wire7325 ) | ( wire7323  &  wire7325 ) ;
 assign wire7314 = ( (~ i_40_)  &  (~ i_31_)  &  (~ i_34_)  &  i_33_ ) ;
 assign wire1271 = ( n_n862  &  n_n860  &  (~ wire166)  &  wire7314 ) ;
 assign wire7308 = ( i_9_  &  (~ i_7_)  &  (~ wire73)  &  wire7306 ) ;
 assign wire1286 = ( n_n998  &  n_n861  &  n_n799  &  n_n710 ) ;
 assign wire1294 = ( (~ i_7_)  &  wire471  &  wire80  &  wire763 ) ;
 assign wire1299 = ( i_16_  &  wire87  &  wire320  &  n_n688 ) ;
 assign wire7291 = ( (~ i_31_)  &  i_33_  &  n_n1047  &  n_n795 ) ;
 assign wire1295 = ( (~ i_40_)  &  wire1299 ) | ( (~ i_40_)  &  wire765  &  wire7291 ) ;
 assign wire7275 = ( (~ i_40_)  &  (~ i_36_)  &  i_38_ ) ;
 assign wire1305 = ( (~ i_7_)  &  wire471  &  wire80  &  wire7275 ) ;
 assign wire1306 = ( n_n888  &  n_n1064  &  n_n700  &  wire7276 ) ;
 assign wire7278 = ( (~ i_39_)  &  (~ i_37_) ) ;
 assign wire1307 = ( n_n998  &  n_n861  &  n_n710  &  wire7278 ) ;
 assign wire1309 = ( n_n710  &  n_n715  &  _10277 ) ;
 assign wire7279 = ( i_40_  &  (~ i_30_)  &  (~ i_39_)  &  i_38_ ) ;
 assign wire7281 = ( i_9_  &  (~ i_7_)  &  (~ i_5_)  &  (~ i_34_) ) ;
 assign wire1316 = ( n_n862  &  _10212 ) | ( n_n862  &  _10213 ) ;
 assign wire1326 = ( i_40_  &  (~ i_36_)  &  i_38_  &  (~ i_37_) ) ;
 assign wire1317 = ( n_n874  &  n_n462 ) | ( n_n874  &  wire1326 ) ;
 assign wire7253 = ( (~ i_9_)  &  i_39_  &  (~ i_16_) ) ;
 assign wire1328 = ( (~ i_36_)  &  wire45  &  wire7253 ) ;
 assign wire1329 = ( (~ i_12_)  &  (~ i_11_)  &  wire45  &  n_n918 ) ;
 assign wire1330 = ( (~ i_38_)  &  (~ i_37_)  &  n_n1006  &  n_n976 ) ;
 assign wire7246 = ( i_0_  &  (~ i_32_)  &  i_33_ ) ;
 assign wire1340 = ( (~ i_40_)  &  (~ i_38_)  &  n_n715  &  wire7246 ) ;
 assign wire1341 = ( n_n998  &  wire808  &  _10207 ) ;
 assign wire1342 = ( n_n966  &  n_n1012  &  wire807 ) ;
 assign wire1343 = ( i_35_  &  (~ i_37_)  &  n_n1074  &  n_n977 ) ;
 assign wire1344 = ( (~ i_40_)  &  i_39_  &  n_n1074  &  n_n698 ) ;
 assign wire7239 = ( i_39_  &  (~ i_32_)  &  i_33_  &  i_38_ ) ;
 assign wire1346 = ( wire7239  &  _10186 ) | ( wire7239  &  _10187 ) ;
 assign wire1347 = ( (~ i_39_)  &  i_38_  &  n_n1074  &  n_n971 ) ;
 assign wire1348 = ( i_39_  &  (~ i_38_)  &  n_n1047  &  n_n700 ) ;
 assign wire7231 = ( (~ i_34_)  &  i_33_  &  i_38_  &  i_37_ ) ;
 assign wire1353 = ( i_5_  &  (~ i_0_)  &  (~ i_32_)  &  wire7231 ) ;
 assign wire1354 = ( (~ i_40_)  &  (~ i_39_)  &  n_n874  &  n_n693 ) ;
 assign wire1362 = ( (~ i_34_)  &  i_36_  &  (~ i_35_)  &  _10141 ) ;
 assign wire7234 = ( n_n1073  &  n_n700 ) | ( n_n1074  &  wire7233 ) ;
 assign wire1366 = ( wire6731  &  _10179 ) | ( wire6731  &  _10180 ) ;
 assign wire7214 = ( (~ i_40_)  &  (~ i_39_)  &  i_38_  &  i_37_ ) | ( (~ i_40_)  &  (~ i_39_)  &  (~ i_38_)  &  (~ i_37_) ) ;
 assign wire1381 = ( (~ i_9_)  &  i_5_  &  (~ i_17_) ) | ( (~ i_9_)  &  i_5_  &  (~ i_16_) ) ;
 assign wire1372 = ( i_32_  &  n_n1047  &  wire7191 ) | ( n_n1047  &  wire7191  &  wire1381 ) ;
 assign wire1374 = ( n_n685  &  (~ n_n1014)  &  n_n1052  &  n_n874 ) ;
 assign wire1375 = ( n_n1074  &  n_n865  &  _10131 ) ;
 assign wire7205 = ( (~ i_40_)  &  i_9_  &  (~ i_7_) ) ;
 assign wire1383 = ( wire320  &  wire383  &  (~ wire166)  &  wire7205 ) ;
 assign wire1386 = ( n_n685  &  n_n1074  &  n_n971  &  n_n1072 ) ;
 assign wire1388 = ( i_11_  &  i_16_  &  i_15_ ) ;
 assign wire1389 = ( i_9_  &  i_12_  &  i_15_ ) ;
 assign wire1390 = ( n_n1074  &  wire779  &  _10082 ) ;
 assign wire7197 = ( (~ i_7_)  &  i_5_  &  (~ i_36_) ) ;
 assign wire1412 = ( (~ i_39_)  &  i_38_  &  n_n966  &  n_n1073 ) ;
 assign wire7181 = ( (~ i_40_)  &  (~ i_39_)  &  (~ i_38_)  &  i_37_ ) ;
 assign wire1415 = ( wire471  &  n_n998  &  wire46  &  wire7181 ) ;
 assign wire1416 = ( _772 ) | ( n_n1066  &  n_n923  &  wire813 ) ;
 assign wire1417 = ( n_n979  &  n_n907  &  wire6716  &  wire342 ) ;
 assign wire1428 = ( n_n1048  &  n_n1047  &  n_n880  &  n_n907 ) ;
 assign wire1429 = ( _785 ) | ( wire378  &  wire76  &  wire801 ) ;
 assign wire1430 = ( _781 ) | ( _782 ) | ( _783 ) ;
 assign wire7164 = ( i_40_  &  i_6_  &  (~ i_38_)  &  i_37_ ) ;
 assign wire1442 = ( (~ i_32_)  &  i_33_  &  n_n1002  &  wire7164 ) ;
 assign wire1444 = ( n_n966  &  n_n1014  &  n_n993  &  n_n884 ) ;
 assign wire7165 = ( i_39_  &  i_12_  &  (~ i_38_)  &  (~ i_37_) ) ;
 assign wire7157 = ( (~ i_34_)  &  n_n968  &  wire46 ) | ( i_34_  &  wire46  &  n_n1073 ) ;
 assign wire1452 = ( n_n973  &  wire7157 ) | ( n_n1074  &  n_n973  &  n_n865 ) ;
 assign wire1453 = ( (~ i_40_)  &  i_39_  &  n_n1074  &  n_n1061 ) ;
 assign wire1454 = ( (~ i_39_)  &  (~ i_38_)  &  n_n1074  &  n_n864 ) ;
 assign wire7063 = ( i_1_  &  (~ i_2_)  &  i_0_ ) ;
 assign wire7148 = ( (~ i_40_)  &  (~ i_39_)  &  i_36_  &  (~ i_38_) ) ;
 assign wire1459 = ( n_n1023  &  n_n1057  &  wire7063  &  wire7148 ) ;
 assign wire1466 = ( _765 ) | ( _766 ) ;
 assign wire1472 = ( n_n1048  &  n_n967  &  n_n1073 ) ;
 assign wire7142 = ( n_n1055  &  n_n1048  &  n_n1047 ) | ( n_n1048  &  n_n1047  &  wire785 ) ;
 assign wire1467 = ( n_n907  &  wire1472 ) | ( n_n907  &  wire7142 ) ;
 assign wire1468 = ( n_n979  &  n_n1001  &  n_n907  &  wire6716 ) ;
 assign wire1496 = ( n_n1074  &  n_n971  &  n_n880  &  n_n629 ) ;
 assign wire1499 = ( wire88  &  n_n998  &  n_n997 ) ;
 assign wire1501 = ( n_n975  &  n_n861  &  n_n991 ) ;
 assign wire7103 = ( n_n1002  &  wire100 ) | ( n_n883  &  wire7102 ) ;
 assign wire7104 = ( n_n977  &  n_n715 ) | ( n_n998  &  wire121 ) ;
 assign wire7105 = ( (~ i_7_)  &  (~ i_5_)  &  (~ i_0_) ) ;
 assign wire7108 = ( (~ i_40_)  &  (~ i_39_)  &  (~ i_35_) ) ;
 assign wire7097 = ( (~ i_7_)  &  (~ i_6_)  &  (~ i_34_) ) ;
 assign wire1522 = ( n_n989  &  n_n983  &  wire445 ) ;
 assign wire7089 = ( n_n977  &  n_n983 ) | ( n_n1023  &  n_n1065 ) ;
 assign wire7090 = ( n_n1066  &  n_n1001 ) | ( n_n976  &  wire121 ) ;
 assign wire1524 = ( n_n1006  &  wire7089 ) | ( n_n1006  &  wire7090 ) ;
 assign wire1525 = ( n_n926  &  n_n1066  &  n_n989 ) ;
 assign wire1539 = ( i_9_  &  (~ i_15_)  &  wire76  &  wire465 ) ;
 assign wire1540 = ( n_n1006  &  n_n1056  &  wire441 ) ;
 assign wire1541 = ( (~ i_12_)  &  (~ i_11_)  &  wire76  &  wire401 ) ;
 assign wire1546 = ( i_40_  &  i_39_  &  (~ i_36_)  &  (~ i_37_) ) ;
 assign wire1547 = ( i_39_  &  (~ i_36_)  &  (~ i_38_)  &  (~ i_37_) ) ;
 assign wire1542 = ( n_n1066  &  n_n989  &  wire1546 ) | ( n_n1066  &  n_n989  &  wire1547 ) ;
 assign wire7073 = ( i_40_  &  (~ i_36_)  &  (~ i_38_) ) ;
 assign wire1548 = ( n_n1066  &  n_n989  &  wire7073 ) ;
 assign wire1550 = ( n_n1074  &  n_n969  &  n_n970 ) ;
 assign wire1551 = ( n_n966  &  n_n1012  &  n_n967 ) ;
 assign wire1552 = ( n_n1074  &  n_n968  &  wire59 ) ;
 assign wire7064 = ( (~ i_40_)  &  (~ i_39_)  &  (~ i_38_)  &  i_37_ ) ;
 assign wire1555 = ( n_n1056  &  n_n1057  &  wire7063  &  wire7064 ) ;
 assign wire1562 = ( (~ n_n1014)  &  n_n1052  &  n_n1057  &  n_n1053 ) ;
 assign wire7067 = ( (~ i_3_)  &  (~ i_4_)  &  wire45 ) ;
 assign wire1557 = ( n_n1067  &  wire1562 ) | ( n_n1067  &  wire797  &  wire7067 ) ;
 assign wire7055 = ( (~ i_12_)  &  (~ i_35_)  &  (~ i_37_) ) | ( (~ i_11_)  &  (~ i_35_)  &  (~ i_37_) ) ;
 assign wire1565 = ( wire76  &  wire7055  &  _9811 ) ;
 assign wire7057 = ( (~ i_14_)  &  i_17_  &  i_16_ ) ;
 assign wire1566 = ( n_n1055  &  n_n1048  &  n_n1047  &  wire7057 ) ;
 assign wire1568 = ( n_n1067  &  n_n1023  &  n_n1065  &  n_n1057 ) ;
 assign wire1577 = ( n_n1055  &  n_n1048  &  n_n1047  &  wire7052 ) ;
 assign wire1578 = ( n_n1073  &  wire76  &  _9825 ) ;
 assign wire7052 = ( i_9_  &  (~ i_12_) ) ;
 assign wire1592 = ( (~ i_22_)  &  wire50  &  wire87  &  wire559 ) ;
 assign wire1620 = ( wire422  &  n_n462  &  n_n801  &  wire375 ) ;
 assign wire7016 = ( i_12_  &  i_16_  &  i_15_ ) ;
 assign wire1624 = ( n_n933  &  n_n1066  &  n_n527  &  wire7016 ) ;
 assign wire7011 = ( i_12_  &  (~ i_11_)  &  i_15_ ) ;
 assign wire1632 = ( n_n1066  &  n_n860  &  n_n927  &  wire7011 ) ;
 assign wire6999 = ( n_n883  &  n_n970 ) | ( n_n969  &  n_n865 ) ;
 assign wire1635 = ( wire555  &  wire6999 ) | ( n_n971  &  n_n1072  &  wire555 ) ;
 assign wire1657 = ( (~ i_18_)  &  wire82 ) | ( (~ i_18_)  &  wire87 ) ;
 assign wire6978 = ( i_12_  &  i_15_  &  n_n793 ) | ( i_11_  &  i_15_  &  n_n793 ) ;
 assign wire6979 = ( n_n791  &  wire6976  &  _9690 ) ;
 assign wire6945 = ( (~ i_39_)  &  (~ i_36_)  &  (~ i_38_)  &  (~ i_37_) ) ;
 assign wire1700 = ( n_n966  &  n_n1012  &  wire6930 ) ;
 assign wire1701 = ( n_n945  &  wire6789  &  wire304 ) ;
 assign wire6930 = ( i_40_  &  i_39_  &  i_22_  &  (~ i_38_) ) ;
 assign wire1704 = ( n_n998  &  n_n973  &  n_n158  &  wire35 ) ;
 assign wire1705 = ( n_n1074  &  n_n330  &  n_n969  &  n_n968 ) ;
 assign wire1707 = ( n_n979  &  n_n978  &  n_n330  &  n_n700 ) ;
 assign wire1708 = ( n_n883  &  n_n998  &  n_n861 ) ;
 assign wire1709 = ( wire50  &  wire6920  &  _9598 ) ;
 assign wire1730 = ( (~ i_7_)  &  wire50  &  wire464  &  n_n1065 ) ;
 assign wire1731 = ( n_n1048  &  n_n1047  &  n_n469  &  wire420 ) ;
 assign wire6890 = ( i_39_  &  (~ i_36_)  &  (~ i_37_) ) ;
 assign wire1741 = ( n_n330  &  n_n1066  &  n_n989  &  wire6890 ) ;
 assign wire1742 = ( n_n979  &  n_n330  &  n_n700  &  wire65 ) ;
 assign wire6874 = ( (~ i_40_)  &  (~ i_36_)  &  i_38_  &  (~ i_37_) ) ;
 assign wire1758 = ( n_n330  &  n_n1066  &  n_n989  &  wire6874 ) ;
 assign wire6842 = ( i_24_  &  i_22_  &  (~ i_19_) ) ;
 assign wire1780 = ( wire512  &  wire614  &  wire6842 ) ;
 assign wire6839 = ( i_24_  &  i_22_  &  (~ i_32_)  &  wire609 ) ;
 assign wire1793 = ( i_11_  &  i_18_  &  (~ i_21_)  &  i_15_ ) ;
 assign wire6841 = ( n_n945  &  wire6789  &  n_n860  &  wire342 ) ;
 assign wire6824 = ( (~ i_39_)  &  (~ i_25_)  &  (~ i_26_)  &  (~ i_38_) ) ;
 assign wire1803 = ( n_n864  &  wire79  &  wire6824 ) ;
 assign wire1804 = ( n_n966  &  n_n1014  &  n_n330  &  n_n993 ) ;
 assign wire1806 = ( n_n1002  &  n_n861  &  n_n710  &  wire100 ) ;
 assign wire1807 = ( n_n709  &  n_n998  &  n_n861  &  n_n710 ) ;
 assign wire1812 = ( wire88  &  n_n997  &  n_n991 ) ;
 assign wire6800 = ( n_n1011  &  n_n1074  &  wire6731  &  wire491 ) ;
 assign wire1821 = ( wire6800  &  _9283 ) | ( wire36  &  wire6800  &  _9284 ) ;
 assign wire1822 = ( n_n1074  &  wire549  &  n_n970 ) ;
 assign wire1832 = ( n_n1072  &  wire42  &  n_n945  &  wire6789 ) ;
 assign wire6801 = ( n_n1011  &  n_n1074  &  wire6731  &  n_n411 ) ;
 assign wire1823 = ( wire48  &  wire1832 ) | ( wire48  &  wire57  &  wire6801 ) ;
 assign wire1839 = ( n_n955  &  _9302 ) | ( n_n955  &  _9303 ) ;
 assign wire1835 = ( wire84  &  wire1839 ) | ( wire84  &  n_n928  &  _9305 ) ;
 assign wire1836 = ( i_12_  &  i_15_  &  wire416  &  n_n928 ) ;
 assign wire6791 = ( n_n945  &  wire6789  &  wire6790 ) ;
 assign wire1845 = ( n_n1048  &  n_n1047  &  (~ wire202)  &  wire458 ) ;
 assign wire1850 = ( n_n979  &  n_n949  &  n_n945 ) | ( n_n979  &  n_n945  &  n_n947 ) ;
 assign wire1847 = ( wire471  &  n_n998  &  wire46  &  wire342 ) ;
 assign wire6780 = ( (~ i_5_)  &  (~ i_32_)  &  (~ i_31_)  &  i_33_ ) ;
 assign wire1860 = ( n_n1002  &  n_n975  &  _9262 ) ;
 assign wire1861 = ( n_n966  &  n_n1012  &  n_n799 ) ;
 assign wire1862 = ( n_n1074  &  wire6731  &  wire120 ) ;
 assign wire1863 = ( n_n966  &  n_n967  &  n_n1073 ) ;
 assign wire1878 = ( n_n966  &  n_n1073  &  wire548 ) ;
 assign wire1871 = ( n_n990  &  n_n861  &  wire94 ) ;
 assign wire1872 = ( wire88  &  n_n1055  &  n_n991 ) ;
 assign wire6766 = ( i_40_  &  i_36_  &  (~ i_38_)  &  i_37_ ) ;
 assign wire6749 = ( i_9_  &  (~ i_5_)  &  i_11_  &  i_15_ ) ;
 assign wire1880 = ( wire45  &  n_n1009  &  wire6749  &  _9057 ) ;
 assign wire6750 = ( i_26_  &  (~ i_38_)  &  (~ i_37_) ) ;
 assign wire1881 = ( (~ i_32_)  &  i_33_  &  n_n1002  &  wire6750 ) ;
 assign wire1882 = ( n_n1074  &  n_n864  &  wire543 ) ;
 assign wire1883 = ( wire363  &  wire1890 ) | ( wire363  &  wire1891 ) | ( wire363  &  wire478 ) ;
 assign wire1884 = ( n_n1074  &  wire66  &  wire6731 ) ;
 assign wire1896 = ( n_n979  &  n_n866  &  n_n907  &  wire6716 ) ;
 assign wire6736 = ( i_25_  &  (~ i_38_)  &  (~ i_37_) ) ;
 assign wire1905 = ( (~ i_32_)  &  i_33_  &  n_n1002  &  wire6736 ) ;
 assign wire1909 = ( wire6739  &  _9110 ) | ( wire6739  &  _9111 ) ;
 assign wire6727 = ( i_12_  &  (~ i_11_)  &  (~ i_32_) ) ;
 assign wire1910 = ( wire325  &  n_n1056  &  wire6727 ) ;
 assign wire6729 = ( (~ i_9_)  &  (~ i_5_)  &  (~ i_16_) ) ;
 assign wire1911 = ( n_n1047  &  wire6728  &  wire6729 ) ;
 assign wire1914 = ( n_n1074  &  n_n970  &  n_n1072 ) ;
 assign wire1926 = ( (~ i_12_)  &  i_11_  &  wire407 ) | ( i_12_  &  (~ i_11_)  &  wire407 ) ;
 assign wire1923 = ( wire363  &  wire1926 ) | ( (~ i_14_)  &  wire363  &  wire686 ) ;
 assign wire1933 = ( n_n979  &  n_n945  &  n_n528  &  wire36 ) ;
 assign wire1935 = ( wire471  &  n_n998  &  wire46  &  wire400 ) ;
 assign wire1936 = ( n_n979  &  n_n907  &  wire6716  &  wire65 ) ;
 assign wire6719 = ( wire1933 ) | ( wire1935 ) | ( wire1936 ) ;
 assign wire6722 = ( n_n1072  &  n_n1073  &  wire670 ) ;
 assign wire6726 = ( _1226 ) | ( _1227 ) ;
 assign wire6746 = ( wire1896 ) | ( n_n907  &  wire6716  &  wire741 ) ;
 assign wire6747 = ( wire6746 ) | ( n_n884  &  wire742 ) ;
 assign wire6753 = ( wire1884 ) | ( n_n1074  &  (~ wire73)  &  wire6722 ) ;
 assign wire6754 = ( wire145 ) | ( wire1881 ) | ( wire1882 ) ;
 assign wire6757 = ( wire6719 ) | ( wire6753 ) | ( _9170 ) ;
 assign wire6764 = ( (~ i_40_)  &  (~ i_39_)  &  n_n985 ) ;
 assign wire6778 = ( wire153 ) | ( wire184 ) | ( wire1860 ) ;
 assign wire6779 = ( wire187 ) | ( wire1861 ) | ( wire1862 ) | ( wire1863 ) ;
 assign wire6786 = ( i_12_  &  (~ i_11_)  &  wire407 ) ;
 assign wire6788 = ( (~ i_12_)  &  i_11_  &  wire407 ) ;
 assign wire6790 = ( i_40_  &  i_39_  &  (~ i_21_)  &  i_38_ ) ;
 assign wire6804 = ( wire145 ) | ( wire241 ) | ( wire1822 ) ;
 assign wire6844 = ( (~ i_17_)  &  (~ i_16_)  &  n_n833 ) ;
 assign wire6845 = ( (~ i_12_)  &  (~ i_31_)  &  wire45  &  wire82 ) ;
 assign wire6849 = ( (~ i_39_)  &  (~ i_38_)  &  i_37_  &  wire94 ) ;
 assign wire6853 = ( n_n785  &  n_n781 ) | ( n_n777  &  wire64 ) ;
 assign wire6854 = ( wire6844  &  wire6845 ) | ( wire106  &  wire6849 ) ;
 assign wire6856 = ( (~ i_9_)  &  (~ i_7_)  &  (~ i_5_)  &  _9411 ) ;
 assign wire6857 = ( (~ i_9_)  &  (~ i_7_)  &  (~ i_5_)  &  _9416 ) ;
 assign wire6860 = ( wire367  &  wire479 ) | ( wire504  &  wire671 ) ;
 assign wire6861 = ( n_n334  &  wire103 ) | ( n_n313  &  wire672 ) ;
 assign wire6863 = ( i_39_  &  (~ i_37_) ) ;
 assign wire6865 = ( i_12_  &  (~ i_18_)  &  i_15_ ) | ( i_11_  &  (~ i_18_)  &  i_15_ ) ;
 assign wire6866 = ( (~ i_9_)  &  (~ i_7_)  &  (~ i_5_)  &  wire6865 ) ;
 assign wire6873 = ( i_21_  &  n_n833 ) ;
 assign wire6877 = ( n_n837  &  wire710 ) | ( wire688  &  wire6873 ) ;
 assign wire6901 = ( wire1730 ) | ( wire422  &  n_n462  &  wire689 ) ;
 assign wire6902 = ( n_n1971 ) | ( wire1731 ) | ( wire711  &  wire429 ) ;
 assign wire6904 = ( n_n1951 ) | ( wire148 ) | ( wire6901 ) | ( wire6902 ) ;
 assign wire6909 = ( wire366  &  wire529 ) | ( wire84  &  wire6856 ) ;
 assign wire6910 = ( wire64  &  n_n771 ) | ( wire84  &  wire6857 ) ;
 assign wire6911 = ( wire386  &  wire132 ) | ( n_n775  &  wire690 ) ;
 assign wire6924 = ( n_n2487 ) | ( n_n2488 ) | ( wire1705 ) | ( wire1708 ) ;
 assign wire6925 = ( wire1704 ) | ( wire1707 ) | ( wire1709 ) ;
 assign wire6927 = ( wire6924 ) | ( wire6925 ) | ( _1045 ) | ( _1046 ) ;
 assign wire6932 = ( n_n469  &  n_n945  &  wire6789 ) ;
 assign wire6948 = ( (~ i_22_)  &  wire82 ) ;
 assign wire6960 = ( n_n862  &  n_n1064  &  wire529 ) | ( n_n862  &  n_n1064  &  wire535 ) ;
 assign wire6961 = ( (~ i_40_)  &  (~ i_38_)  &  wire542 ) | ( (~ i_39_)  &  (~ i_38_)  &  wire542 ) ;
 assign wire6969 = ( (~ i_34_)  &  (~ i_36_)  &  i_35_  &  _9680 ) ;
 assign wire6975 = ( (~ i_39_)  &  (~ i_38_)  &  i_37_  &  wire94 ) ;
 assign wire6980 = ( (~ i_34_)  &  (~ i_36_)  &  i_35_  &  _9700 ) ;
 assign wire6985 = ( n_n1971 ) | ( n_n2487 ) | ( n_n2488 ) ;
 assign wire6993 = ( n_n865  &  _9723 ) | ( n_n865  &  _9724 ) ;
 assign wire7001 = ( n_n1951 ) | ( _968 ) ;
 assign wire7002 = ( wire80  &  n_n926  &  _9533 ) | ( wire80  &  n_n926  &  _9535 ) ;
 assign wire7014 = ( i_9_  &  (~ i_7_)  &  (~ i_5_)  &  i_15_ ) ;
 assign wire7020 = ( n_n998  &  n_n861  &  wire325 ) | ( n_n998  &  n_n861  &  wire556 ) ;
 assign wire7033 = ( wire329  &  wire337 ) | ( (~ i_22_)  &  wire87  &  wire337 ) ;
 assign wire7034 = ( n_n761  &  wire323 ) | ( (~ i_23_)  &  wire323  &  wire370 ) ;
 assign wire7035 = ( wire175 ) | ( wire240 ) ;
 assign wire7038 = ( wire1592 ) | ( wire7033 ) | ( wire7034 ) | ( wire7035 ) ;
 assign wire7044 = ( (~ i_34_)  &  (~ i_36_) ) ;
 assign wire7066 = ( i_9_  &  (~ i_11_) ) ;
 assign wire7069 = ( wire1555 ) | ( n_n1074  &  (~ wire73)  &  wire6722 ) ;
 assign wire7077 = ( wire1548 ) | ( wire1550 ) | ( wire1551 ) | ( wire1552 ) ;
 assign wire7079 = ( i_40_  &  i_6_ ) ;
 assign wire7086 = ( wire1542 ) | ( _856 ) | ( _857 ) ;
 assign wire7087 = ( wire158 ) | ( wire1539 ) | ( wire1540 ) | ( wire1541 ) ;
 assign wire7092 = ( wire1522 ) | ( wire1525 ) | ( n_n980  &  wire560 ) ;
 assign wire7100 = ( (~ i_7_)  &  (~ i_6_)  &  (~ i_34_) ) ;
 assign wire7102 = ( (~ i_34_)  &  i_36_  &  i_37_ ) ;
 assign wire7123 = ( (~ i_28_)  &  (~ i_29_)  &  n_n985  &  wire7121 ) ;
 assign wire7125 = ( i_15_  &  wire1834 ) | ( i_18_  &  i_15_  &  wire42 ) ;
 assign wire7130 = ( i_9_  &  (~ i_5_)  &  (~ i_14_) ) ;
 assign wire7131 = ( n_n1066  &  n_n927  &  wire7130 ) ;
 assign wire7135 = ( wire361  &  wire7123 ) | ( wire777  &  wire7131 ) ;
 assign wire7137 = ( wire333  &  wire36 ) | ( wire92  &  wire461 ) ;
 assign wire7143 = ( wire1468 ) | ( n_n907  &  wire6716  &  wire782 ) ;
 assign wire7151 = ( i_9_  &  (~ i_5_)  &  n_n933  &  n_n1066 ) ;
 assign wire7153 = ( _768 ) | ( wire786  &  wire7151 ) ;
 assign wire7160 = ( _775 ) | ( n_n1074  &  n_n969  &  n_n970 ) ;
 assign wire7161 = ( wire241 ) | ( wire187 ) | ( wire1453 ) | ( wire1454 ) ;
 assign wire7170 = ( wire184 ) | ( wire1442 ) | ( wire1444 ) ;
 assign wire7178 = ( (~ i_34_)  &  (~ i_35_)  &  (~ i_37_) ) ;
 assign wire7180 = ( n_n1048  &  n_n977  &  wire7178 ) ;
 assign wire7184 = ( wire1415 ) | ( wire1417 ) | ( wire814  &  wire7180 ) ;
 assign wire7185 = ( wire1466 ) | ( wire1467 ) | ( wire7143 ) | ( wire7184 ) ;
 assign wire7189 = ( o_15_ ) | ( n_n966  &  n_n862  &  n_n1064 ) ;
 assign wire7208 = ( wire59  &  wire1388 ) | ( wire59  &  wire1389 ) ;
 assign wire7218 = ( wire1372 ) | ( wire7197  &  _10120 ) ;
 assign wire7219 = ( wire1374 ) | ( n_n1047  &  wire7214  &  _10125 ) ;
 assign wire7220 = ( wire183 ) | ( wire251 ) | ( wire1375 ) ;
 assign wire7230 = ( wire1366 ) | ( _10182 ) | ( n_n1073  &  _10181 ) ;
 assign wire7233 = ( (~ i_40_)  &  i_36_  &  (~ i_35_) ) ;
 assign wire7245 = ( wire303 ) | ( wire1346 ) | ( wire1347 ) | ( wire1348 ) ;
 assign wire7252 = ( wire336 ) | ( wire1340 ) | ( wire1341 ) | ( wire1342 ) ;
 assign wire7263 = ( (~ i_34_)  &  (~ i_35_)  &  i_38_ ) ;
 assign wire7265 = ( i_7_  &  i_33_ ) | ( n_n1047  &  wire6728 ) ;
 assign wire7266 = ( n_n1047  &  n_n980 ) | ( n_n980  &  wire7263 ) ;
 assign wire7269 = ( wire1316 ) | ( wire1317 ) | ( wire7265 ) | ( wire7266 ) ;
 assign wire7284 = ( wire1307 ) | ( wire47  &  wire320  &  wire761 ) ;
 assign wire7285 = ( n_n2213 ) | ( wire1306 ) | ( wire1309 ) ;
 assign wire7286 = ( wire1305 ) | ( _625 ) | ( _626 ) ;
 assign wire7293 = ( wire1294 ) | ( n_n1052  &  wire762 ) ;
 assign wire7299 = ( wire1286 ) | ( _620 ) | ( _621 ) ;
 assign wire7304 = ( i_23_  &  i_24_  &  n_n833 ) ;
 assign wire7305 = ( wire50  &  wire35  &  n_n848 ) ;
 assign wire7306 = ( i_15_  &  (~ i_34_)  &  i_33_ ) ;
 assign wire7317 = ( (~ i_39_)  &  (~ i_38_)  &  n_n888 ) ;
 assign wire7333 = ( i_39_  &  i_37_ ) ;
 assign wire7336 = ( n_n2439 ) | ( wire1257 ) | ( wire1262 ) ;
 assign wire7337 = ( wire1253 ) | ( wire1255 ) | ( wire1256 ) ;
 assign wire7339 = ( i_36_  &  wire1251 ) | ( i_36_  &  wire1252 ) ;
 assign wire7341 = ( n_n1777 ) | ( (~ i_7_)  &  wire45  &  wire7339 ) ;
 assign wire7343 = ( wire1238 ) | ( n_n1047  &  _10358 ) ;
 assign wire7344 = ( wire1254 ) | ( wire7336 ) | ( wire7337 ) | ( wire7343 ) ;
 assign wire7348 = ( n_n979  &  wire35  &  n_n848 ) ;
 assign wire7349 = ( i_9_  &  (~ i_7_)  &  (~ i_5_)  &  (~ i_21_) ) ;
 assign wire7353 = ( (~ i_40_)  &  (~ i_38_)  &  wire542 ) | ( (~ i_39_)  &  (~ i_38_)  &  wire542 ) ;
 assign wire7354 = ( n_n1986 ) | ( wire240 ) ;
 assign wire7355 = ( wire245 ) | ( n_n469  &  wire7347  &  wire7348 ) ;
 assign wire7356 = ( n_n1971 ) | ( wire1230 ) | ( _573 ) ;
 assign wire7373 = ( n_n2487 ) | ( n_n2488 ) | ( n_n1990 ) ;
 assign wire7377 = ( n_n862  &  n_n1064  &  wire529 ) | ( n_n862  &  n_n1064  &  wire535 ) ;
 assign wire7378 = ( wire175 ) | ( (~ i_40_)  &  (~ i_38_)  &  wire542 ) ;
 assign wire7411 = ( wire1186 ) | ( wire1189 ) | ( wire406  &  wire467 ) ;
 assign wire7416 = ( (~ i_39_)  &  (~ i_38_)  &  n_n1012  &  wire76 ) ;
 assign wire7420 = ( (~ i_17_)  &  (~ i_16_)  &  wire76 ) ;
 assign wire7421 = ( n_n1072  &  n_n1073  &  wire36 ) ;
 assign wire7423 = ( (~ i_40_)  &  i_38_  &  n_n1073 ) ;
 assign wire7428 = ( i_39_  &  (~ i_36_)  &  (~ i_35_)  &  i_38_ ) ;
 assign wire7430 = ( wire1164 ) | ( wire1165 ) | ( n_n475  &  wire617 ) ;
 assign wire7440 = ( wire1156 ) | ( n_n998  &  wire46  &  wire676 ) ;
 assign wire7441 = ( (~ i_9_)  &  (~ i_5_)  &  wire76 ) ;
 assign wire7442 = ( (~ i_40_)  &  i_36_  &  (~ i_38_)  &  i_37_ ) ;
 assign wire7446 = ( _488 ) | ( n_n1055  &  n_n998  &  _10542 ) ;
 assign wire7450 = ( (~ i_21_)  &  i_15_  &  n_n850  &  wire822 ) ;
 assign wire7456 = ( (~ i_21_)  &  i_15_  &  n_n853  &  wire572 ) ;
 assign wire7458 = ( n_n1971 ) | ( wire48  &  n_n850  &  wire337 ) ;
 assign wire7459 = ( wire365  &  wire337 ) | ( (~ i_22_)  &  wire87  &  wire337 ) ;
 assign wire7460 = ( wire337  &  wire6948 ) | ( wire99  &  wire7456 ) ;
 assign wire7476 = ( (~ i_7_)  &  i_31_  &  wire45 ) ;
 assign wire7487 = ( wire1089 ) | ( wire1090 ) | ( wire1091 ) ;
 assign wire7488 = ( i_9_  &  (~ i_7_)  &  n_n1055  &  n_n1047 ) ;
 assign wire7493 = ( wire1075 ) | ( wire400  &  wire737  &  _10643 ) ;
 assign wire7494 = ( wire7487 ) | ( _430 ) | ( _431 ) | ( _10634 ) ;
 assign wire7495 = ( wire1083 ) | ( wire7493 ) | ( wire692  &  wire7488 ) ;
 assign wire7504 = ( wire182 ) | ( wire301 ) | ( wire1049 ) | ( wire1051 ) ;
 assign wire7506 = ( wire1050 ) | ( wire1112 ) | ( wire1113 ) | ( wire7504 ) ;
 assign wire7518 = ( n_n982  &  n_n998  &  n_n861 ) | ( n_n998  &  n_n861  &  wire325 ) ;
 assign wire7523 = ( i_7_  &  i_33_ ) | ( wire84  &  wire6786 ) ;
 assign wire7524 = ( wire84  &  wire6788 ) | ( wire361  &  wire7123 ) ;
 assign wire7535 = ( (~ i_12_)  &  i_11_  &  wire407  &  wire84 ) | ( i_12_  &  (~ i_11_)  &  wire407  &  wire84 ) ;
 assign wire7538 = ( wire146 ) | ( wire153 ) | ( wire1008 ) | ( wire1010 ) ;
 assign wire7542 = ( i_40_  &  i_39_  &  i_38_  &  n_n968 ) | ( (~ i_40_)  &  (~ i_39_)  &  (~ i_38_)  &  n_n968 ) ;
 assign wire7544 = ( wire333  &  wire581 ) | ( wire583  &  wire7542 ) ;
 assign wire7545 = ( wire473  &  wire7125 ) | ( i_19_  &  wire473  &  wire739 ) ;
 assign wire7554 = ( n_n2439 ) | ( wire985 ) | ( wire987 ) | ( wire988 ) ;
 assign wire7555 = ( wire80  &  n_n926  &  _9533 ) | ( wire80  &  n_n926  &  _9543 ) ;
 assign wire7558 = ( (~ i_23_)  &  n_n469 ) ;
 assign wire7562 = ( (~ i_7_)  &  (~ i_5_)  &  i_12_  &  _10772 ) ;
 assign wire7563 = ( (~ i_40_)  &  (~ i_39_)  &  n_n1009  &  wire422 ) ;
 assign wire7564 = ( i_40_  &  (~ i_39_)  &  n_n1052 ) ;
 assign wire7565 = ( _320 ) | ( n_n862  &  wire529  &  _9615 ) ;
 assign wire7566 = ( wire432  &  wire7562 ) | ( wire408  &  wire7563 ) ;
 assign wire7568 = ( n_n334  &  n_n560 ) | ( n_n525  &  wire7564 ) ;
 assign wire7576 = ( (~ i_7_)  &  (~ i_5_)  &  i_11_  &  _10818 ) ;
 assign wire7588 = ( n_n791  &  wire6976  &  _10837 ) ;
 assign wire7590 = ( wire648  &  wire646 ) | ( wire486  &  wire7588 ) ;
 assign wire7591 = ( wire942 ) | ( wire7590 ) | ( n_n771  &  wire356 ) ;
 assign wire7596 = ( n_n2487 ) | ( n_n2488 ) | ( wire937 ) ;
 assign wire7597 = ( wire940 ) | ( (~ i_36_)  &  wire68  &  n_n329 ) ;
 assign wire7612 = ( wire244 ) | ( wire911 ) | ( n_n334  &  wire103 ) ;
 assign wire7614 = ( wire939 ) | ( wire7596 ) | ( wire7597 ) | ( wire7612 ) ;
 assign wire7625 = ( n_n2836 ) | ( n_n1958 ) | ( n_n1956 ) | ( wire906 ) ;
 assign wire7636 = ( wire890 ) | ( wire894 ) | ( wire7554 ) | ( _10890 ) ;
 assign wire7641 = ( (~ i_39_)  &  (~ i_38_)  &  n_n888 ) ;
 assign wire7645 = ( i_40_  &  i_38_  &  (~ i_37_) ) ;
 assign wire7646 = ( i_11_  &  i_15_  &  wire7645 ) ;
 assign wire7658 = ( wire131 ) | ( n_n2439 ) | ( wire1262 ) ;
 assign wire7659 = ( wire864 ) | ( wire865 ) | ( n_n795  &  wire752 ) ;
 assign wire7661 = ( (~ i_31_)  &  wire45  &  n_n462 ) ;
 assign wire7663 = ( wire860 ) | ( _207 ) | ( _208 ) ;
 assign wire7664 = ( wire244 ) | ( wire859 ) | ( wire102  &  wire7661 ) ;
 assign wire7666 = ( wire357  &  n_n329 ) | ( n_n334  &  n_n560 ) ;
 assign wire7667 = ( wire850 ) | ( _213 ) | ( _214 ) ;
 assign wire7673 = ( wire519 ) | ( wire533 ) | ( wire538 ) ;
 assign wire7676 = ( (~ i_34_)  &  (~ i_36_)  &  i_35_  &  _11002 ) ;
 assign wire7677 = ( n_n966  &  n_n1012  &  n_n973 ) ;
 assign wire7680 = ( wire587  &  wire7676 ) | ( wire364  &  wire7677 ) ;
 assign wire7681 = ( wire7680 ) | ( i_38_  &  (~ i_37_)  &  wire586 ) ;
 assign wire7704 = ( wire154 ) | ( wire309 ) | ( wire310 ) | ( wire312 ) ;
 assign wire7722 = ( (~ i_18_)  &  (~ i_21_)  &  i_15_ ) ;
 assign wire7728 = ( wire276 ) | ( wire303  &  wire655  &  wire7722 ) ;
 assign wire7734 = ( o_15_ ) | ( n_n1074  &  n_n1021  &  wire664 ) ;
 assign wire7747 = ( wire248 ) | ( wire250 ) | ( wire252 ) ;
 assign wire7754 = ( wire153 ) | ( wire229 ) | ( wire232 ) | ( wire235 ) ;
 assign wire7755 = ( wire231 ) | ( wire234 ) | ( wire403  &  wire684 ) ;
 assign wire7757 = ( i_40_  &  i_39_  &  i_36_  &  i_38_ ) ;
 assign wire7761 = ( wire217 ) | ( _124 ) | ( _125 ) ;
 assign wire7762 = ( wire218 ) | ( wire7754 ) | ( wire7755 ) ;
 assign wire7791 = ( wire188 ) | ( wire190 ) | ( wire193 ) ;
 assign wire7811 = ( wire142 ) | ( wire143 ) | ( wire151 ) ;
 assign wire7814 = ( wire144 ) | ( wire7811 ) | ( _35 ) | ( _38 ) ;
 assign _35 = ( wire47  &  wire160 ) | ( wire47  &  _40 ) | ( wire47  &  _41 ) ;
 assign _38 = ( (~ i_39_)  &  wire45  &  n_n1061  &  _10987 ) ;
 assign _40 = ( wire7809  &  wire163 ) | ( wire7809  &  wire164 ) ;
 assign _41 = ( wire7809  &  wire162 ) | ( wire7809  &  _43 ) | ( wire7809  &  _44 ) ;
 assign _43 = ( (~ i_39_)  &  (~ i_36_)  &  (~ i_35_)  &  i_38_ ) ;
 assign _44 = ( (~ i_40_)  &  (~ i_36_)  &  (~ i_35_)  &  i_38_ ) ;
 assign _46 = ( n_n795  &  n_n861  &  wire613 ) | ( n_n795  &  n_n861  &  _11261 ) ;
 assign _53 = ( wire7816  &  wire70  &  _11241 ) ;
 assign _54 = ( wire7816  &  _56 ) | ( wire7816  &  _57 ) ;
 assign _56 = ( wire35  &  n_n945  &  wire6789  &  _11244 ) ;
 assign _57 = ( n_n945  &  wire6789  &  wire7815  &  _11249 ) ;
 assign _60 = ( n_n775  &  _66 ) | ( n_n775  &  n_n860  &  wire104 ) ;
 assign _61 = ( n_n1047  &  wire840  &  wire7817  &  _9420 ) ;
 assign _63 = ( n_n785  &  _66 ) | ( n_n785  &  n_n860  &  wire104 ) ;
 assign _66 = ( n_n860  &  wire38  &  wire7011 ) ;
 assign _78 = ( n_n1074  &  n_n978  &  n_n968  &  _11201 ) ;
 assign _79 = ( n_n1074  &  n_n978  &  n_n968  &  wire420 ) ;
 assign _86 = ( n_n1012  &  wire662  &  _9322 ) ;
 assign _101 = ( n_n985  &  n_n874  &  wire7760  &  _11145 ) ;
 assign _105 = ( n_n1074  &  n_n710  &  n_n1065  &  _11128 ) ;
 assign _110 = ( n_n979  &  n_n1001  &  n_n947  &  wire7399 ) ;
 assign _111 = ( n_n979  &  n_n1001  &  n_n947  &  wire7390 ) ;
 assign _112 = ( n_n979  &  n_n949  &  n_n1001  &  wire7405 ) ;
 assign _113 = ( n_n979  &  n_n969  &  n_n949  &  wire7406 ) ;
 assign _114 = ( n_n979  &  n_n969  &  n_n947  &  wire7390 ) ;
 assign _115 = ( n_n998  &  n_n866  &  wire633  &  _11119 ) ;
 assign _116 = ( n_n977  &  n_n888  &  wire633  &  wire7694 ) ;
 assign _119 = ( n_n979  &  n_n949  &  wire81  &  wire7406 ) ;
 assign _120 = ( n_n979  &  n_n947  &  wire81  &  wire7390 ) ;
 assign _122 = ( n_n979  &  n_n947  &  wire7399  &  _11107 ) ;
 assign _123 = ( n_n979  &  n_n949  &  wire7405  &  _11109 ) ;
 assign _124 = ( n_n1066  &  wire7757  &  _11094 ) | ( n_n1066  &  wire7757  &  _11095 ) ;
 assign _125 = ( n_n1066  &  wire7757  &  _10436 ) | ( n_n1066  &  wire7757  &  _10437 ) ;
 assign _129 = ( wire45  &  n_n973  &  wire7745 ) ;
 assign _130 = ( i_30_  &  (~ i_5_)  &  wire45  &  n_n462 ) ;
 assign _131 = ( wire45  &  wire7743  &  _11079 ) | ( wire45  &  wire7743  &  _11080 ) ;
 assign _132 = ( n_n1066  &  n_n453  &  wire7743 ) | ( n_n1066  &  n_n458  &  wire7743 ) ;
 assign _145 = ( i_39_  &  wire45  &  _9118 ) ;
 assign _148 = ( (~ i_37_)  &  wire45  &  _9118 ) ;
 assign _149 = ( i_38_  &  wire45  &  _9118 ) ;
 assign _158 = ( wire520  &  _11046 ) ;
 assign _159 = ( i_15_  &  _162 ) | ( i_15_  &  _163 ) ;
 assign _162 = ( (~ i_16_)  &  wire445  &  n_n488  &  wire421 ) ;
 assign _163 = ( (~ i_17_)  &  wire45  &  n_n926  &  n_n488 ) ;
 assign _165 = ( n_n979  &  n_n969  &  n_n947  &  n_n791 ) ;
 assign _172 = ( n_n843  &  n_n1057  &  n_n1053  &  wire299 ) ;
 assign _173 = ( n_n843  &  n_n1057  &  n_n1053  &  n_n836 ) ;
 assign _175 = ( wire45  &  n_n492  &  n_n918  &  _11018 ) ;
 assign _176 = ( wire45  &  n_n985  &  n_n488  &  _11020 ) ;
 assign _177 = ( wire45  &  n_n947  &  n_n923  &  _11022 ) ;
 assign _193 = ( wire45  &  n_n1061  &  _10987  &  _10989 ) ;
 assign _195 = ( n_n969  &  n_n888  &  n_n700  &  wire7276 ) ;
 assign _196 = ( n_n330  &  n_n888  &  n_n700  &  _10982 ) ;
 assign _207 = ( n_n330  &  n_n1066  &  n_n989  &  wire1547 ) ;
 assign _208 = ( n_n330  &  n_n1066  &  n_n989  &  wire1546 ) ;
 assign _213 = ( (~ i_13_)  &  wire50  &  wire315  &  wire304 ) ;
 assign _214 = ( (~ i_13_)  &  wire50  &  n_n833  &  wire315 ) ;
 assign _218 = ( wire45  &  wire315  &  _10941 ) ;
 assign _219 = ( wire80  &  wire315  &  _10943 ) ;
 assign _221 = ( wire845  &  _10935 ) | ( _223  &  _10935 ) | ( _224  &  _10935 ) ;
 assign _223 = ( (~ i_7_)  &  (~ i_5_)  &  wire7122  &  _10931 ) ;
 assign _224 = ( (~ i_7_)  &  (~ i_5_)  &  wire45  &  _10933 ) ;
 assign _226 = ( wire7649  &  _231 ) | ( wire44  &  wire7649  &  wire7648 ) ;
 assign _231 = ( n_n411  &  wire1798  &  _10927 ) | ( n_n411  &  _10925  &  _10927 ) ;
 assign _245 = ( n_n1074  &  wire6828  &  wire402 ) | ( n_n1074  &  wire402  &  _10899 ) ;
 assign _250 = ( wire6828  &  wire7630  &  _9558 ) ;
 assign _294 = ( wire325  &  n_n976  &  wire315  &  _10810 ) ;
 assign _295 = ( n_n330  &  n_n989  &  wire445  &  n_n976 ) ;
 assign _297 = ( n_n861  &  n_n710  &  n_n715  &  _10803 ) ;
 assign _320 = ( n_n865  &  n_n843  &  _9179  &  _9806 ) ;
 assign _334 = ( (~ i_22_)  &  wire80  &  wire82  &  wire7145 ) ;
 assign _335 = ( (~ i_22_)  &  wire80  &  wire87  &  wire7145 ) ;
 assign _380 = ( wire1048  &  _10691 ) | ( _384  &  _10691 ) | ( _385  &  _10691 ) ;
 assign _381 = ( wire1046  &  wire7511 ) ;
 assign _384 = ( (~ i_32_)  &  n_n1009  &  n_n1023  &  _9737 ) ;
 assign _385 = ( (~ i_32_)  &  n_n985  &  n_n1023  &  _9445 ) ;
 assign _387 = ( i_20_  &  i_21_  &  wire303  &  _10678 ) ;
 assign _406 = ( n_n985  &  n_n629  &  n_n874  &  _9086 ) ;
 assign _407 = ( n_n1074  &  n_n968  &  n_n629  &  _9131 ) ;
 assign _408 = ( n_n1074  &  n_n1012  &  n_n629  &  _9032 ) ;
 assign _409 = ( (~ i_15_)  &  wire50  &  n_n1052  &  _10651 ) ;
 assign _410 = ( (~ i_15_)  &  wire45  &  n_n1009  &  _10653 ) ;
 assign _430 = ( n_n1001  &  wire38  &  _10613  &  _10615 ) ;
 assign _431 = ( n_n977  &  wire79  &  n_n1073  &  _10617 ) ;
 assign _435 = ( (~ i_7_)  &  (~ i_15_)  &  wire45  &  wire792 ) ;
 assign _440 = ( (~ i_40_)  &  n_n685  &  n_n1074  &  n_n923 ) ;
 assign _441 = ( (~ i_40_)  &  n_n685  &  n_n1052  &  n_n874 ) ;
 assign _452 = ( (~ i_7_)  &  (~ i_15_)  &  wire50  &  n_n833 ) ;
 assign _453 = ( (~ i_15_)  &  _456 ) | ( (~ i_15_)  &  wire715  &  _10584 ) ;
 assign _456 = ( i_40_  &  (~ i_7_)  &  wire45  &  n_n836 ) ;
 assign _479 = ( wire82  &  n_n968  &  wire7452  &  _10552 ) ;
 assign _485 = ( wire87  &  n_n968  &  wire7452  &  _10552 ) ;
 assign _488 = ( i_7_  &  i_33_ ) ;
 assign _494 = ( n_n1023  &  wire681  &  wire7442 ) | ( n_n1023  &  wire7442  &  _10525 ) ;
 assign _512 = ( wire330  &  n_n998  &  n_n949  &  _10507 ) ;
 assign _513 = ( wire330  &  n_n998  &  n_n949  &  n_n791 ) ;
 assign _524 = ( n_n492  &  wire76  &  wire465  &  _10483 ) ;
 assign _525 = ( n_n492  &  wire76  &  wire401  &  _10483 ) ;
 assign _547 = ( wire330  &  n_n998  &  n_n947  &  _10421 ) ;
 assign _554 = ( (~ i_24_)  &  wire50  &  wire82  &  wire54 ) ;
 assign _555 = ( (~ i_24_)  &  wire50  &  wire82  &  wire371 ) ;
 assign _567 = ( n_n842  &  n_n865  &  n_n843  &  _9179 ) ;
 assign _573 = ( n_n865  &  n_n843  &  _9179  &  _9806 ) ;
 assign _593 = ( n_n861  &  n_n991  &  wire767 ) | ( n_n861  &  n_n991  &  _10339 ) ;
 assign _618 = ( wire50  &  wire35  &  n_n528  &  _10305 ) ;
 assign _619 = ( (~ i_13_)  &  wire50  &  n_n528  &  wire315 ) ;
 assign _620 = ( n_n883  &  n_n1047  &  wire1291  &  _10296 ) ;
 assign _621 = ( n_n883  &  n_n1047  &  wire43  &  _10296 ) ;
 assign _625 = ( n_n1012  &  wire488  &  wire7281  &  _10285 ) ;
 assign _626 = ( n_n1047  &  wire488  &  wire494  &  wire7279 ) ;
 assign _713 = ( n_n1047  &  wire7194  &  _10114 ) ;
 assign _714 = ( n_n1047  &  wire7193  &  _10114 ) ;
 assign _722 = ( n_n1047  &  n_n973  &  wire7201  &  _10085 ) ;
 assign _725 = ( n_n1047  &  wire7200  &  wire788  &  _10089 ) ;
 assign _731 = ( (~ i_38_)  &  (~ i_37_)  &  _742 ) | ( (~ i_38_)  &  (~ i_37_)  &  _10093 ) ;
 assign _733 = ( n_n1047  &  n_n967  &  wire7201  &  _10085 ) ;
 assign _742 = ( n_n1047  &  wire1400  &  _10089 ) | ( n_n1047  &  _743  &  _10089 ) ;
 assign _743 = ( i_11_  &  i_16_  &  i_15_ ) ;
 assign _745 = ( i_32_  &  (~ i_33_) ) ;
 assign _765 = ( n_n1067  &  n_n1052  &  n_n1057  &  n_n1053 ) ;
 assign _766 = ( n_n1067  &  n_n1023  &  n_n1065  &  n_n1057 ) ;
 assign _768 = ( n_n926  &  n_n1066  &  wire7132  &  _9971 ) ;
 assign _772 = ( n_n1066  &  n_n928  &  n_n923  &  n_n927 ) ;
 assign _775 = ( n_n1074  &  n_n967  &  n_n968 ) ;
 assign _781 = ( n_n1074  &  n_n969  &  n_n884  &  _10011 ) ;
 assign _782 = ( n_n1074  &  n_n968  &  n_n884  &  _9131 ) ;
 assign _783 = ( n_n1074  &  wire6731  &  n_n978  &  n_n884 ) ;
 assign _785 = ( n_n1012  &  wire76  &  _10009 ) ;
 assign _788 = ( i_40_  &  _791 ) | ( i_40_  &  _792 ) ;
 assign _789 = ( i_40_  &  n_n993  &  wire76  &  _9983 ) ;
 assign _790 = ( i_40_  &  n_n991  &  wire7165  &  _9987 ) ;
 assign _791 = ( i_6_  &  n_n998  &  _9980 ) ;
 assign _792 = ( i_6_  &  n_n1002  &  _9982 ) ;
 assign _805 = ( n_n937  &  wire6907  &  _9425 ) ;
 assign _808 = ( n_n926  &  n_n1066  &  n_n927  &  wire63 ) ;
 assign _809 = ( n_n926  &  n_n933  &  n_n1066  &  n_n928 ) ;
 assign _835 = ( (~ i_7_)  &  _838 ) | ( (~ i_7_)  &  wire7108  &  _9914 ) ;
 assign _836 = ( (~ i_7_)  &  n_n1012  &  n_n1072  &  _9917 ) ;
 assign _838 = ( i_32_  &  (~ i_34_)  &  i_36_ ) | ( i_32_  &  (~ i_34_)  &  i_35_ ) | ( i_32_  &  i_34_  &  (~ i_36_)  &  (~ i_35_) ) ;
 assign _848 = ( (~ i_0_)  &  n_n969  &  n_n865  &  _9905 ) ;
 assign _849 = ( (~ i_0_)  &  n_n991  &  wire400  &  _9907 ) ;
 assign _856 = ( n_n998  &  n_n997  &  wire7079  &  _9879 ) ;
 assign _857 = ( n_n1002  &  wire820  &  wire7079  &  _9883 ) ;
 assign _881 = ( n_n1048  &  n_n1047  &  wire7066  &  _9306 ) ;
 assign _892 = ( i_9_  &  (~ i_14_)  &  i_17_ ) | ( i_9_  &  (~ i_11_)  &  i_17_ ) ;
 assign _893 = ( (~ i_12_)  &  i_17_  &  i_16_ ) | ( (~ i_11_)  &  i_17_  &  i_16_ ) ;
 assign _915 = ( n_n865  &  n_n843  &  _9179  &  _9806 ) ;
 assign _943 = ( n_n1009  &  wire50  &  wire82  &  _9774 ) ;
 assign _954 = ( n_n926  &  wire1624 ) | ( n_n926  &  wire558  &  _9762 ) ;
 assign _959 = ( n_n1009  &  wire1632  &  _9741 ) | ( n_n1009  &  _962  &  _9741 ) ;
 assign _960 = ( n_n1009  &  wire729  &  _9741  &  _9752 ) ;
 assign _962 = ( n_n1066  &  wire78  &  n_n527  &  _9747 ) ;
 assign _968 = ( i_0_  &  wire79  &  n_n1072  &  _9483 ) ;
 assign _970 = ( wire88  &  n_n975  &  wire6938 ) ;
 assign _979 = ( i_0_  &  wire79  &  n_n970  &  _9479 ) ;
 assign _982 = ( n_n685  &  wire6991  &  n_n998  &  _9718 ) ;
 assign _983 = ( n_n685  &  wire6991  &  n_n1002  &  _9721 ) ;
 assign _984 = ( n_n842  &  n_n865  &  n_n843  &  _9179 ) ;
 assign _1021 = ( n_n1009  &  wire50  &  wire87  &  _9636 ) ;
 assign _1045 = ( wire79  &  n_n865  &  wire373  &  _9580 ) ;
 assign _1046 = ( wire6897  &  n_n865  &  wire373  &  _9527 ) ;
 assign _1052 = ( wire79  &  n_n865  &  wire373  &  _9555 ) ;
 assign _1053 = ( wire6828  &  n_n865  &  wire373  &  _9558 ) ;
 assign _1063 = ( i_0_  &  wire79  &  n_n1072  &  _9483 ) ;
 assign _1065 = ( i_0_  &  wire79  &  n_n970  &  _9479 ) ;
 assign _1075 = ( (~ i_23_)  &  wire70  &  wire6841 ) | ( (~ i_23_)  &  wire1793  &  wire6841 ) ;
 assign _1076 = ( (~ i_23_)  &  n_n952  &  wire6839  &  _9451 ) ;
 assign _1080 = ( i_12_  &  i_18_  &  (~ i_21_)  &  i_15_ ) ;
 assign _1081 = ( i_11_  &  (~ i_21_)  &  i_15_  &  i_19_ ) ;
 assign _1171 = ( wire330  &  n_n1002  &  n_n861 ) ;
 assign _1174 = ( (~ i_7_)  &  i_6_  &  wire50  &  wire6766 ) ;
 assign _1178 = ( n_n842  &  n_n1067  &  n_n865  &  _9179 ) ;
 assign _1204 = ( wire45  &  (~ n_n1055)  &  _9118 ) ;
 assign _1213 = ( n_n966  &  n_n969  &  n_n971 ) ;
 assign _1215 = ( n_n1074  &  wire6731  &  n_n884  &  _9080 ) ;
 assign _1216 = ( n_n1009  &  n_n874  &  n_n884  &  _9083 ) ;
 assign _1217 = ( n_n985  &  n_n874  &  n_n884  &  _9086 ) ;
 assign _1218 = ( (~ i_5_)  &  i_31_  &  wire445  &  wire421 ) ;
 assign _1219 = ( (~ i_5_)  &  n_n1047  &  wire55  &  wire6728 ) ;
 assign _1226 = ( wire45  &  n_n1009  &  wire36  &  _9052 ) ;
 assign _1227 = ( wire45  &  n_n1009  &  wire484  &  _9057 ) ;
 assign _9032 = ( (~ i_38_)  &  (~ i_39_) ) ;
 assign _9036 = ( (~ i_12_)  &  i_16_  &  i_15_ ) ;
 assign _9039 = ( i_12_  &  i_17_  &  i_15_ ) | ( i_12_  &  i_16_  &  i_15_ ) ;
 assign _9041 = ( (~ i_12_)  &  i_17_  &  i_15_ ) ;
 assign _9052 = ( i_40_  &  i_39_  &  i_17_  &  i_16_ ) ;
 assign _9057 = ( i_40_  &  i_39_  &  i_17_ ) | ( i_40_  &  i_39_  &  i_16_ ) ;
 assign _9080 = ( (~ i_38_)  &  i_40_ ) ;
 assign _9083 = ( (~ i_39_)  &  (~ i_40_) ) ;
 assign _9086 = ( i_39_  &  i_40_ ) ;
 assign _9110 = ( (~ i_15_)  &  (~ i_32_)  &  (~ i_34_)  &  i_33_ ) ;
 assign _9111 = ( (~ i_12_)  &  (~ i_32_)  &  (~ i_34_)  &  i_33_ ) ;
 assign _9118 = ( (~ i_5_)  &  i_31_  &  (~ i_36_) ) ;
 assign _9119 = ( wire1905 ) | ( _1204 ) | ( _1213 ) ;
 assign _9131 = ( i_38_  &  i_39_ ) ;
 assign _9170 = ( wire1880 ) | ( n_n907  &  wire6716  &  wire637 ) ;
 assign _9179 = ( (~ i_32_)  &  (~ i_34_)  &  i_33_  &  i_38_ ) ;
 assign _9188 = ( i_40_  &  (~ i_7_)  &  i_6_  &  i_39_ ) ;
 assign _9216 = ( wire36  &  i_18_ ) ;
 assign _9236 = ( wire1845 ) | ( wire1847 ) | ( wire6791  &  _9216 ) ;
 assign _9262 = ( i_25_  &  (~ i_32_)  &  i_33_ ) | ( i_26_  &  (~ i_32_)  &  i_33_ ) ;
 assign _9283 = ( (~ i_21_)  &  i_15_  &  n_n951 ) ;
 assign _9284 = ( (~ i_21_)  &  i_18_ ) ;
 assign _9291 = ( (~ i_12_)  &  i_11_  &  wire407 ) | ( i_12_  &  (~ i_11_)  &  wire407 ) ;
 assign _9302 = ( (~ i_12_)  &  i_16_  &  i_15_ ) ;
 assign _9303 = ( (~ i_12_)  &  i_17_  &  i_15_ ) ;
 assign _9305 = ( i_12_  &  i_17_  &  i_15_ ) ;
 assign _9306 = ( (~ i_39_)  &  i_16_  &  (~ i_38_)  &  i_37_ ) ;
 assign _9322 = ( (~ i_40_)  &  i_39_  &  (~ i_38_) ) ;
 assign _9369 = ( i_15_  &  i_12_ ) ;
 assign _9411 = ( i_11_  &  (~ i_17_)  &  i_15_ ) ;
 assign _9416 = ( i_12_  &  (~ i_17_)  &  i_15_ ) ;
 assign _9420 = ( (~ i_39_)  &  (~ i_38_)  &  i_37_ ) ;
 assign _9425 = ( i_40_  &  (~ i_39_)  &  (~ i_38_) ) ;
 assign _9430 = ( wire1780 ) | ( wire6853 ) | ( wire6854 ) ;
 assign _9433 = ( i_24_  &  i_22_  &  n_n793  &  wire607 ) ;
 assign _9445 = ( (~ i_39_)  &  i_40_ ) ;
 assign _9451 = ( (~ i_21_)  &  i_19_  &  n_n793 ) ;
 assign _9473 = ( wire1751 ) | ( n_n1986 ) ;
 assign _9479 = ( i_40_  &  (~ i_39_)  &  i_4_  &  i_38_ ) ;
 assign _9483 = ( i_4_  &  i_36_  &  (~ i_35_)  &  (~ i_37_) ) ;
 assign _9498 = ( wire1749 ) | ( wire1747 ) | ( _1063 ) | ( _1065 ) ;
 assign _9527 = ( (~ i_32_)  &  (~ i_34_)  &  i_33_ ) ;
 assign _9531 = ( wire6886 ) | ( wire6894 ) | ( _9473 ) | ( _9498 ) ;
 assign _9533 = ( i_4_  &  (~ i_7_) ) ;
 assign _9535 = ( i_1_  &  (~ i_7_) ) ;
 assign _9543 = ( i_3_  &  (~ i_7_) ) ;
 assign _9547 = ( i_3_  &  (~ i_7_) ) ;
 assign _9549 = ( i_1_  &  (~ i_7_) ) ;
 assign _9552 = ( wire80  &  n_n833  &  _9547 ) | ( wire80  &  n_n833  &  _9549 ) ;
 assign _9553 = ( wire80  &  n_n926  &  _9533 ) | ( wire80  &  n_n926  &  _9535 ) ;
 assign _9554 = ( n_n1993 ) | ( n_n2213 ) | ( wire1812 ) | ( _9553 ) ;
 assign _9555 = ( i_0_  &  (~ i_4_) ) ;
 assign _9558 = ( (~ i_32_)  &  (~ i_34_)  &  i_33_ ) ;
 assign _9580 = ( i_0_  &  (~ i_1_) ) ;
 assign _9598 = ( (~ i_40_)  &  (~ i_7_)  &  i_39_ ) ;
 assign _9615 = ( (~ i_39_)  &  i_40_ ) ;
 assign _9621 = ( (~ i_23_)  &  (~ i_32_)  &  (~ i_34_)  &  i_33_ ) ;
 assign _9636 = ( (~ i_40_)  &  i_39_  &  (~ i_23_) ) ;
 assign _9680 = ( i_39_  &  i_38_  &  (~ i_37_) ) ;
 assign _9690 = ( i_40_  &  (~ i_34_)  &  (~ i_36_)  &  i_35_ ) ;
 assign _9694 = ( (~ i_34_)  &  (~ i_36_)  &  (~ i_35_)  &  wire400 ) ;
 assign _9700 = ( i_39_  &  i_38_  &  (~ i_37_) ) ;
 assign _9705 = ( wire1653 ) | ( wire6981 ) | ( wire831  &  _9694 ) ;
 assign _9715 = ( n_n1581 ) | ( wire6987 ) | ( n_n1607 ) | ( _9705 ) ;
 assign _9718 = ( (~ i_32_)  &  i_33_  &  (~ i_38_)  &  (~ i_37_) ) ;
 assign _9721 = ( (~ i_32_)  &  i_33_  &  i_38_  &  i_37_ ) ;
 assign _9723 = ( (~ i_40_)  &  (~ i_39_)  &  (~ i_1_)  &  (~ i_38_) ) ;
 assign _9724 = ( (~ i_40_)  &  (~ i_39_)  &  (~ i_4_)  &  (~ i_38_) ) ;
 assign _9728 = ( wire80  &  n_n833  &  _9547 ) | ( wire80  &  n_n833  &  _9549 ) ;
 assign _9732 = ( n_n1990 ) | ( wire7002 ) | ( _970 ) ;
 assign _9735 = ( wire6994 ) | ( wire6998 ) | ( i_2_  &  wire835 ) ;
 assign _9737 = ( i_39_  &  i_40_ ) ;
 assign _9741 = ( i_39_  &  i_40_ ) ;
 assign _9747 = ( i_17_  &  i_16_  &  (~ i_32_)  &  (~ i_31_) ) ;
 assign _9752 = ( i_9_  &  (~ i_7_)  &  (~ i_5_)  &  n_n1066 ) ;
 assign _9755 = ( (~ i_12_)  &  n_n1009  &  wire82  &  _9741 ) ;
 assign _9756 = ( (~ i_12_)  &  n_n926  &  wire82 ) ;
 assign _9762 = ( (~ i_12_)  &  i_11_  &  wire7014 ) | ( i_12_  &  (~ i_11_)  &  wire7014 ) ;
 assign _9769 = ( wire1620 ) | ( wire7020 ) | ( wire319  &  _9755 ) ;
 assign _9770 = ( wire1626 ) | ( _959 ) | ( _960 ) | ( _9769 ) ;
 assign _9774 = ( (~ i_40_)  &  i_39_  &  (~ i_23_) ) ;
 assign _9785 = ( (~ i_34_)  &  (~ i_36_)  &  (~ i_35_)  &  wire400 ) ;
 assign _9794 = ( wire1653 ) | ( wire6981 ) | ( wire831  &  _9785 ) ;
 assign _9797 = ( n_n1628 ) | ( n_n1630 ) | ( n_n1631 ) ;
 assign _9801 = ( i_13_  &  (~ i_32_)  &  i_33_ ) ;
 assign _9806 = ( (~ i_7_)  &  (~ i_3_)  &  i_4_ ) ;
 assign _9811 = ( (~ i_40_)  &  i_9_  &  i_39_  &  i_38_ ) ;
 assign _9823 = ( (~ i_36_)  &  (~ i_35_)  &  (~ i_37_) ) ;
 assign _9825 = ( i_40_  &  i_9_  &  i_39_  &  i_38_ ) ;
 assign _9831 = ( i_9_  &  (~ i_14_)  &  i_16_ ) ;
 assign _9879 = ( i_33_  &  (~ i_32_) ) ;
 assign _9883 = ( i_33_  &  (~ i_32_) ) ;
 assign _9886 = ( i_11_  &  (~ i_32_)  &  i_33_ ) ;
 assign _9905 = ( (~ i_34_)  &  (~ i_7_) ) ;
 assign _9907 = ( (~ i_5_)  &  (~ i_7_) ) ;
 assign _9914 = ( i_32_  &  i_36_  &  (~ i_38_)  &  (~ i_37_) ) ;
 assign _9917 = ( i_34_  &  (~ i_6_) ) ;
 assign _9921 = ( wire7110 ) | ( wire1518 ) | ( _848 ) | ( _849 ) ;
 assign _9935 = ( (~ i_40_)  &  (~ i_39_)  &  (~ i_38_) ) ;
 assign _9966 = ( (~ i_34_)  &  i_33_  &  (~ i_35_) ) ;
 assign _9971 = ( i_17_  &  i_16_  &  (~ i_32_)  &  (~ i_31_) ) ;
 assign _9977 = ( wire7129 ) | ( wire1489 ) ;
 assign _9980 = ( (~ i_32_)  &  i_33_  &  i_38_  &  i_37_ ) ;
 assign _9982 = ( (~ i_32_)  &  i_33_  &  i_38_  &  (~ i_37_) ) ;
 assign _9983 = ( (~ i_15_)  &  (~ i_5_) ) ;
 assign _9987 = ( i_33_  &  (~ i_32_) ) ;
 assign _9989 = ( _790 ) | ( _789 ) ;
 assign _9990 = ( (~ i_40_)  &  (~ i_5_)  &  (~ i_39_)  &  (~ i_15_) ) ;
 assign _9999 = ( wire158 ) | ( n_n1009  &  wire422  &  _9990 ) ;
 assign _10009 = ( i_9_  &  (~ i_5_)  &  i_39_  &  i_38_ ) ;
 assign _10010 = ( wire1428 ) | ( wire140 ) ;
 assign _10011 = ( (~ i_37_)  &  i_35_ ) ;
 assign _10028 = ( wire7170 ) | ( _788 ) | ( _9989 ) | ( _9999 ) ;
 assign _10068 = ( wire156 ) | ( wire1416 ) | ( wire1459 ) | ( wire7153 ) ;
 assign _10069 = ( i_38_  &  (~ i_39_) ) ;
 assign _10072 = ( _745 ) | ( n_n966  &  n_n1073  &  _10069 ) ;
 assign _10073 = ( wire7190 ) | ( wire7139 ) | ( wire7140 ) | ( _9977 ) ;
 assign _10082 = ( (~ i_7_)  &  i_5_  &  (~ i_0_)  &  i_37_ ) ;
 assign _10085 = ( (~ i_7_)  &  (~ i_31_)  &  i_33_ ) ;
 assign _10089 = ( (~ i_7_)  &  (~ i_31_)  &  i_33_ ) ;
 assign _10093 = ( n_n1047  &  wire7201  &  _10089 ) | ( n_n1047  &  wire7200  &  _10089 ) ;
 assign _10114 = ( (~ i_7_)  &  i_5_  &  i_33_ ) ;
 assign _10120 = ( (~ i_14_)  &  (~ i_34_)  &  i_33_  &  (~ i_35_) ) ;
 assign _10125 = ( (~ i_7_)  &  (~ i_31_)  &  i_33_ ) ;
 assign _10131 = ( (~ i_7_)  &  i_5_  &  (~ i_0_)  &  i_38_ ) ;
 assign _10136 = ( wire7211 ) | ( _725 ) | ( wire354  &  wire7208 ) ;
 assign _10141 = ( i_0_  &  (~ i_32_)  &  i_33_ ) ;
 assign _10142 = ( i_39_  &  (~ i_32_)  &  (~ i_34_)  &  i_33_ ) ;
 assign _10143 = ( (~ i_32_)  &  (~ i_34_)  &  i_33_  &  (~ i_38_) ) ;
 assign _10151 = ( n_n970  &  _10142 ) | ( wire6731  &  _10143 ) ;
 assign _10152 = ( _10151 ) | ( i_38_  &  wire1362 ) | ( i_38_  &  wire7234 ) ;
 assign _10173 = ( (~ i_32_)  &  (~ i_34_)  &  i_33_ ) ;
 assign _10177 = ( (~ i_34_)  &  (~ i_36_)  &  i_35_ ) ;
 assign _10178 = ( (~ i_32_)  &  (~ i_34_)  &  i_33_  &  (~ i_38_) ) ;
 assign _10179 = ( (~ i_39_)  &  (~ i_32_)  &  (~ i_34_)  &  i_33_ ) ;
 assign _10180 = ( i_40_  &  (~ i_32_)  &  (~ i_34_)  &  i_33_ ) ;
 assign _10181 = ( (~ i_32_)  &  i_34_  &  i_33_  &  i_38_ ) ;
 assign _10182 = ( wire7227  &  _10177 ) | ( n_n864  &  _10178 ) ;
 assign _10186 = ( (~ i_11_)  &  (~ i_36_)  &  (~ i_35_)  &  (~ i_37_) ) ;
 assign _10187 = ( (~ i_12_)  &  (~ i_36_)  &  (~ i_35_)  &  (~ i_37_) ) ;
 assign _10194 = ( wire806  &  wire805 ) | ( wire748  &  _10173 ) ;
 assign _10207 = ( (~ i_32_)  &  i_33_  &  (~ i_38_)  &  i_37_ ) ;
 assign _10212 = ( (~ i_39_)  &  (~ i_32_)  &  i_34_  &  i_33_ ) ;
 assign _10213 = ( (~ i_40_)  &  (~ i_32_)  &  i_34_  &  i_33_ ) ;
 assign _10233 = ( i_40_  &  i_39_  &  i_38_ ) ;
 assign _10277 = ( (~ i_7_)  &  (~ i_32_)  &  i_33_  &  i_38_ ) ;
 assign _10285 = ( i_38_  &  i_39_ ) ;
 assign _10296 = ( i_33_  &  (~ i_31_) ) ;
 assign _10305 = ( i_15_  &  i_24_ ) ;
 assign _10311 = ( (~ i_36_)  &  (~ i_38_)  &  (~ i_37_) ) ;
 assign _10330 = ( _618 ) | ( _619 ) | ( wire723  &  _10311 ) ;
 assign _10339 = ( (~ i_40_)  &  i_38_  &  i_37_ ) ;
 assign _10358 = ( (~ i_7_)  &  i_32_  &  i_33_ ) ;
 assign _10361 = ( wire1246 ) | ( wire1247 ) | ( wire7341 ) | ( _593 ) ;
 assign _10362 = ( wire7301 ) | ( wire1295 ) | ( wire7293 ) | ( _10330 ) ;
 assign _10388 = ( n_n1986 ) | ( wire1747 ) | ( wire1222 ) | ( _1063 ) ;
 assign _10392 = ( wire80  &  n_n833  &  _9547 ) | ( wire80  &  n_n833  &  _9549 ) ;
 assign _10403 = ( wire245 ) | ( wire176 ) | ( wire7378 ) ;
 assign _10409 = ( wire185 ) | ( n_n1607 ) | ( _9705 ) | ( _10403 ) ;
 assign _10411 = ( n_n2581 ) | ( wire80  &  n_n926  &  _9533 ) ;
 assign _10421 = ( (~ i_22_)  &  (~ i_32_)  &  i_33_ ) ;
 assign _10434 = ( i_39_  &  i_40_ ) ;
 assign _10435 = ( i_2_  &  i_0_  &  (~ i_32_)  &  n_n1066 ) ;
 assign _10436 = ( i_3_  &  i_0_  &  (~ i_32_) ) ;
 assign _10437 = ( i_1_  &  i_0_  &  (~ i_32_) ) ;
 assign _10483 = ( i_15_  &  (~ i_16_) ) ;
 assign _10507 = ( (~ i_22_)  &  (~ i_32_)  &  i_33_ ) ;
 assign _10519 = ( _512 ) | ( _513 ) | ( wire113  &  wire7428 ) ;
 assign _10525 = ( (~ i_1_)  &  i_0_  &  (~ i_32_) ) ;
 assign _10530 = ( (~ i_39_)  &  i_40_ ) ;
 assign _10535 = ( i_3_  &  (~ i_32_)  &  i_33_ ) | ( i_1_  &  (~ i_32_)  &  i_33_ ) ;
 assign _10542 = ( i_4_  &  (~ i_32_)  &  i_33_ ) ;
 assign _10545 = ( wire1155 ) | ( wire1158 ) | ( wire7446 ) ;
 assign _10546 = ( wire7444 ) | ( wire7445 ) | ( wire7440 ) | ( _10545 ) ;
 assign _10547 = ( n_n1414 ) | ( n_n1412 ) | ( wire7412 ) | ( _10546 ) ;
 assign _10549 = ( i_24_  &  (~ i_22_)  &  n_n1074  &  wire87 ) ;
 assign _10552 = ( i_24_  &  (~ i_32_)  &  (~ i_34_)  &  i_33_ ) ;
 assign _10554 = ( i_24_  &  (~ i_32_)  &  (~ i_34_)  &  i_33_ ) ;
 assign _10561 = ( i_38_  &  i_39_ ) ;
 assign _10584 = ( i_40_  &  (~ i_7_)  &  (~ i_32_) ) ;
 assign _10586 = ( _452 ) | ( n_n1066  &  n_n668  &  wire713 ) ;
 assign _10588 = ( (~ i_7_)  &  (~ i_34_)  &  (~ i_36_)  &  (~ i_35_) ) ;
 assign _10607 = ( (~ i_7_)  &  i_5_  &  (~ i_39_)  &  (~ i_0_) ) ;
 assign _10613 = ( (~ i_7_)  &  (~ i_34_)  &  (~ i_36_)  &  (~ i_35_) ) ;
 assign _10615 = ( (~ i_11_)  &  i_9_ ) ;
 assign _10617 = ( (~ i_11_)  &  i_9_ ) ;
 assign _10634 = ( wire1088 ) | ( wire1092 ) ;
 assign _10636 = ( (~ i_40_)  &  i_9_  &  i_39_  &  i_38_ ) ;
 assign _10643 = ( (~ i_7_)  &  (~ i_34_)  &  (~ i_36_)  &  (~ i_35_) ) ;
 assign _10651 = ( (~ i_40_)  &  (~ i_7_)  &  (~ i_39_) ) ;
 assign _10653 = ( (~ i_40_)  &  (~ i_7_)  &  (~ i_39_) ) ;
 assign _10657 = ( (~ i_32_)  &  (~ i_34_)  &  i_33_ ) ;
 assign _10668 = ( (~ i_7_)  &  i_5_  &  (~ i_0_)  &  i_38_ ) ;
 assign _10677 = ( i_23_  &  i_24_  &  i_22_  &  i_15_ ) ;
 assign _10678 = ( _10677  &  wire35 ) ;
 assign _10691 = ( i_24_  &  wire731  &  wire7511 ) ;
 assign _10693 = ( i_24_  &  (~ i_32_)  &  (~ i_34_)  &  i_33_ ) ;
 assign _10696 = ( (~ i_7_)  &  (~ i_5_)  &  i_12_ ) ;
 assign _10699 = ( i_20_  &  i_21_  &  i_22_  &  i_15_ ) ;
 assign _10704 = ( (~ i_7_)  &  (~ i_5_)  &  i_11_ ) ;
 assign _10705 = ( wire1044 ) | ( wire7518 ) | ( i_25_  &  wire575 ) ;
 assign _10712 = ( i_12_  &  i_17_  &  i_15_ ) ;
 assign _10718 = ( (~ i_21_)  &  i_15_  &  n_n951 ) ;
 assign _10723 = ( (~ i_30_)  &  (~ i_32_)  &  (~ i_31_)  &  n_n1066 ) ;
 assign _10724 = ( wire156 ) | ( wire6907  &  n_n935  &  _9425 ) ;
 assign _10772 = ( (~ i_23_)  &  (~ i_21_)  &  i_15_ ) ;
 assign _10803 = ( i_39_  &  (~ i_40_) ) ;
 assign _10804 = ( i_10_  &  i_27_  &  (~ i_39_)  &  i_38_ ) ;
 assign _10809 = ( wire925 ) | ( wire926 ) | ( wire928 ) | ( wire929 ) ;
 assign _10810 = ( (~ i_31_)  &  (~ i_32_) ) ;
 assign _10818 = ( (~ i_23_)  &  (~ i_21_)  &  i_15_ ) ;
 assign _10830 = ( (~ i_36_)  &  (~ i_35_)  &  (~ i_37_) ) ;
 assign _10837 = ( (~ i_18_)  &  (~ i_34_)  &  (~ i_36_)  &  i_35_ ) ;
 assign _10867 = ( i_40_  &  (~ i_7_)  &  (~ i_32_)  &  i_33_ ) ;
 assign _10875 = ( (~ i_7_)  &  i_25_ ) | ( (~ i_7_)  &  (~ i_26_) ) ;
 assign _10886 = ( (~ i_7_)  &  (~ i_36_)  &  i_37_ ) ;
 assign _10890 = ( wire7555 ) | ( wire50  &  n_n693  &  _10875 ) ;
 assign _10896 = ( i_0_  &  (~ i_1_) ) ;
 assign _10897 = ( wire79  &  wire7630  &  _9555 ) | ( wire79  &  wire7630  &  _10896 ) ;
 assign _10899 = ( (~ i_7_)  &  i_1_  &  i_0_ ) ;
 assign _10903 = ( wire131 ) | ( wire893 ) | ( _250 ) | ( _10897 ) ;
 assign _10904 = ( n_n1957 ) | ( wire904 ) | ( wire905 ) | ( wire7625 ) ;
 assign _10925 = ( i_11_  &  i_18_  &  i_15_ ) | ( i_11_  &  i_15_  &  i_19_ ) ;
 assign _10927 = ( i_9_  &  (~ i_7_)  &  (~ i_5_) ) ;
 assign _10931 = ( (~ i_34_)  &  i_33_  &  (~ i_35_)  &  i_29_ ) ;
 assign _10933 = ( i_30_  &  (~ i_31_)  &  (~ i_29_) ) ;
 assign _10935 = ( (~ i_40_)  &  i_39_  &  (~ i_38_)  &  i_37_ ) ;
 assign _10941 = ( i_40_  &  (~ i_39_)  &  (~ i_31_) ) ;
 assign _10943 = ( i_40_  &  i_39_  &  (~ i_13_) ) ;
 assign _10946 = ( (~ i_36_)  &  (~ i_38_)  &  i_37_ ) ;
 assign _10973 = ( wire849 ) | ( _221 ) | ( (~ i_40_)  &  wire843 ) ;
 assign _10982 = ( (~ i_39_)  &  i_40_ ) ;
 assign _10987 = ( (~ i_10_)  &  (~ i_7_) ) | ( (~ i_7_)  &  (~ i_27_) ) ;
 assign _10989 = ( (~ i_39_)  &  (~ i_40_) ) ;
 assign _10991 = ( wire227 ) | ( wire869 ) | ( wire872 ) | ( _193 ) ;
 assign _11002 = ( i_40_  &  (~ i_38_)  &  i_37_ ) ;
 assign _11007 = ( wire7654 ) | ( wire7658 ) | ( wire7659 ) | ( _10991 ) ;
 assign _11009 = ( n_n1330 ) | ( n_n1332 ) | ( wire7681 ) | ( _11007 ) ;
 assign _11018 = ( i_15_  &  (~ i_16_) ) ;
 assign _11020 = ( i_15_  &  (~ i_16_) ) ;
 assign _11022 = ( (~ i_11_)  &  (~ i_9_) ) ;
 assign _11043 = ( wire286 ) | ( wire288 ) | ( wire289 ) ;
 assign _11046 = ( i_9_  &  i_17_  &  i_15_ ) | ( i_9_  &  i_16_  &  i_15_ ) ;
 assign _11057 = ( wire279 ) | ( n_n1068  &  wire520 ) ;
 assign _11058 = ( wire287 ) | ( wire7728 ) | ( _11043 ) | ( _11057 ) ;
 assign _11060 = ( (~ i_15_)  &  (~ i_32_)  &  (~ i_34_)  &  i_33_ ) ;
 assign _11064 = ( (~ i_14_)  &  (~ i_32_)  &  (~ i_34_)  &  i_33_ ) ;
 assign _11066 = ( i_3_  &  (~ i_32_)  &  i_33_ ) | ( i_4_  &  (~ i_32_)  &  i_33_ ) ;
 assign _11073 = ( i_39_  &  (~ i_32_)  &  (~ i_34_)  &  i_33_ ) ;
 assign _11074 = ( (~ i_12_)  &  (~ i_32_)  &  (~ i_34_)  &  i_33_ ) ;
 assign _11076 = ( n_n970  &  _11073 ) | ( wire6739  &  _11074 ) ;
 assign _11079 = ( i_0_  &  i_1_ ) ;
 assign _11080 = ( i_0_  &  i_4_ ) ;
 assign _11089 = ( i_2_  &  (~ i_32_)  &  i_33_ ) ;
 assign _11092 = ( (~ i_5_)  &  i_28_ ) | ( (~ i_5_)  &  i_29_ ) ;
 assign _11094 = ( i_4_  &  i_0_  &  (~ i_32_) ) ;
 assign _11095 = ( i_2_  &  i_0_  &  (~ i_32_) ) ;
 assign _11099 = ( _129 ) | ( _130 ) | ( _131 ) | ( _132 ) ;
 assign _11107 = ( (~ i_38_)  &  (~ i_39_) ) ;
 assign _11109 = ( (~ i_38_)  &  (~ i_39_) ) ;
 assign _11112 = ( i_39_  &  (~ i_12_)  &  i_11_  &  i_38_ ) | ( i_39_  &  i_12_  &  (~ i_11_)  &  i_38_ ) ;
 assign _11116 = ( wire451 ) | ( wire454 ) | ( _122 ) | ( _123 ) ;
 assign _11119 = ( (~ i_22_)  &  (~ i_32_)  &  i_33_ ) ;
 assign _11124 = ( _113 ) | ( _114 ) | ( _115 ) | ( _116 ) ;
 assign _11128 = ( i_39_  &  i_40_ ) ;
 assign _11145 = ( (~ i_39_)  &  i_40_ ) ;
 assign _11153 = ( (~ i_25_)  &  (~ i_32_)  &  i_33_ ) ;
 assign _11155 = ( i_1_  &  (~ i_32_)  &  i_33_ ) ;
 assign _11161 = ( wire7692 ) | ( wire446 ) | ( _11116 ) | ( _11124 ) ;
 assign _11170 = ( (~ i_7_)  &  (~ i_39_)  &  i_25_ ) ;
 assign _11184 = ( i_13_  &  (~ i_36_)  &  (~ i_38_)  &  i_37_ ) ;
 assign _11201 = ( (~ i_7_)  &  (~ i_5_)  &  i_24_ ) ;
 assign _11220 = ( wire191 ) | ( wire192 ) | ( _78 ) | ( _79 ) ;
 assign _11232 = ( n_n785  &  wire463 ) | ( n_n785  &  wire840  &  wire7817 ) ;
 assign _11234 = ( (~ i_21_)  &  i_15_  &  wire469  &  n_n428 ) ;
 assign _11241 = ( n_n945  &  wire6789  &  n_n860 ) ;
 assign _11244 = ( i_18_  &  (~ i_21_)  &  i_15_  &  i_19_ ) ;
 assign _11249 = ( i_11_  &  i_18_  &  i_15_ ) ;
 assign _11256 = ( (~ i_7_)  &  (~ i_39_)  &  (~ i_26_) ) ;
 assign _11261 = ( (~ i_40_)  &  i_34_  &  (~ i_36_)  &  (~ i_35_) ) ;
 assign _11278 = ( (~ i_17_)  &  (~ i_16_)  &  i_31_  &  (~ i_36_) ) ;


endmodule

