module spla_mapped (
	i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_14_, i_3_, 
	i_13_, i_4_, i_12_, i_1_, i_11_, i_2_, i_0_, i_15_, o_1_, o_19_, 
	o_2_, o_0_, o_29_, o_39_, o_38_, o_25_, o_12_, o_37_, o_26_, o_11_, 
	o_36_, o_27_, o_14_, o_35_, o_28_, o_13_, o_34_, o_21_, o_16_, o_40_, 
	o_33_, o_22_, o_15_, o_32_, o_23_, o_18_, o_31_, o_24_, o_17_, o_43_, 
	o_30_, o_44_, o_41_, o_42_, o_20_, o_45_, o_10_, o_9_, o_7_, o_8_, 
	o_5_, o_6_, o_3_, o_4_);

input i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_14_, i_3_, i_13_, i_4_, i_12_, i_1_, i_11_, i_2_, i_0_, i_15_;

output o_1_, o_19_, o_2_, o_0_, o_29_, o_39_, o_38_, o_25_, o_12_, o_37_, o_26_, o_11_, o_36_, o_27_, o_14_, o_35_, o_28_, o_13_, o_34_, o_21_, o_16_, o_40_, o_33_, o_22_, o_15_, o_32_, o_23_, o_18_, o_31_, o_24_, o_17_, o_43_, o_30_, o_44_, o_41_, o_42_, o_20_, o_45_, o_10_, o_9_, o_7_, o_8_, o_5_, o_6_, o_3_, o_4_;

wire wire5057, wire16872, n_n5144, wire736, wire16876, n_n162, wire16877, wire16898, wire5026, wire5027, wire16911, n_n4721, wire16933, n_n4399, n_n17, n_n159, n_n4103, n_n4102, wire17601, wire17602, n_n4, wire17604, wire17612, wire17849, wire17861, wire17862, wire17876, wire17877, wire17913, wire17915, wire18141, wire18142, wire18148, n_n2998, wire18154, wire18155, wire18167, wire18212, wire18213, wire18214, wire18292, wire18297, n_n10, wire185, wire270, wire18299, n_n2721, wire3442, wire18310, wire18311, n_n135, wire267, wire3439, n_n259, wire18323, wire18329, wire18330, n_n14, wire18354, wire18355, n_n3166, wire18437, wire18490, wire18499, wire18512, wire18526, wire18565, wire3194, wire18568, wire18572, n_n16, n_n2748, wire18621, wire18623, wire18682, wire18683, wire18685, n_n4845, wire18795, wire2962, wire18802, wire18803, wire18807, wire18809, wire19030, wire19349, wire19459, wire19869, wire19914, n_n5, wire19922, wire19928, n_n275, wire441, wire19941, wire19946, n_n219, n_n218, wire428, n_n184, n_n163, wire725, n_n35, wire729, n_n65, n_n71, n_n124, n_n9, wire343, n_n48, n_n220, n_n38, wire244, wire5024, n_n373, wire140, n_n39, wire5022, n_n374, n_n134, n_n132, n_n969, wire1595, n_n54, n_n52, n_n519, n_n4597, n_n156, n_n205, n_n211, wire390, n_n177, wire719, wire393, wire712, wire714, n_n31, n_n30, wire143, wire154, wire47, n_n4161, n_n170, wire720, wire722, wire715, wire132, wire723, wire730, wire727, wire137, n_n4449, wire1864, wire17164, wire599, wire146, wire131, wire695, wire17198, wire17213, n_n2239, wire4643, wire17249, wire17256, wire17257, wire4561, wire4562, wire17303, wire17305, wire17322, n_n2249, wire17341, wire17342, n_n2265, n_n2266, wire17379, n_n2234, n_n4120, wire4434, wire17420, n_n4106, n_n19, n_n111, n_n7241, n_n7240, n_n51, wire747, n_n13, wire717, n_n149, wire77, wire431, wire529, wire568, wire569, n_n53, n_n3825, wire4060, wire17726, wire17729, n_n3795, n_n3800, n_n3802, wire17798, n_n3787, wire17831, wire17832, wire17836, wire17839, wire721, wire728, wire157, n_n157, wire213, n_n36, n_n34, wire597, wire620, n_n2630, wire17884, n_n2622, n_n3467, wire17934, wire17935, n_n3454, n_n3473, wire17958, wire17959, wire17968, n_n3456, n_n7263, n_n161, n_n7265, n_n7267, wire3628, wire3629, wire18150, wire253, n_n4308, n_n6271, n_n126, n_n6267, n_n47, wire152, wire4260, wire17554, n_n3085, n_n6266, n_n6270, n_n6269, n_n6268, wire245, n_n5052, n_n41, n_n40, n_n57, wire144, n_n5055, wire122, wire3469, wire751, wire18298, wire525, n_n200, n_n33, wire1417, wire55, wire149, wire127, n_n2728, wire675, wire3451, wire18301, wire18302, wire126, wire587, wire172, wire147, wire158, wire133, wire767, n_n6, n_n3389, n_n191, wire145, wire388, wire770, n_n3179, wire18375, n_n144, n_n7346, n_n3, n_n2, wire430, wire708, n_n18, n_n5319, wire17587, wire684, n_n197, n_n212, n_n4441, wire575, wire18577, wire18578, n_n2754, wire18593, wire18594, n_n2747, n_n101, n_n42, wire3128, wire18624, wire18625, wire18626, n_n4755, wire381, n_n43, wire63, wire48, wire662, wire18711, wire18712, wire18719, wire2977, wire18783, wire18789, wire18790, n_n6005, wire17072, wire419, wire445, wire446, wire3470, wire18360, wire18361, wire95, n_n799, wire2310, wire19504, wire777, wire776, wire775, n_n7252, wire389, wire3248, wire454, wire742, wire779, wire783, wire781, wire707, n_n46, n_n199, wire726, wire724, wire168, n_n138, n_n216, wire214, n_n5107, n_n108, n_n148, wire90, n_n5000, wire98, n_n102, n_n1434, wire118, n_n1408, wire120, wire179, wire324, wire18720, wire789, n_n117, n_n1426, n_n89, wire93, wire241, wire273, wire791, wire53, n_n77, n_n1416, wire117, wire281, wire294, wire793, n_n125, wire85, wire142, wire422, wire150, wire80, wire78, n_n55, wire252, wire796, wire207, n_n150, n_n1520, wire155, wire205, wire215, wire17490, wire800, wire234, wire86, wire84, wire799, wire181, wire134, wire156, wire458, wire176, wire123, wire541, wire4393, n_n3912, n_n123, wire570, wire60, n_n1700, wire220, wire803, wire17470, wire17471, wire4829, n_n214, wire4354, wire4355, n_n1624, wire17479, wire17486, n_n4112, n_n155, n_n1594, wire17082, wire808, wire180, n_n4904, wire447, wire4320, n_n5037, n_n5033, wire219, wire108, n_n4903, wire1844, wire4935, wire544, wire17501, wire716, wire718, wire52, wire129, n_n4622, wire182, n_n5060, n_n130, n_n3276, n_n83, n_n6445, n_n7242, n_n68, wire344, wire462, wire817, wire130, wire188, n_n59, wire226, wire820, wire4558, wire17307, wire4554, wire17314, wire304, wire306, wire824, wire4701, wire17178, n_n2253, n_n61, wire228, n_n147, n_n63, wire351, wire377, wire139, n_n213, wire257, wire313, n_n129, n_n166, n_n127, n_n82, wire190, wire334, wire836, n_n139, wire260, wire373, wire2900, wire18865, wire18866, n_n1870, n_n95, wire74, wire136, wire840, wire18857, wire18874, n_n1800, wire68, n_n112, n_n113, wire227, wire232, wire844, wire845, wire542, wire850, wire849, n_n5109, wire677, wire75, wire19119, wire852, n_n140, n_n142, wire290, wire856, n_n116, wire255, wire199, wire402, wire19640, wire19641, wire859, wire743, n_n103, n_n207, n_n173, n_n169, n_n204, n_n151, n_n141, n_n115, n_n209, n_n178, n_n183, n_n90, n_n70, n_n62, n_n189, n_n122, n_n185, n_n84, n_n136, n_n210, n_n172, n_n58, n_n118, n_n32, n_n186, n_n107, n_n198, n_n168, n_n176, n_n60, n_n12, wire151, wire94, wire184, wire268, wire18738, wire860, wire81, n_n1442, wire111, wire162, wire164, wire341, wire863, wire206, wire243, wire368, wire18752, wire865, wire153, n_n4686, wire247, wire135, wire704, n_n4231, wire218, wire248, n_n4460, n_n4900, wire867, n_n4518, wire1224, wire17100, wire532, wire4739, wire4740, wire17102, wire594, wire660, wire17521, wire17522, n_n4116, wire104, n_n5111, n_n5113, wire868, n_n7254, n_n7248, n_n3562, wire3601, wire18168, wire18169, n_n3398, wire481, wire3594, wire18172, wire18173, wire18174, n_n3050, wire124, wire128, wire875, wire18180, n_n3033, wire711, wire87, wire877, n_n2948, wire16880, n_n231, wire308, wire887, wire189, wire299, wire896, wire894, wire561, wire4658, wire4659, wire17217, wire899, wire200, wire201, wire902, wire376, n_n201, wire904, wire2861, wire18892, n_n1862, wire911, wire18901, n_n1799, wire246, wire254, wire913, n_n2881, wire69, n_n1708, wire223, wire239, wire916, wire51, n_n1717, wire564, wire924, wire2610, wire19138, n_n1170, wire70, wire233, wire251, wire925, wire928, n_n4674, n_n78, n_n974, n_n215, wire933, n_n7260, n_n7266, wire19929, wire19933, wire551, n_n202, n_n72, n_n131, n_n182, n_n143, n_n137, n_n128, n_n190, n_n196, n_n64, n_n175, n_n171, n_n7264, n_n74, wire566, wire670, n_n4808, wire683, wire524, wire672, n_n4564, wire709, n_n4169, wire942, wire359, n_n1514, wire432, wire17034, wire17035, n_n4996, n_n4994, wire511, wire946, wire449, wire656, wire17410, wire443, n_n4240, wire4965, wire4966, n_n4154, wire654, wire739, wire279, n_n4602, wire605, wire59, n_n5075, wire54, wire498, wire951, n_n6492, n_n3413, wire546, wire674, n_n3889, wire671, wire463, wire960, wire959, wire1730, wire18555, wire4485, wire4486, wire17367, wire17368, wire968, wire115, wire116, wire371, wire17253, wire971, n_n5739, wire17258, wire17259, wire17260, n_n2340, n_n5743, wire440, wire973, wire4619, wire17268, wire366, wire17272, wire975, wire979, wire978, wire362, n_n2310, wire17333, wire397, wire229, wire265, wire989, wire988, wire302, wire303, wire316, wire18831, wire993, wire18832, wire685, n_n5011, wire110, n_n1517, wire457, wire572, wire1003, wire1006, n_n832, wire1012, wire291, wire297, wire19621, wire1017, n_n56, n_n133, wire198, wire18773, wire1021, wire186, wire217, wire18780, wire1023, wire256, wire216, wire1022, wire224, n_n4981, wire208, wire225, wire148, wire17083, wire1030, n_n4620, wire1173, wire17528, n_n4131, wire17534, n_n4109, wire249, wire571, wire17033, wire549, n_n4476, wire537, wire4842, wire17007, wire621, wire17553, n_n3417, n_n6384, n_n3419, wire1036, n_n3421, wire391, wire1041, wire1044, wire1049, wire4481, wire17374, wire526, wire4531, wire17329, wire374, wire1056, wire4505, wire4506, wire4508, wire4509, n_n2257, wire1060, wire263, wire17361, wire1064, wire250, wire1069, wire62, n_n5019, wire19179, wire1070, wire65, wire1902, wire16987, wire760, wire1072, wire385, wire19196, wire19197, wire1075, wire277, wire1077, wire276, wire211, wire271, wire1079, n_n972, wire1084, wire1089, wire1087, wire1090, wire3433, wire3434, wire18316, n_n164, n_n5103, wire212, n_n5067, wire221, wire298, wire1096, wire591, wire515, wire4948, wire657, wire1789, wire17013, n_n4424, wire518, wire57, wire653, wire694, wire17018, wire17019, n_n4404, wire666, wire17050, wire17064, n_n4312, wire141, wire258, wire125, n_n4566, wire46, n_n1553, wire209, n_n5059, n_n5058, wire577, wire1115, wire1114, wire1116, wire1117, wire1120, wire358, wire17395, wire1124, wire1126, wire292, wire311, wire317, wire319, wire1129, wire321, wire326, wire327, wire1132, wire197, wire203, wire309, wire323, wire1135, wire1136, wire83, wire384, wire1143, wire330, wire1145, wire19221, wire1147, wire1150, wire1152, wire500, wire1154, wire1153, n_n3415, wire1160, wire1159, n_n7262, n_n73, n_n1606, wire100, wire1170, n_n3979, wire361, wire363, wire426, wire442, wire1174, wire1177, wire1176, wire1179, wire1178, wire655, wire1190, wire1189, wire1188, wire380, wire18986, wire1194, wire364, wire1197, wire1196, wire1195, wire18834, wire1401, wire331, n_n1826, wire1200, wire1199, wire18961, wire18962, wire18966, n_n1803, wire18981, wire312, wire1201, wire261, wire264, wire375, wire19001, wire1205, wire1207, wire92, wire19413, wire19414, wire1211, n_n1542, n_n4641, wire693, wire169, wire19320, wire1214, wire274, wire1216, wire1218, wire2083, n_n369, wire335, wire652, wire1229, wire18706, n_n3054, n_n2770, wire1234, wire412, wire1239, wire18938, wire18939, n_n3638, wire1242, wire1244, wire1243, wire1246, n_n1811, wire1247, wire1251, wire1255, wire1257, wire4869, n_n817, wire167, wire2329, wire2331, wire19480, wire19481, wire320, wire19660, wire1259, wire195, wire19663, wire1261, wire1260, wire1263, wire686, wire1271, n_n4692, wire1277, wire175, wire383, wire1279, wire1285, wire1287, wire1286, wire473, wire19253, wire1290, wire19250, wire1289, wire19260, wire1292, wire557, wire1294, wire1293, n_n1566, wire88, wire1295, n_n1575, wire349, wire1297, wire19464, wire1302, wire19469, wire1305, wire329, wire1311, wire171, n_n2859, n_n4657, wire160, wire174, wire651, n_n3570, n_n3573, wire1319, wire4182, n_n3823, wire222, wire1321, wire1326, n_n5070, wire3496, wire3497, wire18272, wire18273, n_n3037, wire469, wire1331, wire673, wire18283, n_n3029, wire1336, wire173, n_n2733, wire1341, wire378, wire1345, wire1343, wire1342, wire165, wire1347, wire280, wire1346, wire2302, wire2303, wire19510, n_n784, wire629, wire2308, wire19506, wire19516, n_n752, wire166, wire269, wire275, wire278, wire1354, wire1357, wire282, wire283, wire1363, wire296, wire262, wire332, wire342, wire1366, wire1367, wire479, n_n3525, wire1375, n_n3561, n_n3578, wire4067, wire17716, wire17717, wire1378, wire18454, wire18455, n_n3180, wire1381, wire1383, wire18461, n_n3170, wire1386, wire1390, wire1389, wire170, wire18534, wire1395, wire1404, wire1405, wire2080, n_n371, wire1416, wire1415, wire1414, wire759, wire645, wire664, wire394, wire240, wire187, wire210, wire17741, wire1420, n_n3592, wire648, wire681, wire17766, wire17767, n_n3834, n_n3601, wire504, n_n3833, wire1425, wire1427, wire1432, wire19099, wire1436, wire1437, wire19599, wire19600, n_n772, wire235, wire236, wire1444, wire325, n_n326, wire19701, wire1446, wire497, wire1450, wire636, wire18253, wire1459, wire1463, wire4223, wire17588, n_n2956, wire1465, wire1470, wire1469, wire401, wire1477, wire1476, wire1480, wire1479, wire1478, wire336, wire19895, wire1483, wire161, wire1482, wire16886, n_n5021, wire565, wire1488, wire579, wire1489, wire3985, wire17787, n_n3514, wire1491, wire17793, n_n3511, wire690, wire1493, wire1496, wire230, wire1498, wire347, wire352, wire1497, wire1500, wire1499, wire1503, wire1504, wire357, wire19328, wire1507, wire314, wire1510, wire259, wire337, wire19831, wire1513, wire338, wire1512, wire689, wire1519, wire1520, wire370, wire18367, n_n3176, wire1524, wire1527, wire315, wire1537, wire19442, wire19443, wire1539, n_n1163, wire348, wire1544, wire1553, wire1556, wire1558, wire1560, wire1562, wire295, wire333, wire19882, wire1568, wire1570, wire560, wire688, wire289, wire18426, wire1576, n_n3555, wire1580, wire1579, wire1578, wire19318, wire1581, wire1582, wire19835, wire1587, wire19901, wire1590, wire19905, wire1592, wire121, wire434, wire538, wire539, wire17918, wire17919, wire17920, wire17921, wire1601, n_n2777, wire1602, wire607, wire640, wire584, wire107, wire339, wire19523, wire1605, wire19767, wire1613, wire99, wire1617, wire18028, n_n3485, wire698, wire3820, wire17926, n_n3510, wire1625, wire578, wire3177, wire18581, wire18582, wire18583, wire1627, wire17880, wire17881, wire642, wire322, wire1628, wire407, wire1630, wire163, wire194, wire1632, n_n765, wire635, wire1633, wire19556, wire19557, wire19560, wire346, wire19796, wire1636, wire1640, wire1639, wire19786, wire19787, wire19793, n_n302, wire354, wire1641, wire19799, wire19812, wire17960, wire242, wire272, wire17944, wire1648, wire17947, wire17948, n_n3470, n_n2642, wire18611, wire1655, wire1658, wire2232, wire19569, wire1659, wire19574, wire1668, wire1666, wire19846, wire18122, n_n3501, wire18125, n_n3500, wire19577, wire1674, wire2218, wire19584, n_n834, wire1675, wire19587, wire19588, wire19591, wire19582, wire19596, wire415, wire1684, wire1689, wire696, n_n3542, wire3767, wire17979, wire17980, n_n3482, wire18032, n_n3487, wire18039, n_n3460, wire1695, wire1704, wire19624, wire1706, wire1709, wire1708, wire1707, wire2182, wire19614, wire19617, wire19619, wire1717, wire1716, wire1720, wire18657, wire1723, wire606, wire1729, wire17896, wire17897, wire17898, n_n2626, wire19013, wire1735, wire1739, wire1738, wire1741, wire237, wire1740, wire19633, wire1743, wire1742, wire1949, wire1748, wire1747, wire18044, n_n3492, wire18049, wire18050, wire18051, n_n3491, wire1751, wire18057, wire18058, n_n3462, wire18063, wire18064, n_n3489, wire18078, n_n3451, wire1754, wire1753, wire19630, wire1756, wire19654, wire1758, wire19856, wire1761, wire18978, wire1766, wire19672, wire1775, wire1779, wire1778, wire1777, wire1780, wire3403, wire18342, wire18345, wire1782, wire1786, wire19021, wire19023, n_n1801, wire4974, wire16952, wire16953, wire16954, n_n4419, wire202, wire307, wire17339, wire1794, wire17149, wire18004, wire1807, wire19500, wire1809, wire18007, wire1811, wire18014, wire1812, wire17903, wire1814, wire49, wire50, wire56, wire72, wire79, wire82, wire438, wire399, wire340, wire284, wire177, wire183, wire425, wire192, wire193, wire424, wire196, wire204, wire293, wire300, wire301, wire305, wire310, wire318, wire328, wire345, wire369, wire372, wire398, wire400, wire405, wire406, wire408, wire409, wire410, wire414, wire416, wire418, wire1840, wire16980, wire1853, wire1862, wire815, wire1128, wire1209, wire1253, wire1409, wire1550, wire1557, wire138, wire439, wire467, wire499, wire19899, wire507, wire510, wire513, wire520, wire552, wire19888, wire556, wire1906, wire1907, wire19879, wire1910, wire1912, wire1914, wire1940, wire19848, wire1945, wire19850, wire1951, wire1960, wire1961, wire1962, wire1968, wire1971, wire1972, wire19827, wire1976, wire1979, wire19770, wire1982, wire1983, wire1987, wire1990, wire19766, wire1991, wire19760, wire1992, wire1995, wire1996, wire1997, wire19759, wire1998, wire1999, wire2000, wire2004, wire19780, wire2026, wire19782, wire19783, wire2027, wire19778, wire2032, wire2041, wire2045, wire19727, wire19728, wire2062, wire19724, wire2068, wire2070, wire2078, wire19716, wire2079, wire19714, wire2099, wire2108, wire2119, wire2124, wire2125, wire2130, wire2134, wire2136, wire2139, wire2141, wire2146, wire2149, wire2153, wire2155, wire2156, wire2157, wire2163, wire2169, wire2174, wire2176, wire2179, wire19620, wire2180, wire2181, wire19605, wire2190, wire19607, wire19608, wire2191, wire19602, wire2195, wire2197, wire2205, wire19535, wire2269, wire19530, wire2277, wire19531, wire2278, wire19528, wire19529, wire2282, wire2283, wire2287, wire2290, wire2293, wire19519, wire2294, wire2295, wire2296, wire19486, wire2323, wire2324, wire19472, wire2335, wire2340, wire2343, wire2344, wire2345, wire2349, wire2350, wire19461, wire2351, wire19447, wire19448, wire2352, wire19449, wire19450, wire2353, wire19440, wire19441, wire19438, wire2359, wire19426, wire2364, wire19427, wire2365, wire2370, wire19424, wire2372, wire2374, wire19411, wire19412, wire2382, wire2384, wire2393, wire2398, wire2404, wire19387, wire2407, wire2410, wire2415, wire2417, wire2418, wire2424, wire2427, wire2428, wire2435, wire19339, wire2442, wire2448, wire19337, wire2449, wire2451, wire2452, wire2462, wire2463, wire19315, wire2464, wire19312, wire2468, wire2475, wire2480, wire19297, wire2481, wire19295, wire2487, wire2489, wire19290, wire19291, wire2490, wire19279, wire2493, wire2498, wire19246, wire2518, wire19245, wire2523, wire19243, wire2525, wire2526, wire2532, wire2537, wire2545, wire2548, wire19204, wire2557, wire2559, wire2560, wire19194, wire2565, wire2567, wire2568, wire2578, wire2579, wire2584, wire2588, wire2594, wire2598, wire19150, wire2599, wire2614, wire2615, wire19128, wire19129, wire2618, wire2630, wire19113, wire2634, wire19110, wire2635, wire2636, wire2645, wire2646, wire2657, wire2666, wire2669, wire2676, wire2679, wire2691, wire2692, wire19043, wire2700, wire19038, wire2703, wire2704, wire2705, wire19016, wire2712, wire2717, wire2720, wire2721, wire2724, wire2726, wire2728, wire19008, wire2729, wire2730, wire19006, wire2731, wire2733, wire2738, wire2739, wire18993, wire2740, wire2743, wire18992, wire2744, wire2748, wire18956, wire2775, wire18958, wire18959, wire2776, wire18944, wire18945, wire2785, wire2791, wire2797, wire2801, wire2802, wire2808, wire2809, wire2814, wire2815, wire2817, wire2825, wire18921, wire2828, wire2831, wire2842, wire2843, wire18894, wire2853, wire2865, wire2866, wire2870, wire18879, wire2875, wire2897, wire18859, wire18852, wire2910, wire18847, wire2914, wire2915, wire2939, wire18824, wire2940, wire18821, wire2943, wire2944, wire18810, wire2952, wire18811, wire2953, wire2958, wire2959, wire2964, wire18784, wire2970, wire2974, wire2975, wire2979, wire18771, wire2981, wire2995, wire3001, wire3006, wire3013, wire18744, wire3014, wire3015, wire3044, wire3059, wire3060, wire18696, wire3066, wire3067, wire3068, wire3069, wire3078, wire18687, wire3079, wire3080, wire18686, wire3081, wire3102, wire3111, wire3113, wire3123, wire3124, wire3135, wire18617, wire3136, wire18609, wire3142, wire3143, wire3154, wire3155, wire3195, wire3201, wire18529, wire3219, wire3222, wire18528, wire3223, wire3225, wire3229, wire3234, wire3244, wire3245, wire3256, wire3257, wire3258, wire3264, wire3271, wire3275, wire3279, wire18457, wire3280, wire3312, wire18416, wire3313, wire3325, wire3337, wire18394, wire3338, wire18386, wire3342, wire3353, wire3374, wire3375, wire3385, wire3392, wire3397, wire3404, wire3409, wire3415, wire3425, wire3435, wire3437, wire3438, wire3471, wire3479, wire3498, wire3515, wire18260, wire3516, wire3520, wire3524, wire3526, wire3531, wire3533, wire3550, wire3551, wire3563, wire18194, wire3570, wire3575, wire3580, wire18188, wire3581, wire3588, wire3607, wire3621, wire18157, wire3622, wire3624, wire3643, wire18117, wire3653, wire18111, wire18102, wire18103, wire18104, wire3662, wire18092, wire3665, wire18087, wire18088, wire3671, wire3676, wire18067, wire18068, wire18069, wire3685, wire18053, wire3690, wire3696, wire3700, wire3701, wire3702, wire3710, wire3723, wire3747, wire17993, wire3755, wire3759, wire3773, wire3774, wire3810, wire17940, wire17941, wire17942, wire3811, wire3828, wire17909, wire3829, wire17901, wire3835, wire3836, wire3850, wire3851, wire3866, wire3886, wire3887, wire3895, wire3896, wire3897, wire3899, wire3900, wire3901, wire3957, wire17808, wire3958, wire3964, wire3973, wire3990, wire17781, wire3991, wire3996, wire3998, wire4013, wire4020, wire4021, wire4026, wire4027, wire17739, wire4043, wire4048, wire4064, wire4065, wire4080, wire4088, wire4102, wire4103, wire4104, wire4113, wire4130, wire4143, wire4151, wire17632, wire4158, wire4159, wire4172, wire4185, wire4217, wire17591, wire4220, wire4221, wire4228, wire4229, wire4230, wire17569, wire4233, wire17570, wire4234, wire4252, wire4253, wire4263, wire4285, wire17535, wire4286, wire4291, wire4323, wire17468, wire4324, wire4343, wire17480, wire4344, wire4382, wire17447, wire4395, wire17448, wire4396, wire17428, wire4419, wire4427, wire4429, wire17391, wire4453, wire4454, wire4458, wire4459, wire17385, wire4470, wire4474, wire4475, wire4491, wire4496, wire17357, wire4500, wire4504, wire17349, wire17350, wire17352, wire17353, wire17343, wire4510, wire4520, wire17336, wire4523, wire4526, wire17324, wire4539, wire17317, wire4544, wire17319, wire4545, wire4548, wire4549, wire4550, wire4551, wire17310, wire4568, wire4569, wire17292, wire4572, wire17294, wire17295, wire4573, wire4576, wire17287, wire4581, wire4591, wire4602, wire4628, wire4638, wire4639, wire4644, wire4649, wire17224, wire4651, wire4655, wire17215, wire4662, wire4663, wire4669, wire4671, wire4676, wire4684, wire4685, wire4735, wire4743, wire4750, wire4752, wire4753, wire4765, wire4768, wire4780, wire4786, wire4805, wire4818, wire17089, wire4819, wire4820, wire4821, wire17074, wire4822, wire4827, wire4828, wire4831, wire4832, wire4838, wire4839, wire4857, wire4858, wire4859, wire17052, wire4860, wire4863, wire4888, wire4890, wire4891, wire4900, wire4904, wire4905, wire4908, wire4919, wire4924, wire4933, wire4937, wire4941, wire16988, wire4942, wire4950, wire16972, wire4953, wire16964, wire4961, wire16946, wire4982, wire4986, wire16940, wire4993, wire4998, wire16908, wire16909, wire5067, wire5068, wire16861, wire16857, wire16863, wire16865, wire16867, wire16871, wire16884, wire16885, wire16888, wire16889, wire16890, wire16892, wire16896, wire16910, wire16924, wire16929, wire16930, wire16936, wire16941, wire16943, wire16950, wire16957, wire16960, wire16962, wire16966, wire16968, wire16976, wire16990, wire16991, wire16993, wire16994, wire16995, wire16996, wire16997, wire17001, wire17003, wire17016, wire17028, wire17038, wire17039, wire17041, wire17042, wire17044, wire17045, wire17047, wire17053, wire17055, wire17056, wire17058, wire17060, wire17061, wire17063, wire17067, wire17071, wire17076, wire17079, wire17093, wire17094, wire17096, wire17106, wire17108, wire17109, wire17114, wire17115, wire17116, wire17117, wire17119, wire17121, wire17122, wire17123, wire17125, wire17127, wire17128, wire17129, wire17134, wire17136, wire17137, wire17140, wire17141, wire17145, wire17146, wire17152, wire17153, wire17154, wire17156, wire17158, wire17166, wire17170, wire17172, wire17174, wire17181, wire17184, wire17185, wire17187, wire17191, wire17193, wire17196, wire17201, wire17202, wire17203, wire17206, wire17209, wire17212, wire17220, wire17226, wire17231, wire17239, wire17241, wire17243, wire17245, wire17246, wire17247, wire17251, wire17265, wire17266, wire17271, wire17275, wire17276, wire17280, wire17281, wire17284, wire17285, wire17288, wire17289, wire17290, wire17291, wire17297, wire17298, wire17299, wire17301, wire17309, wire17325, wire17337, wire17338, wire17359, wire17360, wire17363, wire17364, wire17365, wire17377, wire17382, wire17383, wire17384, wire17388, wire17389, wire17390, wire17392, wire17393, wire17394, wire17397, wire17398, wire17400, wire17405, wire17417, wire17418, wire17433, wire17434, wire17435, wire17436, wire17439, wire17440, wire17441, wire17443, wire17446, wire17450, wire17452, wire17453, wire17454, wire17456, wire17457, wire17458, wire17459, wire17462, wire17465, wire17467, wire17469, wire17484, wire17493, wire17499, wire17504, wire17505, wire17507, wire17509, wire17513, wire17516, wire17518, wire17537, wire17541, wire17542, wire17543, wire17545, wire17548, wire17549, wire17550, wire17555, wire17557, wire17558, wire17559, wire17560, wire17562, wire17565, wire17568, wire17574, wire17575, wire17578, wire17579, wire17581, wire17585, wire17592, wire17593, wire17594, wire17596, wire17599, wire17605, wire17606, wire17608, wire17610, wire17622, wire17626, wire17627, wire17629, wire17631, wire17635, wire17638, wire17639, wire17640, wire17646, wire17647, wire17650, wire17651, wire17654, wire17656, wire17659, wire17660, wire17662, wire17663, wire17667, wire17668, wire17672, wire17674, wire17677, wire17679, wire17681, wire17684, wire17685, wire17686, wire17688, wire17690, wire17691, wire17692, wire17693, wire17695, wire17696, wire17698, wire17700, wire17701, wire17704, wire17705, wire17706, wire17708, wire17709, wire17710, wire17712, wire17721, wire17725, wire17732, wire17735, wire17740, wire17744, wire17746, wire17748, wire17750, wire17753, wire17757, wire17760, wire17761, wire17764, wire17765, wire17772, wire17773, wire17776, wire17778, wire17779, wire17783, wire17786, wire17796, wire17800, wire17801, wire17806, wire17810, wire17813, wire17816, wire17817, wire17818, wire17819, wire17821, wire17822, wire17824, wire17825, wire17826, wire17827, wire17830, wire17837, wire17840, wire17844, wire17845, wire17850, wire17852, wire17853, wire17854, wire17858, wire17864, wire17865, wire17868, wire17870, wire17872, wire17873, wire17887, wire17889, wire17891, wire17893, wire17894, wire17906, wire17908, wire17911, wire17916, wire17931, wire17955, wire17963, wire17964, wire17965, wire17976, wire17985, wire17987, wire17988, wire17989, wire17995, wire17996, wire17999, wire18000, wire18001, wire18003, wire18010, wire18012, wire18013, wire18017, wire18018, wire18019, wire18021, wire18023, wire18026, wire18027, wire18035, wire18036, wire18071, wire18074, wire18075, wire18076, wire18085, wire18089, wire18096, wire18097, wire18098, wire18106, wire18107, wire18120, wire18128, wire18129, wire18132, wire18134, wire18136, wire18145, wire18158, wire18159, wire18160, wire18161, wire18163, wire18164, wire18178, wire18182, wire18185, wire18187, wire18190, wire18191, wire18193, wire18196, wire18201, wire18202, wire18205, wire18209, wire18210, wire18220, wire18221, wire18222, wire18232, wire18234, wire18237, wire18238, wire18243, wire18245, wire18252, wire18264, wire18266, wire18268, wire18269, wire18270, wire18278, wire18287, wire18290, wire18294, wire18295, wire18300, wire18307, wire18318, wire18321, wire18324, wire18325, wire18328, wire18334, wire18348, wire18353, wire18358, wire18370, wire18371, wire18372, wire18388, wire18393, wire18397, wire18398, wire18401, wire18403, wire18409, wire18411, wire18414, wire18418, wire18420, wire18422, wire18429, wire18433, wire18434, wire18445, wire18452, wire18471, wire18474, wire18475, wire18476, wire18482, wire18487, wire18488, wire18492, wire18493, wire18495, wire18496, wire18504, wire18507, wire18509, wire18510, wire18533, wire18537, wire18541, wire18546, wire18548, wire18562, wire18564, wire18575, wire18576, wire18586, wire18587, wire18588, wire18596, wire18598, wire18600, wire18602, wire18603, wire18605, wire18607, wire18608, wire18614, wire18616, wire18619, wire18631, wire18632, wire18637, wire18638, wire18641, wire18642, wire18646, wire18650, wire18652, wire18655, wire18656, wire18663, wire18665, wire18668, wire18669, wire18670, wire18671, wire18677, wire18679, wire18688, wire18691, wire18692, wire18694, wire18701, wire18702, wire18703, wire18704, wire18705, wire18709, wire18714, wire18715, wire18718, wire18726, wire18732, wire18735, wire18737, wire18749, wire18750, wire18755, wire18757, wire18760, wire18761, wire18763, wire18767, wire18768, wire18770, wire18776, wire18777, wire18786, wire18788, wire18793, wire18801, wire18804, wire18812, wire18815, wire18816, wire18826, wire18828, wire18833, wire18837, wire18838, wire18839, wire18841, wire18845, wire18846, wire18850, wire18854, wire18855, wire18871, wire18877, wire18878, wire18882, wire18883, wire18884, wire18885, wire18889, wire18890, wire18891, wire18895, wire18911, wire18913, wire18914, wire18916, wire18917, wire18918, wire18919, wire18922, wire18923, wire18924, wire18925, wire18926, wire18928, wire18930, wire18931, wire18932, wire18934, wire18936, wire18941, wire18943, wire18947, wire18949, wire18951, wire18955, wire18965, wire18968, wire18969, wire18970, wire18971, wire18972, wire18973, wire18976, wire18985, wire18991, wire18998, wire19003, wire19005, wire19010, wire19011, wire19015, wire19025, wire19027, wire19031, wire19034, wire19048, wire19050, wire19054, wire19057, wire19062, wire19063, wire19069, wire19076, wire19077, wire19078, wire19079, wire19083, wire19084, wire19087, wire19089, wire19090, wire19098, wire19103, wire19104, wire19106, wire19109, wire19118, wire19123, wire19125, wire19127, wire19130, wire19134, wire19146, wire19147, wire19148, wire19153, wire19158, wire19164, wire19169, wire19178, wire19182, wire19186, wire19189, wire19190, wire19193, wire19200, wire19202, wire19208, wire19210, wire19212, wire19213, wire19216, wire19220, wire19227, wire19232, wire19234, wire19238, wire19239, wire19241, wire19249, wire19256, wire19263, wire19268, wire19270, wire19272, wire19273, wire19276, wire19278, wire19281, wire19285, wire19286, wire19294, wire19301, wire19302, wire19304, wire19306, wire19307, wire19308, wire19309, wire19310, wire19316, wire19317, wire19324, wire19325, wire19326, wire19332, wire19338, wire19343, wire19344, wire19346, wire19347, wire19351, wire19354, wire19355, wire19359, wire19362, wire19363, wire19364, wire19366, wire19368, wire19369, wire19370, wire19376, wire19380, wire19381, wire19389, wire19393, wire19395, wire19396, wire19400, wire19401, wire19402, wire19403, wire19405, wire19406, wire19409, wire19423, wire19429, wire19431, wire19437, wire19454, wire19455, wire19456, wire19466, wire19471, wire19479, wire19485, wire19491, wire19494, wire19496, wire19497, wire19498, wire19499, wire19513, wire19520, wire19521, wire19527, wire19536, wire19538, wire19539, wire19541, wire19542, wire19543, wire19544, wire19545, wire19548, wire19549, wire19552, wire19567, wire19576, wire19580, wire19581, wire19589, wire19603, wire19610, wire19612, wire19613, wire19623, wire19629, wire19636, wire19638, wire19644, wire19645, wire19646, wire19647, wire19648, wire19650, wire19652, wire19653, wire19656, wire19658, wire19659, wire19666, wire19667, wire19668, wire19670, wire19671, wire19674, wire19676, wire19677, wire19680, wire19687, wire19691, wire19693, wire19694, wire19695, wire19698, wire19702, wire19704, wire19706, wire19707, wire19708, wire19710, wire19717, wire19718, wire19722, wire19725, wire19726, wire19730, wire19731, wire19733, wire19734, wire19735, wire19738, wire19739, wire19746, wire19747, wire19750, wire19752, wire19756, wire19757, wire19758, wire19765, wire19769, wire19775, wire19777, wire19779, wire19792, wire19800, wire19801, wire19802, wire19803, wire19804, wire19807, wire19808, wire19813, wire19823, wire19825, wire19828, wire19829, wire19830, wire19834, wire19837, wire19839, wire19841, wire19842, wire19843, wire19845, wire19858, wire19861, wire19867, wire19875, wire19876, wire19878, wire19880, wire19884, wire19886, wire19887, wire19890, wire19891, wire19893, wire19898, wire19904, wire19907, wire19909, wire19910, wire19911, wire19917, wire19920, wire19923, wire19925, wire19926, wire19930, wire19938, wire19939, wire19943, wire19944, _86, _87, _143, _217, _252, _255, _285, _288, _314, _317, _360, _409, _422, _425, _453, _461, _462, _465, _499, _511, _596, _635, _636, _696, _699, _745, _778, _823, _969, _976, _1018, _1021, _1126, _1129, _1208, _1211, _1239, _1242, _1262, _1263, _1264, _1265, _1289, _1307, _1308, _1347, _1401, _1404, _1411, _1414, _1455, _1516, _1517, _1519, _1533, _1544, _1549, _1581, _1643, _1648, _1676, _1679, _1721, _1845, _1846, _1848, _1849, _1862, _1871, _1972, _1978, _1990, _1992, _1993, _2020, _2023, _2026, _2056, _2059, _2060, _2071, _2123, _2126, _2182, _2199, _2250, _2264, _2265, _2270, _2332, _2335, _2519, _2561, _2581, _2591, _2594, _2597, _2661, _2679, _2726, _2729, _2737, _2738, _2740, _2752, _2775, _2778, _2781, _2784, _2787, _2858, _2863, _2866, _2884, _2890, _2894, _2901, _2906, _2909, _2912, _2919, _2938, _2970, _2973, _2976, _2981, _2990, _2993, _3004, _3007, _3035, _3077, _3082, _3089, _3092, _3095, _3098, _3109, _3110, _3112, _3127, _3149, _3158, _3273, _3304, _3312, _3332, _3335, _3344, _3392, _3429, _3430, _3440, _3486, _3568, _3637, _3638, _3639, _3809, _3810, _3811, _3812, _3827, _3899, _3948, _4048, _4072, _4088, _4188, _4253, _4363, _4473, _4479, _4492, _4495, _4527, _4585, _4657, _4707, _4718, _4739, _4740, _4890, _4924, _4944, _4984, _4987, _4992, _5193, _5201, _5204, _5207, _5208, _5289, _5329, _5528, _5529, _5561, _5601, _5628, _5825, _5873, _5959, _5996, _28911, _28939, _29017, _29024, _29028, _29046, _29052, _29053, _29117, _29131, _29155, _29156, _29181, _29189, _29191, _29192, _29193, _29197, _29204, _29206, _29207, _29210, _29212, _29222, _29234, _29252, _29269, _29274, _29276, _29298, _29305, _29309, _29313, _29315, _29327, _29332, _29343, _29353, _29356, _29375, _29379, _29381, _29383, _29386, _29424, _29427, _29429, _29431, _29448, _29458, _29464, _29471, _29472, _29474, _29477, _29478, _29479, _29480, _29539, _29544, _29545, _29607, _29608, _29611, _29613, _29641, _29643, _29645, _29649, _29651, _29653, _29659, _29694, _29711, _29722, _29731, _29755, _29771, _29772, _29782, _29784, _29832, _29849, _29851, _29864, _29870, _29885, _29886, _29890, _29895, _29896, _29897, _29898, _29899, _29900, _29904, _29913, _29934, _29936, _29938, _29962, _29963, _30001, _30030, _30031, _30032, _30036, _30037, _30039, _30040, _30042, _30050, _30071, _30073, _30076, _30081, _30087, _30101, _30102, _30108, _30113, _30119, _30120, _30153, _30155, _30162, _30163, _30166, _30172, _30175, _30176, _30194, _30195, _30198, _30203, _30206, _30217, _30218, _30221, _30224, _30229, _30240, _30242, _30244, _30248, _30250, _30273, _30296, _30322, _30323, _30347, _30353, _30358, _30359, _30362, _30371, _30385, _30386, _30390, _30391, _30395, _30401, _30404, _30450, _30453, _30455, _30457, _30468, _30471, _30482, _30484, _30488, _30490, _30491, _30495, _30497, _30546, _30549, _30553, _30557, _30561, _30565, _30568, _30569, _30571, _30578, _30595, _30599, _30604, _30607, _30622, _30623, _30650, _30652, _30656, _30657, _30659, _30665, _30668, _30673, _30694, _30702, _30703, _30710, _30763, _30765, _30792, _30794, _30798, _30799, _30811, _30816, _30817, _30819, _30821, _30824, _30833, _30839, _30848, _30850, _30851, _30861, _30865, _30866, _30869, _30896, _30923, _30926, _30948, _30950, _30958, _30959, _30964, _30973, _30974, _30980, _30983, _30984, _30987, _30988, _31018, _31021, _31022, _31026, _31044, _31045, _31049, _31050, _31059, _31078, _31080, _31081, _31082, _31115, _31116, _31117, _31127, _31128, _31132, _31135, _31139, _31143, _31145, _31151, _31153, _31166, _31167, _31173, _31175, _31176, _31182, _31186, _31188, _31190, _31193, _31195, _31197, _31199, _31203, _31214, _31216, _31219, _31221, _31223, _31229, _31237, _31238, _31243, _31251, _31262, _31264, _31266, _31270, _31272, _31276, _31278, _31279, _31280, _31283, _31285, _31286, _31297, _31298, _31302, _31305, _31318, _31319, _31321, _31328, _31330, _31334, _31338, _31340, _31342, _31343, _31356, _31360, _31365, _31368, _31372, _31374, _31376, _31377, _31378, _31381, _31382, _31392, _31423, _31433, _31435, _31437, _31442, _31445, _31446, _31450, _31455, _31468, _31494, _31496, _31512, _31554, _31555, _31567, _31569, _31572, _31586, _31588, _31592, _31594, _31600, _31614, _31615, _31624, _31632, _31662, _31663, _31664, _31754, _31770, _31801, _31819, _31826, _31830, _31832, _31833, _31834, _31883, _31887, _31890, _31892, _31894, _31899, _31900, _31910, _31923, _31932, _31940, _31946, _31961, _31977, _31978, _31998, _32003, _32019, _32025, _32040, _32062, _32066, _32068, _32081, _32090, _32094, _32108, _32110, _32114, _32115, _32140, _32141, _32149, _32161, _32183, _32185, _32227, _32230, _32240, _32241, _32250, _32288, _32293, _32297, _32302, _32304, _32314, _32327, _32330, _32331, _32341, _32343, _32344, _32351, _32363, _32372, _32380, _32382, _32401, _32406, _32408, _32410, _32412, _32417, _32419, _32421, _32426, _32437, _32442, _32447, _32450, _32452, _32454, _32472, _32474, _32477, _32478, _32488, _32495, _32504, _32509, _32510, _32514, _32515, _32516, _32521, _32526, _32529, _32536, _32540, _32541, _32548, _32550, _32554, _32558, _32562, _32577, _32580, _32583, _32603, _32625, _32636, _32643, _32647, _32649, _32651, _32652, _32654, _32657, _32665, _32666, _32675, _32677, _32682, _32695, _32697, _32719, _32764, _32769, _32771, _32772, _32802, _32808, _32812, _32815, _32818, _32832, _32837, _32839, _32841, _32844, _32845, _32856, _32877, _32880, _32881, _32918, _32919, _32920, _32999, _33004, _33013, _33033, _33038, _33048, _33099, _33101, _33104, _33117, _33122, _33138, _33161, _33162, _33163, _33164, _33165, _33185, _33212, _33214, _33216, _33217, _33218, _33220, _33223, _33239, _33261, _33275, _33286, _33287, _33291, _33293, _33351, _33353, _33354, _33361, _33362, _33400, _33401, _33461, _33464, _33477, _33487, _33489, _33493, _33495, _33496, _33497, _33528, _33535, _33537, _33543, _33561, _33568, _33578, _33612, _33614, _33626, _33656, _33658, _33659, _33662, _33670, _33681, _33709, _33710;

assign o_1_ = ( wire388 ) | ( wire16865 ) | ( wire16867 ) | ( _28939 ) ;
 assign o_19_ = ( n_n5144 ) | ( wire736  &  wire16876 ) ;
 assign o_2_ = ( wire16877 ) | ( wire736  &  n_n162 ) ;
 assign o_0_ = ( n_n231 ) | ( wire16886 ) | ( _5996 ) | ( _29024 ) ;
 assign o_29_ = ( wire5026 ) | ( wire5027 ) | ( wire16911 ) ;
 assign o_39_ = ( n_n4721 ) | ( wire16933 ) ;
 assign o_38_ = ( _29478 ) | ( _29479 ) ;
 assign o_25_ = ( n_n5144 ) | ( n_n159  &  _29480 ) ;
 assign o_12_ = ( wire17405 ) | ( _30030 ) | ( _30032 ) ;
 assign o_37_ = ( n_n4103 ) | ( n_n4102 ) | ( _30250 ) ;
 assign o_26_ = ( wire17601 ) | ( wire17602 ) | ( _30296 ) ;
 assign o_11_ = ( wire17604 ) | ( wire17612 ) | ( _4363 ) ;
 assign o_36_ = ( wire17849 ) | ( wire17698 ) | ( wire17779 ) | ( _30457 ) ;
 assign o_27_ = ( wire17861 ) | ( wire17862 ) | ( _30599 ) ;
 assign o_14_ = ( wire17876 ) | ( wire17877 ) | ( wire17913 ) | ( wire17915 ) ;
 assign o_35_ = ( n_n3451 ) | ( _30821 ) | ( _30869 ) ;
 assign o_28_ = ( n_n2998 ) | ( wire18154 ) | ( wire18155 ) | ( wire18167 ) ;
 assign o_13_ = ( wire18213 ) | ( n_n3033 ) | ( _30950 ) | ( _30959 ) ;
 assign o_34_ = ( n_n3029 ) | ( wire18290 ) | ( _31045 ) | ( _31059 ) ;
 assign o_21_ = ( wire18299 ) | ( n_n10  &  wire185 ) | ( n_n10  &  wire270 ) ;
 assign o_16_ = ( n_n2721 ) | ( wire3442 ) | ( wire18310 ) | ( wire18311 ) ;
 assign o_40_ = ( n_n5144 ) | ( wire3439 ) | ( n_n135  &  wire267 ) ;
 assign o_33_ = ( n_n259 ) | ( wire18323 ) | ( wire18329 ) | ( wire18330 ) ;
 assign o_22_ = ( n_n5144 ) | ( _31116 ) | ( wire267  &  _31115 ) ;
 assign o_15_ = ( wire18354 ) | ( wire18355 ) | ( _31145 ) ;
 assign o_32_ = ( n_n3170 ) | ( wire18488 ) | ( _31280 ) | ( _31283 ) ;
 assign o_23_ = ( wire18495 ) | ( wire18507 ) | ( _31321 ) | ( _31328 ) ;
 assign o_18_ = ( wire18548 ) | ( wire18562 ) | ( _31378 ) | ( _31381 ) ;
 assign o_31_ = ( wire3194 ) | ( wire18568 ) | ( wire18572 ) ;
 assign o_24_ = ( n_n5144 ) | ( n_n159  &  _31392 ) ;
 assign o_17_ = ( n_n2748 ) | ( wire18621 ) | ( wire18623 ) ;
 assign o_43_ = ( wire18685 ) | ( _31496 ) ;
 assign o_30_ = ( wire18292 ) | ( n_n3033 ) | ( _30950 ) | ( _31555 ) ;
 assign o_44_ = ( n_n4845 ) | ( wire18795 ) | ( wire18737 ) | ( _31600 ) ;
 assign o_41_ = ( n_n5144 ) | ( wire2962 ) ;
 assign o_42_ = ( wire18802 ) | ( wire18803 ) | ( wire18807 ) ;
 assign o_20_ = ( n_n5144 ) | ( wire736  &  wire18809 ) ;
 assign o_45_ = ( wire18437 ) | ( wire18490 ) | ( _31664 ) ;
 assign o_10_ = ( wire19030 ) | ( wire19025 ) | ( _31890 ) | ( _32185 ) ;
 assign o_9_ = ( wire19349 ) | ( wire19459 ) | ( _32697 ) ;
 assign o_7_ = ( wire19677 ) | ( wire19680 ) | ( _33101 ) | ( _33165 ) ;
 assign o_8_ = ( i_3_  &  (~ i_1_)  &  i_2_  &  (~ i_0_) ) | ( i_3_  &  (~ i_1_)  &  (~ i_2_)  &  (~ i_0_) ) ;
 assign o_5_ = ( wire19813 ) | ( wire19861 ) | ( _33537 ) | ( _33662 ) ;
 assign o_6_ = ( wire19922 ) | ( _86 ) | ( _87 ) ;
 assign o_3_ = ( n_n259 ) | ( wire18323 ) | ( wire19928 ) ;
 assign o_4_ = ( n_n275 ) | ( wire441 ) | ( wire19941 ) | ( wire19946 ) ;
 assign wire5057 = ( n_n35  &  wire5067  &  wire16861 ) | ( n_n35  &  wire5068  &  wire16861 ) ;
 assign wire16872 = ( wire428 ) | ( wire16871 ) ;
 assign n_n5144 = ( i_2_  &  (~ i_0_) ) | ( i_3_  &  (~ i_1_)  &  (~ i_2_)  &  (~ i_0_) ) ;
 assign wire736 = ( n_n184  &  n_n163  &  wire725  &  n_n35 ) ;
 assign wire16876 = ( i_5_  &  i_3_  &  (~ i_4_) ) ;
 assign n_n162 = ( i_5_  &  (~ i_3_)  &  (~ i_4_) ) ;
 assign wire16877 = ( n_n5144 ) | ( n_n184  &  wire725  &  wire16857 ) ;
 assign wire16898 = ( i_2_  &  (~ i_0_) ) | ( i_3_  &  (~ i_1_)  &  (~ i_2_)  &  i_0_ ) | ( i_3_  &  (~ i_1_)  &  (~ i_2_)  &  (~ i_0_) ) ;
 assign wire5026 = ( n_n5  &  n_n65 ) | ( n_n65  &  wire398 ) | ( n_n65  &  wire16908 ) ;
 assign wire5027 = ( n_n5  &  wire343 ) | ( wire343  &  wire16908 ) | ( wire343  &  wire16909 ) ;
 assign wire16911 = ( wire16910 ) | ( _5959 ) | ( n_n12  &  _29046 ) ;
 assign n_n4721 = ( wire244  &  n_n39 ) | ( n_n38  &  wire1595 ) | ( n_n39  &  wire1595 ) ;
 assign wire16933 = ( n_n373 ) | ( n_n374 ) | ( wire16929 ) | ( wire16930 ) ;
 assign n_n4399 = ( wire17149 ) | ( wire17121 ) | ( wire17140 ) | ( _29343 ) ;
 assign n_n17 = ( i_7_  &  (~ i_6_) ) ;
 assign n_n159 = ( i_1_  &  (~ i_2_)  &  (~ i_0_) ) ;
 assign n_n4103 = ( n_n4112 ) | ( wire17513 ) | ( _30101 ) | ( _30102 ) ;
 assign n_n4102 = ( n_n4109 ) | ( wire17565 ) | ( _30162 ) | ( _30163 ) ;
 assign wire17601 = ( wire4228 ) | ( wire4229 ) | ( wire17599 ) ;
 assign wire17602 = ( wire4217 ) | ( wire4221 ) | ( wire17592 ) | ( wire17593 ) ;
 assign n_n4 = ( n_n159  &  n_n35  &  n_n111 ) ;
 assign wire17604 = ( n_n4  &  n_n71 ) | ( n_n13  &  wire1496 ) ;
 assign wire17612 = ( wire17605 ) | ( wire17606 ) | ( wire17608 ) | ( wire17610 ) ;
 assign wire17849 = ( wire17844 ) | ( wire17845 ) | ( _30561 ) ;
 assign wire17861 = ( wire3900 ) | ( wire3901 ) | ( wire17852 ) | ( wire17853 ) ;
 assign wire17862 = ( wire3895 ) | ( wire3896 ) | ( wire3897 ) | ( wire17854 ) ;
 assign wire17876 = ( wire584 ) | ( wire3866 ) | ( wire17872 ) | ( wire17873 ) ;
 assign wire17877 = ( wire17868 ) | ( wire17870 ) | ( _30607 ) ;
 assign wire17913 = ( wire3828 ) | ( wire3829 ) | ( wire17911 ) ;
 assign wire17915 = ( n_n2622 ) | ( wire3836 ) | ( wire17906 ) | ( wire17908 ) ;
 assign wire18141 = ( n_n3482 ) | ( wire3773 ) | ( _30665 ) | ( _30668 ) ;
 assign wire18142 = ( wire18000 ) | ( wire18001 ) | ( wire18026 ) | ( wire18027 ) ;
 assign wire18148 = ( n_n3454 ) | ( n_n3456 ) | ( wire18145 ) | ( _30866 ) ;
 assign n_n2998 = ( wire3628 ) | ( wire3629 ) | ( wire18150 ) ;
 assign wire18154 = ( wire3624 ) | ( n_n218  &  n_n19  &  n_n157 ) ;
 assign wire18155 = ( n_n7241 ) | ( n_n17  &  wire743 ) | ( n_n17  &  wire1524 ) ;
 assign wire18167 = ( wire3621 ) | ( wire3622 ) | ( wire18163 ) | ( wire18164 ) ;
 assign wire18212 = ( wire18209 ) | ( wire18210 ) | ( n_n46  &  wire1271 ) ;
 assign wire18213 = ( wire18185 ) | ( wire18187 ) | ( _30926 ) ;
 assign wire18214 = ( wire18212 ) | ( wire18185 ) | ( wire18187 ) | ( _30926 ) ;
 assign wire18292 = ( n_n3029 ) | ( wire18245 ) | ( _31044 ) | ( _31045 ) ;
 assign wire18297 = ( wire3469 ) | ( wire3470 ) | ( wire18294 ) | ( wire18295 ) ;
 assign n_n10 = ( n_n162  &  n_n159  &  n_n161 ) ;
 assign wire185 = ( wire729  &  n_n149 ) | ( wire730  &  n_n149 ) | ( wire717  &  n_n149 ) ;
 assign wire270 = ( wire729  &  n_n191 ) | ( wire730  &  n_n191 ) | ( wire717  &  n_n191 ) ;
 assign wire18299 = ( n_n5144 ) | ( n_n51  &  wire751 ) | ( n_n51  &  wire18298 ) ;
 assign n_n2721 = ( wire675 ) | ( wire3451 ) | ( wire18301 ) | ( wire18302 ) ;
 assign wire3442 = ( n_n162  &  n_n220  &  n_n200  &  wire767 ) ;
 assign wire18310 = ( wire587 ) | ( wire18307 ) | ( n_n32  &  wire124 ) ;
 assign wire18311 = ( n_n2728 ) | ( wire18300 ) | ( _31082 ) ;
 assign n_n135 = ( (~ i_9_)  &  (~ i_10_)  &  (~ i_11_)  &  wire725 ) ;
 assign wire267 = ( n_n159  &  n_n111  &  wire747 ) | ( n_n159  &  n_n111  &  n_n126 ) ;
 assign wire3439 = ( wire185  &  n_n6 ) | ( wire270  &  n_n6 ) | ( n_n6  &  wire372 ) ;
 assign n_n259 = ( wire3433 ) | ( wire3434 ) | ( wire18316 ) ;
 assign wire18323 = ( n_n7252 ) | ( wire389 ) | ( wire3425 ) | ( wire18321 ) ;
 assign wire18329 = ( wire3415 ) | ( wire18325 ) | ( n_n10  &  wire145 ) ;
 assign wire18330 = ( wire3437 ) | ( wire3438 ) | ( wire18328 ) ;
 assign n_n14 = ( n_n159  &  n_n48  &  n_n161 ) ;
 assign wire18354 = ( wire3385 ) | ( wire18348 ) | ( _3158 ) | ( _31132 ) ;
 assign wire18355 = ( wire18353 ) | ( _3149 ) | ( _31139 ) | ( _31143 ) ;
 assign n_n3166 = ( n_n3179 ) | ( n_n3176 ) | ( _31175 ) | ( _31176 ) ;
 assign wire18437 = ( wire18403 ) | ( wire18422 ) | ( _31223 ) ;
 assign wire18490 = ( n_n3170 ) | ( wire18452 ) | ( _31279 ) | ( _31280 ) ;
 assign wire18499 = ( wire454 ) | ( wire3245 ) | ( wire18496 ) ;
 assign wire18512 = ( wire708 ) | ( wire3234 ) | ( wire18510 ) ;
 assign wire18526 = ( wire3225 ) | ( _2912 ) | ( _2919 ) | ( _31330 ) ;
 assign wire18565 = ( wire4323 ) | ( wire4324 ) | ( wire18564 ) ;
 assign wire3194 = ( i_7_  &  i_6_  &  n_n159  &  _31382 ) ;
 assign wire18568 = ( n_n5144 ) | ( n_n159  &  n_n218  &  n_n18 ) ;
 assign wire18572 = ( wire430 ) | ( n_n5319 ) | ( wire684 ) | ( wire3195 ) ;
 assign n_n16 = ( (~ i_7_)  &  i_6_ ) ;
 assign n_n2748 = ( n_n4441 ) | ( wire575 ) | ( wire18577 ) | ( wire18578 ) ;
 assign wire18621 = ( wire3135 ) | ( wire3136 ) | ( wire18619 ) ;
 assign wire18623 = ( n_n2747 ) | ( wire3143 ) | ( wire18614 ) | ( wire18616 ) ;
 assign wire18682 = ( wire4933 ) | ( _31433 ) | ( n_n101  &  _29383 ) ;
 assign wire18683 = ( wire18638 ) | ( wire18677 ) | ( _31442 ) ;
 assign wire18685 = ( wire18655 ) | ( wire18656 ) | ( wire18670 ) | ( wire18671 ) ;
 assign n_n4845 = ( wire2977 ) | ( wire18783 ) | ( wire18789 ) | ( wire18790 ) ;
 assign wire18795 = ( wire18682 ) | ( wire18683 ) | ( wire18685 ) | ( wire18793 ) ;
 assign wire2962 = ( n_n162  &  n_n184  &  n_n163  &  n_n161 ) ;
 assign wire18802 = ( wire4354 ) | ( wire4355 ) | ( wire4827 ) | ( wire4828 ) ;
 assign wire18803 = ( n_n6271 ) | ( n_n6267 ) | ( n_n6270 ) | ( n_n6269 ) ;
 assign wire18807 = ( wire419 ) | ( wire445 ) | ( wire18801 ) | ( wire18804 ) ;
 assign wire18809 = ( (~ i_5_)  &  i_3_  &  i_4_ ) ;
 assign wire19030 = ( n_n1800 ) | ( n_n1799 ) | ( n_n1801 ) | ( wire19027 ) ;
 assign wire19349 = ( wire19212 ) | ( wire19278 ) | ( _32454 ) ;
 assign wire19459 = ( wire19127 ) | ( wire19454 ) | ( _32695 ) ;
 assign wire19869 = ( wire19738 ) | ( wire19739 ) | ( wire19757 ) | ( wire19758 ) ;
 assign wire19914 = ( wire19893 ) | ( wire19909 ) | ( _33658 ) | ( _33659 ) ;
 assign n_n5 = ( n_n159  &  n_n124  &  n_n111 ) ;
 assign wire19922 = ( wire454 ) | ( wire19920 ) | ( wire742  &  wire779 ) ;
 assign wire19928 = ( wire467 ) | ( wire19925 ) | ( wire19926 ) ;
 assign n_n275 = ( wire525 ) | ( n_n7266 ) | ( wire19929 ) | ( wire19933 ) ;
 assign wire441 = ( _33710 ) | ( n_n3  &  wire95 ) | ( n_n3  &  _33709 ) ;
 assign wire19941 = ( n_n7260 ) | ( wire439 ) | ( wire19938 ) | ( wire19939 ) ;
 assign wire19946 = ( wire707 ) | ( wire138 ) | ( wire19944 ) ;
 assign n_n219 = ( (~ i_1_)  &  (~ i_2_)  &  i_0_ ) ;
 assign n_n218 = ( (~ i_5_)  &  (~ i_3_)  &  i_4_ ) ;
 assign wire428 = ( (~ i_7_)  &  i_6_  &  n_n219  &  n_n218 ) | ( i_7_  &  (~ i_6_)  &  n_n219  &  n_n218 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n219  &  n_n218 ) ;
 assign n_n184 = ( (~ i_9_)  &  (~ i_10_)  &  (~ i_11_) ) ;
 assign n_n163 = ( i_1_  &  (~ i_2_)  &  i_0_ ) ;
 assign wire725 = ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  (~ i_15_) ) ;
 assign n_n35 = ( (~ i_7_)  &  (~ i_8_)  &  (~ i_6_) ) ;
 assign wire729 = ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  (~ i_15_) ) ;
 assign n_n65 = ( (~ i_9_)  &  i_10_  &  (~ i_11_)  &  wire729 ) ;
 assign n_n71 = ( i_9_  &  i_10_  &  (~ i_11_)  &  wire729 ) ;
 assign n_n124 = ( (~ i_7_)  &  (~ i_8_)  &  i_6_ ) ;
 assign n_n9 = ( n_n162  &  n_n159  &  n_n124 ) ;
 assign wire343 = ( i_9_  &  i_10_  &  (~ i_11_)  &  wire729 ) | ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire729 ) ;
 assign n_n48 = ( i_5_  &  (~ i_3_)  &  i_4_ ) ;
 assign n_n220 = ( (~ i_1_)  &  (~ i_2_)  &  (~ i_0_) ) ;
 assign n_n38 = ( n_n124  &  n_n48  &  n_n220 ) ;
 assign wire244 = ( n_n156  &  wire720 ) | ( n_n156  &  wire723 ) | ( n_n156  &  wire727 ) ;
 assign wire5024 = ( n_n39  &  wire235 ) | ( n_n39  &  wire236 ) ;
 assign n_n373 = ( wire5024 ) | ( n_n38  &  wire244 ) ;
 assign wire140 = ( i_15_  &  n_n156  &  n_n205 ) | ( (~ i_15_)  &  n_n156  &  n_n205 ) | ( (~ i_15_)  &  n_n156  &  n_n211 ) ;
 assign n_n39 = ( n_n48  &  n_n220  &  n_n126 ) ;
 assign wire5022 = ( n_n38  &  wire235 ) | ( n_n38  &  wire236 ) ;
 assign n_n374 = ( wire5022 ) | ( wire140  &  n_n39 ) ;
 assign n_n134 = ( i_9_  &  (~ i_10_)  &  i_11_  &  wire719 ) ;
 assign n_n132 = ( (~ i_9_)  &  (~ i_10_)  &  i_11_  &  wire719 ) ;
 assign n_n969 = ( n_n39  &  n_n134 ) | ( n_n38  &  n_n132 ) | ( n_n39  &  n_n132 ) ;
 assign wire1595 = ( wire132 ) | ( wire46 ) | ( wire280 ) | ( wire121 ) ;
 assign n_n54 = ( i_9_  &  i_10_  &  (~ i_11_)  &  wire728 ) ;
 assign n_n52 = ( (~ i_9_)  &  i_10_  &  (~ i_11_)  &  wire728 ) ;
 assign n_n519 = ( n_n39  &  n_n54 ) | ( n_n38  &  n_n52 ) | ( n_n39  &  n_n52 ) ;
 assign n_n4597 = ( n_n38  &  n_n134 ) | ( n_n38  &  n_n132 ) | ( n_n39  &  n_n132 ) ;
 assign n_n156 = ( i_9_  &  i_10_  &  (~ i_11_) ) ;
 assign n_n205 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_ ) ;
 assign n_n211 = ( i_14_  &  (~ i_13_)  &  (~ i_12_) ) ;
 assign wire390 = ( n_n39  &  n_n54 ) | ( n_n38  &  n_n52 ) ;
 assign n_n177 = ( i_9_  &  (~ i_10_)  &  i_11_ ) ;
 assign wire719 = ( i_14_  &  i_13_  &  i_12_  &  i_15_ ) ;
 assign wire393 = ( n_n38  &  n_n177  &  wire719 ) ;
 assign wire712 = ( n_n38  &  n_n54 ) | ( n_n39  &  n_n52 ) ;
 assign wire714 = ( i_8_  &  (~ i_1_)  &  (~ i_2_)  &  (~ i_0_) ) ;
 assign n_n31 = ( (~ i_7_)  &  (~ i_6_)  &  n_n162  &  wire714 ) ;
 assign n_n30 = ( n_n162  &  n_n35  &  n_n220 ) ;
 assign wire143 = ( wire717  &  n_n216 ) | ( n_n216  &  wire716 ) | ( n_n216  &  wire718 ) ;
 assign wire154 = ( wire723  &  n_n216 ) | ( wire730  &  n_n216 ) | ( wire727  &  n_n216 ) ;
 assign wire47 = ( wire720  &  n_n216 ) | ( wire722  &  n_n216 ) | ( wire715  &  n_n216 ) ;
 assign n_n4161 = ( n_n30  &  wire143 ) | ( n_n30  &  wire154 ) | ( n_n30  &  wire47 ) ;
 assign n_n170 = ( (~ i_9_)  &  (~ i_10_)  &  i_11_ ) ;
 assign wire720 = ( i_14_  &  (~ i_13_)  &  i_12_  &  i_15_ ) ;
 assign wire722 = ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  i_15_ ) ;
 assign wire715 = ( i_14_  &  i_13_  &  (~ i_12_)  &  i_15_ ) ;
 assign wire132 = ( n_n170  &  wire720 ) | ( n_n170  &  wire722 ) | ( n_n170  &  wire715 ) ;
 assign wire723 = ( i_14_  &  i_13_  &  (~ i_12_)  &  (~ i_15_) ) ;
 assign wire730 = ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  (~ i_15_) ) ;
 assign wire727 = ( i_14_  &  i_13_  &  i_12_  &  (~ i_15_) ) ;
 assign wire137 = ( n_n177  &  wire723 ) | ( n_n177  &  wire730 ) | ( n_n177  &  wire727 ) ;
 assign n_n4449 = ( n_n31  &  wire168 ) | ( n_n31  &  wire74 ) | ( n_n31  &  wire68 ) ;
 assign wire1864 = ( wire168 ) | ( wire74 ) | ( wire68 ) | ( wire151 ) ;
 assign wire17164 = ( n_n31  &  wire181 ) | ( n_n31  &  wire151 ) ;
 assign wire599 = ( n_n4449 ) | ( wire17164 ) | ( n_n30  &  wire1864 ) ;
 assign wire146 = ( n_n177  &  wire717 ) | ( n_n177  &  wire716 ) | ( n_n177  &  wire718 ) ;
 assign wire131 = ( wire729  &  n_n177 ) | ( n_n177  &  wire726 ) | ( n_n177  &  wire724 ) ;
 assign wire695 = ( n_n31  &  wire146 ) | ( n_n31  &  wire131 ) ;
 assign wire17198 = ( wire17196 ) | ( _5193 ) | ( wire176  &  _29653 ) ;
 assign wire17213 = ( wire4671 ) | ( wire17203 ) | ( wire17206 ) | ( wire17212 ) ;
 assign n_n2239 = ( wire4658 ) | ( wire4659 ) | ( wire17217 ) ;
 assign wire4643 = ( n_n162  &  n_n35  &  n_n220  &  wire899 ) ;
 assign wire17249 = ( wire4639 ) | ( wire17241 ) | ( wire17246 ) | ( wire17247 ) ;
 assign wire17256 = ( n_n71  &  n_n125 ) | ( n_n125  &  wire115 ) | ( n_n125  &  wire17253 ) ;
 assign wire17257 = ( wire17251 ) | ( n_n123  &  wire971 ) | ( n_n123  &  wire1176 ) ;
 assign wire4561 = ( wire243  &  wire979 ) | ( wire729  &  n_n199  &  wire979 ) ;
 assign wire4562 = ( n_n34  &  wire164 ) | ( n_n34  &  wire358 ) ;
 assign wire17303 = ( wire4568 ) | ( wire4569 ) | ( wire17299 ) | ( wire17301 ) ;
 assign wire17305 = ( wire17289 ) | ( wire17290 ) | ( wire17297 ) | ( wire17298 ) ;
 assign wire17322 = ( wire4545 ) | ( wire4548 ) | ( wire4549 ) ;
 assign n_n2249 = ( n_n2310 ) | ( wire17333 ) | ( wire4526 ) | ( _4924 ) ;
 assign wire17341 = ( n_n41  &  wire51 ) | ( n_n41  &  wire202 ) | ( n_n41  &  wire17339 ) ;
 assign wire17342 = ( wire4520 ) | ( wire17338 ) | ( n_n40  &  wire1794 ) ;
 assign n_n2265 = ( wire4485 ) | ( wire4486 ) | ( wire17367 ) | ( wire17368 ) ;
 assign n_n2266 = ( wire4481 ) | ( wire17374 ) | ( n_n212  &  wire1049 ) ;
 assign wire17379 = ( wire4474 ) | ( wire4475 ) | ( wire17377 ) ;
 assign n_n2234 = ( n_n2265 ) | ( n_n2266 ) | ( wire17379 ) ;
 assign n_n4120 = ( n_n4161 ) | ( wire449 ) | ( wire656 ) | ( wire17410 ) ;
 assign wire4434 = ( _4492 ) | ( n_n33  &  wire234 ) | ( n_n33  &  wire84 ) ;
 assign wire17420 = ( wire443 ) | ( wire17417 ) | ( wire17418 ) ;
 assign n_n4106 = ( wire599 ) | ( n_n4120 ) | ( wire4434 ) | ( wire17420 ) ;
 assign n_n19 = ( (~ i_1_)  &  i_2_  &  i_0_ ) ;
 assign n_n111 = ( (~ i_5_)  &  (~ i_3_)  &  (~ i_4_) ) ;
 assign n_n7241 = ( (~ i_7_)  &  (~ i_6_)  &  n_n19  &  n_n111 ) ;
 assign n_n7240 = ( (~ i_7_)  &  i_6_  &  n_n19  &  n_n111 ) ;
 assign n_n51 = ( (~ i_9_)  &  i_10_  &  (~ i_11_)  &  wire725 ) ;
 assign wire747 = ( (~ i_7_)  &  i_8_  &  (~ i_6_) ) ;
 assign n_n13 = ( n_n159  &  n_n111  &  wire747 ) ;
 assign wire717 = ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  i_15_ ) ;
 assign n_n149 = ( (~ i_9_)  &  i_10_  &  (~ i_11_) ) ;
 assign wire77 = ( wire730  &  n_n149 ) | ( wire717  &  n_n149 ) ;
 assign wire431 = ( i_7_  &  i_6_  &  n_n19  &  n_n111 ) | ( i_7_  &  (~ i_6_)  &  n_n19  &  n_n111 ) ;
 assign wire529 = ( i_7_  &  (~ i_6_)  &  n_n159  &  n_n111 ) ;
 assign wire568 = ( i_7_  &  i_6_  &  n_n219  &  n_n111 ) | ( i_7_  &  (~ i_6_)  &  n_n219  &  n_n111 ) ;
 assign wire569 = ( (~ i_7_)  &  i_6_  &  n_n219  &  n_n111 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n219  &  n_n111 ) ;
 assign n_n53 = ( i_9_  &  i_10_  &  (~ i_11_)  &  wire725 ) ;
 assign n_n3825 = ( n_n3578 ) | ( wire4067 ) | ( wire17716 ) | ( wire17717 ) ;
 assign wire4060 = ( _4048 ) | ( wire241  &  n_n112 ) | ( wire273  &  n_n112 ) ;
 assign wire17726 = ( wire515 ) | ( wire4064 ) | ( wire4065 ) | ( wire17725 ) ;
 assign wire17729 = ( n_n101  &  wire181 ) | ( n_n101  &  wire1378 ) | ( n_n108  &  wire1378 ) ;
 assign n_n3795 = ( n_n3825 ) | ( wire4060 ) | ( wire17726 ) | ( wire17729 ) ;
 assign n_n3800 = ( wire449 ) | ( wire656 ) | ( wire3985 ) | ( wire17787 ) ;
 assign n_n3802 = ( n_n3514 ) | ( wire17793 ) | ( n_n30  &  wire1491 ) ;
 assign wire17798 = ( n_n3511 ) | ( wire3973 ) | ( wire17796 ) ;
 assign n_n3787 = ( n_n3800 ) | ( n_n3802 ) | ( wire17798 ) ;
 assign wire17831 = ( n_n36  &  wire52 ) | ( n_n36  &  wire129 ) ;
 assign wire17832 = ( wire146  &  n_n34 ) | ( wire131  &  n_n34 ) ;
 assign wire17836 = ( n_n3525 ) | ( wire17822 ) | ( n_n34  &  wire129 ) ;
 assign wire17839 = ( wire17825 ) | ( wire17826 ) | ( wire17830 ) | ( wire17837 ) ;
 assign wire721 = ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  i_15_ ) ;
 assign wire728 = ( i_14_  &  (~ i_13_)  &  i_12_  &  (~ i_15_) ) ;
 assign wire157 = ( n_n156  &  wire719 ) | ( n_n156  &  wire721 ) | ( n_n156  &  wire728 ) ;
 assign n_n157 = ( (~ i_7_)  &  (~ i_6_) ) ;
 assign wire213 = ( i_8_  &  n_n162  &  n_n220  &  n_n157 ) | ( (~ i_8_)  &  n_n162  &  n_n220  &  n_n157 ) ;
 assign n_n36 = ( (~ i_7_)  &  (~ i_6_)  &  n_n218  &  wire714 ) ;
 assign n_n34 = ( n_n218  &  n_n35  &  n_n220 ) ;
 assign wire597 = ( wire432 ) | ( wire17034 ) | ( wire17035 ) ;
 assign wire620 = ( n_n4460 ) | ( wire17033 ) ;
 assign n_n2630 = ( wire17880 ) | ( wire17881 ) | ( n_n34  &  wire1627 ) ;
 assign wire17884 = ( wire642 ) | ( wire17028 ) | ( _30623 ) ;
 assign n_n2622 = ( wire597 ) | ( wire620 ) | ( n_n2630 ) | ( wire17884 ) ;
 assign n_n3467 = ( wire449 ) | ( wire656 ) | ( wire3820 ) | ( wire17926 ) ;
 assign wire17934 = ( n_n3510 ) | ( n_n31  &  wire1625 ) ;
 assign wire17935 = ( n_n4449 ) | ( n_n3514 ) | ( n_n3511 ) | ( wire17931 ) ;
 assign n_n3454 = ( n_n3467 ) | ( wire17934 ) | ( wire17935 ) ;
 assign n_n3473 = ( wire458 ) | ( n_n3525 ) | ( wire584 ) | ( wire17960 ) ;
 assign wire17958 = ( _30824 ) | ( wire154  &  n_n36 ) | ( wire47  &  n_n36 ) ;
 assign wire17959 = ( n_n4460 ) | ( wire17955 ) | ( n_n36  &  wire151 ) ;
 assign wire17968 = ( wire642 ) | ( wire17963 ) | ( wire17964 ) | ( wire17965 ) ;
 assign n_n3456 = ( n_n3473 ) | ( wire17958 ) | ( wire17959 ) | ( wire17968 ) ;
 assign n_n7263 = ( (~ i_7_)  &  (~ i_6_)  &  n_n219  &  n_n48 ) ;
 assign n_n161 = ( i_7_  &  (~ i_8_)  &  i_6_ ) ;
 assign n_n7265 = ( i_7_  &  (~ i_6_)  &  n_n219  &  n_n218 ) ;
 assign n_n7267 = ( (~ i_7_)  &  (~ i_6_)  &  n_n219  &  n_n218 ) ;
 assign wire3628 = ( n_n10  &  wire253 ) | ( wire253  &  n_n12 ) ;
 assign wire3629 = ( n_n9  &  n_n151 ) | ( n_n6  &  n_n151 ) | ( n_n151  &  n_n12 ) ;
 assign wire18150 = ( n_n9  &  wire717  &  n_n149 ) | ( n_n9  &  wire717  &  n_n191 ) ;
 assign wire253 = ( (~ i_9_)  &  i_10_  &  (~ i_11_)  &  wire717 ) | ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire717 ) ;
 assign n_n4308 = ( n_n48  &  n_n220  &  wire157  &  n_n161 ) ;
 assign n_n6271 = ( n_n124  &  n_n220  &  n_n177  &  n_n111 ) ;
 assign n_n126 = ( (~ i_7_)  &  i_8_  &  i_6_ ) ;
 assign n_n6267 = ( n_n220  &  n_n156  &  n_n111  &  n_n126 ) ;
 assign n_n47 = ( i_7_  &  i_6_  &  n_n48  &  wire714 ) ;
 assign wire152 = ( wire725  &  n_n149 ) | ( n_n149  &  wire721 ) | ( n_n149  &  wire728 ) ;
 assign wire4260 = ( n_n46  &  wire173 ) | ( n_n46  &  wire204 ) ;
 assign wire17554 = ( n_n47  &  _30153 ) | ( wire719  &  n_n47  &  _30155 ) ;
 assign n_n3085 = ( wire4260 ) | ( wire17554 ) | ( n_n47  &  wire152 ) ;
 assign n_n6266 = ( n_n220  &  n_n177  &  n_n111  &  n_n126 ) ;
 assign n_n6270 = ( n_n220  &  n_n170  &  n_n111  &  n_n126 ) ;
 assign n_n6269 = ( n_n124  &  n_n220  &  n_n111  &  n_n149 ) ;
 assign n_n6268 = ( n_n124  &  n_n220  &  n_n170  &  n_n111 ) ;
 assign wire245 = ( wire719  &  n_n149 ) | ( n_n149  &  wire721 ) | ( n_n149  &  wire728 ) ;
 assign n_n5052 = ( n_n17  &  n_n48  &  wire714  &  wire245 ) ;
 assign n_n41 = ( i_7_  &  (~ i_6_)  &  n_n48  &  wire714 ) ;
 assign n_n40 = ( n_n48  &  n_n220  &  n_n200 ) ;
 assign n_n57 = ( i_9_  &  (~ i_10_)  &  i_11_  &  wire725 ) ;
 assign wire144 = ( n_n156  &  wire719 ) | ( n_n156  &  wire728 ) ;
 assign n_n5055 = ( n_n40  &  n_n57 ) | ( n_n41  &  wire144 ) ;
 assign wire122 = ( wire725  &  n_n156 ) | ( n_n156  &  wire721 ) ;
 assign wire3469 = ( wire152  &  n_n40 ) | ( wire719  &  n_n149  &  n_n40 ) ;
 assign wire751 = ( n_n159  &  n_n218  &  n_n126 ) ;
 assign wire18298 = ( n_n159  &  n_n218  &  wire747 ) ;
 assign wire525 = ( wire725  &  n_n149  &  wire751 ) | ( wire725  &  n_n149  &  wire18298 ) ;
 assign n_n200 = ( i_7_  &  (~ i_8_)  &  (~ i_6_) ) ;
 assign n_n33 = ( n_n162  &  n_n220  &  n_n200 ) ;
 assign wire1417 = ( n_n184  &  wire725 ) | ( n_n184  &  wire719 ) | ( n_n184  &  wire728 ) ;
 assign wire55 = ( wire720  &  n_n149 ) | ( wire722  &  n_n149 ) | ( wire715  &  n_n149 ) ;
 assign wire149 = ( wire729  &  n_n170 ) | ( n_n170  &  wire726 ) | ( n_n170  &  wire724 ) ;
 assign wire127 = ( wire723  &  n_n149 ) | ( wire730  &  n_n149 ) | ( wire727  &  n_n149 ) ;
 assign n_n2728 = ( n_n33  &  wire55 ) | ( n_n33  &  wire149 ) | ( n_n33  &  wire127 ) ;
 assign wire675 = ( n_n33  &  wire150 ) | ( n_n33  &  wire129 ) ;
 assign wire3451 = ( n_n33  &  wire63 ) | ( n_n33  &  wire52 ) ;
 assign wire18301 = ( n_n33  &  wire48 ) | ( n_n33  &  n_n128 ) | ( n_n33  &  wire173 ) ;
 assign wire18302 = ( wire130  &  n_n32 ) | ( wire139  &  n_n32 ) | ( n_n32  &  wire128 ) ;
 assign wire126 = ( n_n170  &  wire723 ) | ( n_n170  &  wire730 ) | ( n_n170  &  wire727 ) ;
 assign wire587 = ( wire132  &  n_n33 ) | ( n_n33  &  wire126 ) ;
 assign wire172 = ( wire725  &  n_n191 ) | ( wire721  &  n_n191 ) | ( wire728  &  n_n191 ) ;
 assign wire147 = ( n_n170  &  wire717 ) | ( n_n170  &  wire716 ) | ( n_n170  &  wire718 ) ;
 assign wire158 = ( wire729  &  n_n149 ) | ( n_n149  &  wire726 ) | ( n_n149  &  wire724 ) ;
 assign wire133 = ( wire717  &  n_n149 ) | ( n_n149  &  wire716 ) | ( n_n149  &  wire718 ) ;
 assign wire767 = ( wire172 ) | ( wire147 ) | ( wire158 ) | ( wire133 ) ;
 assign n_n6 = ( n_n159  &  n_n35  &  n_n48 ) ;
 assign n_n3389 = ( i_7_  &  i_6_  &  n_n219  &  n_n111 ) | ( (~ i_7_)  &  i_6_  &  n_n219  &  n_n111 ) | ( i_7_  &  (~ i_6_)  &  n_n219  &  n_n111 ) ;
 assign n_n191 = ( i_9_  &  (~ i_10_)  &  (~ i_11_) ) ;
 assign wire145 = ( wire729  &  n_n191 ) | ( wire730  &  n_n191 ) ;
 assign wire388 = ( (~ i_7_)  &  i_6_  &  n_n162  &  n_n219 ) | ( i_7_  &  (~ i_6_)  &  n_n162  &  n_n219 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n162  &  n_n219 ) ;
 assign wire770 = ( wire729  &  n_n156 ) | ( n_n156  &  wire730 ) | ( n_n156  &  wire717 ) ;
 assign n_n3179 = ( wire3469 ) | ( wire3470 ) | ( wire18360 ) | ( wire18361 ) ;
 assign wire18375 = ( wire3550 ) | ( wire3551 ) | ( wire18370 ) | ( wire18371 ) ;
 assign n_n144 = ( (~ i_9_)  &  i_10_  &  (~ i_11_)  &  wire717 ) ;
 assign n_n7346 = ( i_7_  &  i_6_  &  n_n159  &  n_n218 ) ;
 assign n_n3 = ( n_n159  &  n_n218  &  n_n124 ) ;
 assign n_n2 = ( n_n159  &  n_n218  &  n_n35 ) ;
 assign wire430 = ( i_7_  &  (~ i_6_)  &  n_n159  &  n_n218 ) ;
 assign wire708 = ( wire430 ) | ( wire77  &  n_n2 ) ;
 assign n_n18 = ( i_7_  &  i_6_ ) ;
 assign n_n5319 = ( (~ i_7_)  &  (~ i_6_)  &  n_n159  &  _31153 ) ;
 assign wire17587 = ( i_7_  &  (~ i_5_)  &  i_6_ ) ;
 assign wire684 = ( i_3_  &  i_4_  &  n_n159  &  wire17587 ) ;
 assign n_n197 = ( n_n218  &  n_n220  &  n_n200 ) ;
 assign n_n212 = ( i_7_  &  (~ i_6_)  &  n_n218  &  wire714 ) ;
 assign n_n4441 = ( n_n4518 ) | ( wire17100 ) | ( n_n197  &  wire1224 ) ;
 assign wire575 = ( wire4739 ) | ( wire4740 ) | ( wire17102 ) ;
 assign wire18577 = ( n_n2777 ) | ( wire18575 ) ;
 assign wire18578 = ( wire18576 ) | ( n_n197  &  wire1602 ) ;
 assign n_n2754 = ( wire3177 ) | ( wire18581 ) | ( wire18582 ) | ( wire18583 ) ;
 assign wire18593 = ( wire594 ) | ( wire681 ) | ( wire504 ) | ( wire18586 ) ;
 assign wire18594 = ( n_n2770 ) | ( n_n3601 ) | ( wire18587 ) | ( wire18588 ) ;
 assign n_n2747 = ( n_n2754 ) | ( wire18593 ) | ( wire18594 ) ;
 assign n_n101 = ( n_n162  &  n_n124  &  n_n220 ) ;
 assign n_n42 = ( n_n162  &  n_n220  &  n_n161 ) ;
 assign wire3128 = ( n_n42  &  wire130 ) | ( n_n42  &  wire124 ) ;
 assign wire18624 = ( n_n42  &  wire139 ) | ( n_n43  &  wire139 ) ;
 assign wire18625 = ( n_n43  &  wire52 ) | ( n_n43  &  wire129 ) ;
 assign wire18626 = ( n_n43  &  wire124 ) | ( n_n42  &  wire128 ) | ( n_n43  &  wire128 ) ;
 assign n_n4755 = ( wire3128 ) | ( wire18624 ) | ( wire18625 ) | ( wire18626 ) ;
 assign wire381 = ( wire725  &  n_n156 ) | ( n_n156  &  wire721 ) | ( n_n156  &  wire728 ) ;
 assign n_n43 = ( i_7_  &  i_6_  &  n_n162  &  wire714 ) ;
 assign wire63 = ( wire723  &  n_n191 ) | ( wire730  &  n_n191 ) | ( wire727  &  n_n191 ) ;
 assign wire48 = ( wire720  &  n_n191 ) | ( wire722  &  n_n191 ) | ( wire715  &  n_n191 ) ;
 assign wire662 = ( n_n43  &  wire63 ) | ( n_n43  &  wire48 ) ;
 assign wire18711 = ( n_n5058 ) | ( wire3550 ) | ( wire3551 ) | ( wire4900 ) ;
 assign wire18712 = ( n_n5055 ) | ( wire18709 ) | ( n_n40  &  wire182 ) ;
 assign wire18719 = ( n_n3054 ) | ( wire18701 ) | ( wire18702 ) | ( wire18718 ) ;
 assign wire2977 = ( n_n162  &  n_n35  &  n_n220  &  wire1023 ) ;
 assign wire18783 = ( wire2979 ) | ( n_n31  &  wire1022 ) | ( n_n31  &  wire1263 ) ;
 assign wire18789 = ( wire18786 ) | ( _31572 ) | ( wire1096  &  _31567 ) ;
 assign wire18790 = ( wire18776 ) | ( wire18777 ) | ( wire18788 ) ;
 assign n_n6005 = ( n_n220  &  n_n111  &  n_n149  &  n_n200 ) ;
 assign wire17072 = ( i_7_  &  i_8_  &  (~ i_6_) ) ;
 assign wire419 = ( n_n220  &  n_n156  &  n_n111  &  wire17072 ) ;
 assign wire445 = ( n_n220  &  n_n177  &  n_n111  &  wire17072 ) ;
 assign wire446 = ( n_n220  &  n_n170  &  n_n111  &  n_n200 ) ;
 assign wire3470 = ( wire725  &  n_n156  &  _31049 ) | ( n_n156  &  wire721  &  _31049 ) ;
 assign wire18360 = ( n_n5055 ) | ( wire245  &  n_n41 ) | ( n_n41  &  wire150 ) ;
 assign wire18361 = ( n_n5059 ) | ( n_n5058 ) | ( wire18358 ) ;
 assign wire95 = ( n_n156  &  wire730 ) | ( n_n156  &  wire717 ) ;
 assign n_n799 = ( wire2329 ) | ( wire2331 ) | ( wire19480 ) | ( wire19481 ) ;
 assign wire2310 = ( n_n30  &  wire111 ) | ( n_n30  &  wire297 ) | ( n_n30  &  wire19500 ) ;
 assign wire19504 = ( wire2324 ) | ( wire19491 ) | ( wire19498 ) | ( wire19499 ) ;
 assign wire777 = ( i_9_  &  (~ i_10_)  &  i_11_  &  wire719 ) | ( i_9_  &  i_10_  &  (~ i_11_)  &  wire719 ) | ( (~ i_9_)  &  i_10_  &  (~ i_11_)  &  wire719 ) ;
 assign wire776 = ( i_9_  &  (~ i_10_)  &  i_11_  &  wire719 ) | ( i_9_  &  i_10_  &  (~ i_11_)  &  wire719 ) | ( (~ i_9_)  &  i_10_  &  (~ i_11_)  &  wire719 ) | ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire719 ) ;
 assign wire775 = ( (~ i_9_)  &  (~ i_10_)  &  i_11_  &  wire719 ) | ( (~ i_9_)  &  (~ i_10_)  &  (~ i_11_)  &  wire719 ) ;
 assign n_n7252 = ( i_7_  &  i_6_  &  n_n162  &  n_n219 ) ;
 assign wire389 = ( i_7_  &  i_6_  &  n_n162  &  n_n19 ) | ( (~ i_7_)  &  i_6_  &  n_n162  &  n_n19 ) | ( i_7_  &  (~ i_6_)  &  n_n162  &  n_n19 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n162  &  n_n19 ) ;
 assign wire3248 = ( i_7_  &  i_6_  &  n_n159  &  n_n111 ) ;
 assign wire454 = ( wire3248 ) | ( n_n5  &  wire77 ) ;
 assign wire742 = ( n_n159  &  n_n111  &  n_n126 ) ;
 assign wire779 = ( (~ i_9_)  &  i_10_  &  (~ i_11_)  &  wire725 ) | ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire725 ) | ( (~ i_9_)  &  (~ i_10_)  &  (~ i_11_)  &  wire725 ) ;
 assign wire783 = ( n_n159  &  n_n111  &  wire747 ) | ( n_n159  &  n_n111  &  n_n126 ) ;
 assign wire781 = ( (~ i_9_)  &  i_10_  &  (~ i_11_)  &  wire725 ) | ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire725 ) ;
 assign wire707 = ( wire430 ) | ( wire185  &  n_n2 ) ;
 assign n_n46 = ( n_n48  &  n_n220  &  n_n161 ) ;
 assign n_n199 = ( (~ i_9_)  &  i_10_  &  i_11_ ) ;
 assign wire726 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  (~ i_15_) ) ;
 assign wire724 = ( (~ i_14_)  &  i_13_  &  i_12_  &  (~ i_15_) ) ;
 assign wire168 = ( wire729  &  n_n199 ) | ( n_n199  &  wire726 ) | ( n_n199  &  wire724 ) ;
 assign n_n138 = ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire719 ) ;
 assign n_n216 = ( i_9_  &  i_10_  &  i_11_ ) ;
 assign wire214 = ( wire725  &  n_n216 ) | ( wire721  &  n_n216 ) ;
 assign n_n5107 = ( n_n47  &  n_n138 ) | ( n_n46  &  wire214 ) ;
 assign n_n108 = ( n_n162  &  n_n220  &  n_n126 ) ;
 assign n_n148 = ( (~ i_9_)  &  i_10_  &  (~ i_11_)  &  wire720 ) ;
 assign wire90 = ( wire729  &  n_n156 ) | ( n_n156  &  wire726 ) ;
 assign n_n5000 = ( n_n101  &  n_n148 ) | ( n_n108  &  wire90 ) ;
 assign wire98 = ( wire720  &  n_n191 ) | ( wire715  &  n_n191 ) ;
 assign n_n102 = ( i_9_  &  i_10_  &  i_11_  &  wire729 ) ;
 assign n_n1434 = ( n_n31  &  wire98 ) | ( n_n30  &  n_n102 ) ;
 assign wire118 = ( wire720  &  n_n149 ) | ( wire715  &  n_n149 ) ;
 assign n_n1408 = ( n_n71  &  n_n31 ) | ( n_n30  &  wire118 ) ;
 assign wire120 = ( n_n177  &  wire717 ) | ( n_n177  &  wire726 ) | ( n_n177  &  wire724 ) ;
 assign wire179 = ( n_n177  &  wire730 ) | ( n_n177  &  wire716 ) | ( n_n177  &  wire718 ) ;
 assign wire324 = ( n_n177  &  wire722 ) | ( n_n177  &  wire723 ) | ( n_n177  &  wire727 ) ;
 assign wire18720 = ( wire729  &  n_n177 ) | ( n_n177  &  wire720 ) | ( n_n177  &  wire715 ) ;
 assign wire789 = ( wire120 ) | ( wire179 ) | ( wire324 ) | ( wire18720 ) ;
 assign n_n117 = ( (~ i_9_)  &  (~ i_10_)  &  (~ i_11_)  &  wire729 ) ;
 assign n_n1426 = ( n_n30  &  wire98 ) | ( n_n31  &  n_n117 ) ;
 assign n_n89 = ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire729 ) ;
 assign wire93 = ( wire717  &  n_n191 ) | ( n_n191  &  wire726 ) | ( n_n191  &  wire724 ) ;
 assign wire241 = ( wire730  &  n_n191 ) | ( n_n191  &  wire716 ) | ( n_n191  &  wire718 ) ;
 assign wire273 = ( wire722  &  n_n191 ) | ( wire723  &  n_n191 ) | ( wire727  &  n_n191 ) ;
 assign wire791 = ( n_n89 ) | ( wire93 ) | ( wire241 ) | ( wire273 ) ;
 assign wire53 = ( n_n170  &  wire720 ) | ( n_n170  &  wire715 ) ;
 assign n_n77 = ( (~ i_9_)  &  (~ i_10_)  &  i_11_  &  wire729 ) ;
 assign n_n1416 = ( n_n31  &  wire53 ) | ( n_n30  &  n_n77 ) ;
 assign wire117 = ( n_n170  &  wire717 ) | ( n_n170  &  wire726 ) | ( n_n170  &  wire724 ) ;
 assign wire281 = ( n_n170  &  wire730 ) | ( n_n170  &  wire716 ) | ( n_n170  &  wire718 ) ;
 assign wire294 = ( n_n170  &  wire722 ) | ( n_n170  &  wire723 ) | ( n_n170  &  wire727 ) ;
 assign wire793 = ( wire53 ) | ( wire117 ) | ( wire281 ) | ( wire294 ) ;
 assign n_n125 = ( n_n218  &  n_n220  &  n_n126 ) ;
 assign wire85 = ( wire722  &  n_n216 ) | ( wire715  &  n_n216 ) | ( wire727  &  n_n216 ) ;
 assign wire142 = ( wire723  &  n_n216 ) | ( wire730  &  n_n216 ) | ( n_n216  &  wire716 ) ;
 assign wire422 = ( n_n125  &  wire85 ) | ( n_n125  &  wire142 ) ;
 assign wire150 = ( wire725  &  n_n170 ) | ( n_n170  &  wire721 ) | ( n_n170  &  wire728 ) ;
 assign wire80 = ( n_n177  &  wire719 ) | ( n_n177  &  wire728 ) ;
 assign wire78 = ( wire725  &  n_n177 ) | ( n_n177  &  wire721 ) ;
 assign n_n55 = ( (~ i_9_)  &  (~ i_10_)  &  i_11_  &  wire725 ) ;
 assign wire252 = ( wire719  &  n_n170 ) | ( n_n170  &  wire721 ) | ( n_n170  &  wire728 ) ;
 assign wire796 = ( wire80 ) | ( wire78 ) | ( n_n55 ) | ( wire252 ) ;
 assign wire207 = ( wire720  &  n_n149 ) | ( wire727  &  n_n149 ) ;
 assign n_n150 = ( i_9_  &  i_10_  &  (~ i_11_)  &  wire726 ) ;
 assign n_n1520 = ( n_n38  &  wire207 ) | ( n_n39  &  n_n150 ) ;
 assign wire155 = ( n_n156  &  wire723 ) | ( n_n156  &  wire730 ) | ( n_n156  &  wire716 ) ;
 assign wire205 = ( n_n156  &  wire717 ) | ( n_n156  &  wire724 ) | ( n_n156  &  wire718 ) ;
 assign wire215 = ( n_n156  &  wire722 ) | ( n_n156  &  wire715 ) | ( n_n156  &  wire727 ) ;
 assign wire17490 = ( wire729  &  n_n156 ) | ( n_n156  &  wire720 ) | ( n_n156  &  wire726 ) ;
 assign wire800 = ( wire155 ) | ( wire205 ) | ( wire215 ) | ( wire17490 ) ;
 assign wire234 = ( wire723  &  n_n149 ) | ( wire730  &  n_n149 ) | ( n_n149  &  wire716 ) ;
 assign wire86 = ( wire729  &  n_n216 ) | ( wire726  &  n_n216 ) ;
 assign wire84 = ( wire722  &  n_n149 ) | ( wire715  &  n_n149 ) | ( wire727  &  n_n149 ) ;
 assign wire799 = ( n_n148 ) | ( wire234 ) | ( wire86 ) | ( wire84 ) ;
 assign wire181 = ( wire729  &  n_n216 ) | ( wire726  &  n_n216 ) | ( wire724  &  n_n216 ) ;
 assign wire134 = ( n_n156  &  wire720 ) | ( n_n156  &  wire722 ) | ( n_n156  &  wire715 ) ;
 assign wire156 = ( n_n156  &  wire723 ) | ( n_n156  &  wire730 ) | ( n_n156  &  wire727 ) ;
 assign wire458 = ( n_n36  &  wire134 ) | ( n_n36  &  wire156 ) ;
 assign wire176 = ( wire729  &  n_n156 ) | ( n_n156  &  wire726 ) | ( n_n156  &  wire724 ) ;
 assign wire123 = ( n_n156  &  wire717 ) | ( n_n156  &  wire716 ) | ( n_n156  &  wire718 ) ;
 assign wire541 = ( n_n36  &  wire176 ) | ( n_n36  &  wire123 ) ;
 assign wire4393 = ( wire90  &  n_n123 ) | ( wire155  &  n_n123 ) | ( wire205  &  n_n123 ) ;
 assign n_n3912 = ( wire4393 ) | ( wire719  &  n_n216  &  n_n125 ) ;
 assign n_n123 = ( n_n218  &  n_n124  &  n_n220 ) ;
 assign wire570 = ( wire90  &  n_n125 ) | ( n_n125  &  wire205 ) ;
 assign wire60 = ( wire729  &  n_n149 ) | ( n_n149  &  wire726 ) ;
 assign n_n1700 = ( n_n148  &  n_n125 ) | ( n_n123  &  wire60 ) ;
 assign wire220 = ( wire717  &  n_n149 ) | ( n_n149  &  wire724 ) | ( n_n149  &  wire718 ) ;
 assign wire803 = ( wire234 ) | ( wire84 ) | ( wire60 ) | ( wire220 ) ;
 assign wire17470 = ( n_n53  &  n_n108 ) | ( n_n101  &  wire218 ) ;
 assign wire17471 = ( wire157  &  n_n108 ) | ( n_n101  &  wire141 ) ;
 assign wire4829 = ( n_n47  &  wire142 ) | ( n_n47  &  wire86 ) | ( n_n47  &  wire180 ) ;
 assign n_n214 = ( i_9_  &  i_10_  &  i_11_  &  wire720 ) ;
 assign wire4354 = ( n_n220  &  n_n156  &  n_n111  &  n_n200 ) ;
 assign wire4355 = ( n_n220  &  n_n111  &  n_n149  &  wire17072 ) ;
 assign n_n1624 = ( wire4354 ) | ( wire4355 ) | ( n_n47  &  n_n214 ) ;
 assign wire17479 = ( n_n4996 ) | ( n_n4994 ) | ( n_n101  &  wire946 ) ;
 assign wire17486 = ( wire4343 ) | ( wire17484 ) | ( _4718 ) | ( _30071 ) ;
 assign n_n4112 = ( wire17486 ) | ( _30039 ) | ( _30040 ) | ( _30073 ) ;
 assign n_n155 = ( i_9_  &  i_10_  &  (~ i_11_)  &  wire720 ) ;
 assign n_n1594 = ( n_n47  &  wire60 ) | ( n_n46  &  n_n155 ) ;
 assign wire17082 = ( n_n4641 ) | ( n_n47  &  wire1840 ) ;
 assign wire808 = ( n_n148 ) | ( wire234 ) | ( wire84 ) | ( wire220 ) ;
 assign wire180 = ( wire717  &  n_n216 ) | ( wire724  &  n_n216 ) | ( n_n216  &  wire718 ) ;
 assign n_n4904 = ( n_n108  &  wire85 ) | ( n_n108  &  wire142 ) | ( n_n108  &  wire180 ) ;
 assign wire447 = ( n_n220  &  n_n156  &  n_n111  &  n_n161 ) ;
 assign wire4320 = ( n_n220  &  n_n111  &  n_n149  &  wire16987 ) ;
 assign n_n5037 = ( wire447 ) | ( wire4320 ) | ( n_n108  &  n_n214 ) ;
 assign n_n5033 = ( n_n108  &  wire86 ) | ( n_n101  &  n_n198 ) ;
 assign wire219 = ( wire722  &  n_n199 ) | ( wire715  &  n_n199 ) | ( wire727  &  n_n199 ) ;
 assign wire108 = ( wire723  &  n_n199 ) | ( wire730  &  n_n199 ) | ( n_n199  &  wire716 ) ;
 assign n_n4903 = ( n_n5033 ) | ( n_n101  &  wire219 ) | ( n_n101  &  wire108 ) ;
 assign wire1844 = ( wire219 ) | ( wire108 ) | ( wire258 ) | ( wire16980 ) ;
 assign wire4935 = ( n_n101  &  n_n214 ) | ( n_n101  &  wire70 ) | ( n_n101  &  wire258 ) ;
 assign wire544 = ( wire4935 ) | ( n_n108  &  wire1844 ) ;
 assign wire17501 = ( wire17493 ) | ( wire17499 ) | ( _30087 ) ;
 assign wire716 = ( (~ i_14_)  &  i_13_  &  i_12_  &  i_15_ ) ;
 assign wire718 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  i_15_ ) ;
 assign wire52 = ( wire717  &  n_n191 ) | ( n_n191  &  wire716 ) | ( n_n191  &  wire718 ) ;
 assign wire129 = ( wire729  &  n_n191 ) | ( n_n191  &  wire726 ) | ( n_n191  &  wire724 ) ;
 assign n_n4622 = ( n_n17  &  n_n48  &  wire714  &  wire142 ) ;
 assign wire182 = ( n_n177  &  wire719 ) | ( n_n177  &  wire721 ) | ( n_n177  &  wire728 ) ;
 assign n_n5060 = ( n_n17  &  n_n48  &  wire714  &  wire182 ) ;
 assign n_n130 = ( i_9_  &  i_10_  &  (~ i_11_)  &  wire719 ) ;
 assign n_n3276 = ( (~ i_7_)  &  i_6_  &  n_n48  &  n_n19 ) | ( i_7_  &  (~ i_6_)  &  n_n48  &  n_n19 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n48  &  n_n19 ) ;
 assign n_n83 = ( i_9_  &  (~ i_10_)  &  i_11_  &  wire729 ) ;
 assign n_n6445 = ( wire729  &  n_n177  &  n_n41 ) ;
 assign n_n7242 = ( i_7_  &  i_6_  &  n_n48  &  n_n19 ) ;
 assign n_n68 = ( (~ i_9_)  &  i_10_  &  (~ i_11_)  &  wire730 ) ;
 assign wire344 = ( i_9_  &  i_10_  &  (~ i_11_)  &  wire730 ) | ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire730 ) ;
 assign wire462 = ( i_7_  &  i_6_  &  n_n218  &  n_n19 ) | ( i_7_  &  (~ i_6_)  &  n_n218  &  n_n19 ) ;
 assign wire817 = ( i_5_  &  (~ i_3_)  &  i_4_ ) | ( (~ i_5_)  &  (~ i_3_)  &  (~ i_4_) ) ;
 assign wire130 = ( n_n184  &  wire729 ) | ( n_n184  &  wire726 ) | ( n_n184  &  wire724 ) ;
 assign wire188 = ( i_8_  &  n_n17  &  n_n218  &  n_n220 ) | ( (~ i_8_)  &  n_n17  &  n_n218  &  n_n220 ) ;
 assign n_n59 = ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire725 ) ;
 assign wire226 = ( i_8_  &  n_n218  &  n_n220  &  n_n157 ) | ( (~ i_8_)  &  n_n218  &  n_n220  &  n_n157 ) ;
 assign wire820 = ( (~ i_9_)  &  i_10_  &  i_11_  &  wire725 ) | ( i_9_  &  (~ i_10_)  &  i_11_  &  wire725 ) | ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire725 ) ;
 assign wire4558 = ( n_n218  &  wire714  &  n_n157  &  wire820 ) ;
 assign wire17307 = ( wire725  &  n_n34  &  n_n191 ) | ( wire725  &  n_n34  &  n_n216 ) ;
 assign wire4554 = ( _4984 ) | ( n_n34  &  wire115 ) | ( n_n34  &  wire17310 ) ;
 assign wire17314 = ( n_n36  &  n_n63 ) | ( n_n36  &  wire115 ) | ( n_n36  &  wire17309 ) ;
 assign wire304 = ( i_15_  &  n_n184  &  n_n211 ) | ( (~ i_15_)  &  n_n184  &  n_n211 ) | ( i_15_  &  n_n184  &  n_n204 ) ;
 assign wire306 = ( i_15_  &  n_n211  &  n_n191 ) | ( (~ i_15_)  &  n_n211  &  n_n191 ) | ( i_15_  &  n_n191  &  n_n204 ) ;
 assign wire824 = ( wire129 ) | ( wire130 ) | ( wire304 ) | ( wire306 ) ;
 assign wire4701 = ( n_n47  &  wire304 ) | ( n_n47  &  wire306 ) | ( n_n47  &  wire200 ) ;
 assign wire17178 = ( n_n47  &  wire129 ) | ( n_n47  &  wire130 ) ;
 assign n_n2253 = ( wire4701 ) | ( wire17178 ) | ( n_n46  &  wire824 ) ;
 assign n_n61 = ( (~ i_9_)  &  i_10_  &  i_11_  &  wire725 ) ;
 assign wire228 = ( i_8_  &  n_n162  &  n_n16  &  n_n220 ) | ( (~ i_8_)  &  n_n162  &  n_n16  &  n_n220 ) ;
 assign n_n147 = ( (~ i_9_)  &  i_10_  &  (~ i_11_)  &  wire722 ) ;
 assign n_n63 = ( i_9_  &  i_10_  &  i_11_  &  wire725 ) ;
 assign wire351 = ( wire730  &  n_n149 ) | ( wire717  &  n_n149 ) | ( n_n149  &  wire724 ) ;
 assign wire377 = ( n_n156  &  wire730 ) | ( n_n156  &  wire717 ) | ( n_n156  &  wire724 ) ;
 assign wire139 = ( n_n184  &  wire717 ) | ( n_n184  &  wire716 ) | ( n_n184  &  wire718 ) ;
 assign n_n213 = ( i_14_  &  i_13_  &  (~ i_12_) ) ;
 assign wire257 = ( i_15_  &  n_n191  &  n_n213 ) | ( (~ i_15_)  &  n_n191  &  n_n213 ) ;
 assign wire313 = ( i_15_  &  n_n184  &  n_n213 ) | ( (~ i_15_)  &  n_n184  &  n_n213 ) ;
 assign n_n129 = ( i_9_  &  i_10_  &  (~ i_11_)  &  wire721 ) ;
 assign n_n166 = ( (~ i_9_)  &  (~ i_10_)  &  i_11_  &  wire716 ) ;
 assign n_n127 = ( (~ i_9_)  &  i_10_  &  (~ i_11_)  &  wire721 ) ;
 assign n_n82 = ( (~ i_9_)  &  (~ i_10_)  &  i_11_  &  wire715 ) ;
 assign wire190 = ( i_8_  &  n_n17  &  n_n48  &  n_n220 ) | ( (~ i_8_)  &  n_n17  &  n_n48  &  n_n220 ) ;
 assign wire334 = ( i_8_  &  n_n16  &  n_n48  &  n_n220 ) | ( (~ i_8_)  &  n_n16  &  n_n48  &  n_n220 ) ;
 assign wire836 = ( n_n177  &  wire715 ) | ( n_n170  &  wire715 ) | ( n_n177  &  wire716 ) ;
 assign n_n139 = ( (~ i_9_)  &  i_10_  &  i_11_  &  wire721 ) ;
 assign wire260 = ( n_n156  &  wire723 ) | ( n_n156  &  wire716 ) | ( n_n156  &  wire718 ) ;
 assign wire373 = ( wire729  &  n_n156 ) | ( n_n156  &  wire717 ) ;
 assign wire2900 = ( n_n40  &  wire345 ) | ( n_n156  &  wire715  &  n_n40 ) ;
 assign wire18865 = ( n_n36  &  n_n102 ) | ( n_n38  &  n_n73 ) ;
 assign wire18866 = ( n_n34  &  wire136 ) | ( n_n36  &  wire364 ) ;
 assign n_n1870 = ( wire18865 ) | ( wire18866 ) | ( wire143  &  n_n36 ) ;
 assign n_n95 = ( (~ i_9_)  &  i_10_  &  i_11_  &  wire729 ) ;
 assign wire74 = ( wire717  &  n_n199 ) | ( n_n199  &  wire716 ) | ( n_n199  &  wire718 ) ;
 assign wire136 = ( i_15_  &  n_n199  &  n_n213 ) | ( (~ i_15_)  &  n_n199  &  n_n213 ) ;
 assign wire840 = ( wire257 ) | ( n_n95 ) | ( wire74 ) | ( wire136 ) ;
 assign wire18857 = ( wire18854 ) | ( wire18855 ) | ( n_n39  &  wire836 ) ;
 assign wire18874 = ( n_n1870 ) | ( wire18871 ) | ( _2199 ) | ( _31940 ) ;
 assign n_n1800 = ( wire18874 ) | ( _31899 ) | ( _31900 ) | ( _31946 ) ;
 assign wire68 = ( wire723  &  n_n199 ) | ( wire730  &  n_n199 ) | ( wire727  &  n_n199 ) ;
 assign n_n112 = ( n_n218  &  n_n220  &  n_n161 ) ;
 assign n_n113 = ( i_7_  &  i_6_  &  n_n218  &  wire714 ) ;
 assign wire227 = ( n_n156  &  wire720 ) | ( n_n156  &  wire715 ) | ( n_n156  &  wire727 ) ;
 assign wire232 = ( i_15_  &  n_n156  &  n_n205 ) | ( (~ i_15_)  &  n_n156  &  n_n205 ) | ( i_15_  &  n_n156  &  n_n204 ) ;
 assign wire844 = ( wire127 ) | ( wire155 ) | ( wire227 ) | ( wire232 ) ;
 assign wire845 = ( wire721  &  n_n199 ) | ( wire728  &  n_n199 ) | ( wire721  &  n_n216 ) | ( wire728  &  n_n216 ) ;
 assign wire542 = ( n_n34  &  wire127 ) | ( n_n36  &  n_n148 ) ;
 assign wire850 = ( n_n149  &  wire721 ) | ( n_n149  &  wire728 ) ;
 assign wire849 = ( n_n156  &  wire721 ) | ( n_n149  &  wire721 ) | ( n_n156  &  wire728 ) | ( n_n149  &  wire728 ) ;
 assign n_n5109 = ( n_n65  &  n_n46 ) | ( n_n47  &  wire118 ) ;
 assign wire677 = ( n_n47  &  wire127 ) | ( n_n47  &  wire133 ) ;
 assign wire75 = ( wire717  &  n_n149 ) | ( n_n149  &  wire718 ) ;
 assign wire19119 = ( wire727  &  n_n149 ) | ( n_n149  &  wire726 ) ;
 assign wire852 = ( wire118 ) | ( wire234 ) | ( wire75 ) | ( wire19119 ) ;
 assign n_n140 = ( (~ i_9_)  &  i_10_  &  i_11_  &  wire719 ) ;
 assign n_n142 = ( i_9_  &  i_10_  &  i_11_  &  wire719 ) ;
 assign wire290 = ( n_n156  &  wire722 ) | ( n_n156  &  wire727 ) | ( n_n156  &  wire716 ) ;
 assign wire856 = ( wire290 ) | ( n_n156  &  wire720 ) | ( n_n156  &  wire715 ) ;
 assign n_n116 = ( (~ i_9_)  &  (~ i_10_)  &  (~ i_11_)  &  wire719 ) ;
 assign wire255 = ( i_8_  &  n_n16  &  n_n218  &  n_n220 ) | ( (~ i_8_)  &  n_n16  &  n_n218  &  n_n220 ) ;
 assign wire199 = ( wire722  &  n_n149 ) | ( wire727  &  n_n149 ) | ( n_n149  &  wire716 ) ;
 assign wire402 = ( wire719  &  n_n199 ) | ( n_n156  &  wire724 ) ;
 assign wire19640 = ( i_9_  &  i_10_  &  i_11_  &  wire719 ) | ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire719 ) ;
 assign wire19641 = ( wire720  &  n_n149 ) | ( wire715  &  n_n149 ) | ( n_n149  &  wire724 ) ;
 assign wire859 = ( wire199 ) | ( wire402 ) | ( wire19640 ) | ( wire19641 ) ;
 assign wire743 = ( (~ i_1_)  &  (~ i_2_)  &  i_0_  &  _30896 ) ;
 assign n_n103 = ( i_9_  &  i_10_  &  i_11_  &  wire724 ) ;
 assign n_n207 = ( (~ i_14_)  &  i_13_  &  i_12_ ) ;
 assign n_n173 = ( i_9_  &  (~ i_10_)  &  i_11_  &  wire716 ) ;
 assign n_n169 = ( (~ i_9_)  &  (~ i_10_)  &  i_11_  &  wire720 ) ;
 assign n_n204 = ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_) ) ;
 assign n_n151 = ( i_9_  &  i_10_  &  (~ i_11_)  &  wire717 ) ;
 assign n_n141 = ( i_9_  &  i_10_  &  i_11_  &  wire721 ) ;
 assign n_n115 = ( (~ i_9_)  &  (~ i_10_)  &  (~ i_11_)  &  wire721 ) ;
 assign n_n209 = ( i_14_  &  i_13_  &  i_12_ ) ;
 assign n_n178 = ( (~ i_9_)  &  (~ i_10_)  &  (~ i_11_)  &  wire726 ) ;
 assign n_n183 = ( (~ i_9_)  &  (~ i_10_)  &  (~ i_11_)  &  wire720 ) ;
 assign n_n90 = ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire724 ) ;
 assign n_n70 = ( (~ i_9_)  &  i_10_  &  (~ i_11_)  &  wire715 ) ;
 assign n_n62 = ( (~ i_9_)  &  i_10_  &  i_11_  &  wire728 ) ;
 assign n_n189 = ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire722 ) ;
 assign n_n122 = ( (~ i_9_)  &  (~ i_10_)  &  (~ i_11_)  &  wire715 ) ;
 assign n_n185 = ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire726 ) ;
 assign n_n84 = ( i_9_  &  (~ i_10_)  &  i_11_  &  wire724 ) ;
 assign n_n136 = ( (~ i_9_)  &  (~ i_10_)  &  (~ i_11_)  &  wire728 ) ;
 assign n_n210 = ( i_9_  &  i_10_  &  i_11_  &  wire722 ) ;
 assign n_n172 = ( i_9_  &  (~ i_10_)  &  i_11_  &  wire717 ) ;
 assign n_n58 = ( i_9_  &  (~ i_10_)  &  i_11_  &  wire728 ) ;
 assign n_n118 = ( (~ i_9_)  &  (~ i_10_)  &  (~ i_11_)  &  wire724 ) ;
 assign n_n32 = ( i_7_  &  (~ i_6_)  &  n_n162  &  wire714 ) ;
 assign n_n186 = ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire717 ) ;
 assign n_n107 = ( i_9_  &  i_10_  &  i_11_  &  wire715 ) ;
 assign n_n198 = ( (~ i_9_)  &  i_10_  &  i_11_  &  wire720 ) ;
 assign n_n168 = ( (~ i_9_)  &  (~ i_10_)  &  i_11_  &  wire722 ) ;
 assign n_n176 = ( i_9_  &  (~ i_10_)  &  i_11_  &  wire720 ) ;
 assign n_n60 = ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire728 ) ;
 assign n_n12 = ( n_n159  &  n_n124  &  n_n48 ) ;
 assign wire151 = ( wire720  &  n_n199 ) | ( wire722  &  n_n199 ) | ( wire715  &  n_n199 ) ;
 assign wire94 = ( n_n184  &  wire717 ) | ( n_n184  &  wire726 ) | ( n_n184  &  wire724 ) ;
 assign wire184 = ( n_n184  &  wire730 ) | ( n_n184  &  wire716 ) | ( n_n184  &  wire718 ) ;
 assign wire268 = ( n_n184  &  wire722 ) | ( n_n184  &  wire723 ) | ( n_n184  &  wire727 ) ;
 assign wire18738 = ( n_n184  &  wire729 ) | ( n_n184  &  wire720 ) | ( n_n184  &  wire715 ) ;
 assign wire860 = ( wire94 ) | ( wire184 ) | ( wire268 ) | ( wire18738 ) ;
 assign wire81 = ( wire720  &  n_n199 ) | ( wire715  &  n_n199 ) ;
 assign n_n1442 = ( n_n31  &  n_n102 ) | ( n_n30  &  wire81 ) ;
 assign wire111 = ( wire720  &  n_n216 ) | ( wire715  &  n_n216 ) ;
 assign wire162 = ( wire730  &  n_n216 ) | ( n_n216  &  wire716 ) | ( n_n216  &  wire718 ) ;
 assign wire164 = ( wire717  &  n_n216 ) | ( wire726  &  n_n216 ) | ( wire724  &  n_n216 ) ;
 assign wire341 = ( wire722  &  n_n216 ) | ( wire723  &  n_n216 ) | ( wire727  &  n_n216 ) ;
 assign wire863 = ( wire111 ) | ( wire162 ) | ( wire164 ) | ( wire341 ) ;
 assign wire206 = ( wire730  &  n_n199 ) | ( n_n199  &  wire716 ) | ( n_n199  &  wire718 ) ;
 assign wire243 = ( wire717  &  n_n199 ) | ( n_n199  &  wire726 ) | ( n_n199  &  wire724 ) ;
 assign wire368 = ( wire722  &  n_n199 ) | ( wire723  &  n_n199 ) | ( wire727  &  n_n199 ) ;
 assign wire18752 = ( wire729  &  n_n199 ) | ( wire720  &  n_n199 ) | ( wire715  &  n_n199 ) ;
 assign wire865 = ( wire206 ) | ( wire243 ) | ( wire368 ) | ( wire18752 ) ;
 assign wire153 = ( wire725  &  n_n199 ) | ( wire721  &  n_n199 ) ;
 assign n_n4686 = ( n_n212  &  n_n140 ) | ( n_n197  &  wire153 ) ;
 assign wire247 = ( wire725  &  n_n199 ) | ( wire721  &  n_n199 ) | ( wire728  &  n_n199 ) ;
 assign wire135 = ( wire719  &  n_n199 ) | ( wire728  &  n_n199 ) ;
 assign wire704 = ( n_n212  &  n_n63 ) | ( n_n197  &  wire135 ) ;
 assign n_n4231 = ( n_n4686 ) | ( wire704 ) | ( n_n212  &  wire247 ) ;
 assign wire218 = ( wire719  &  n_n199 ) | ( wire721  &  n_n199 ) | ( wire728  &  n_n199 ) ;
 assign wire248 = ( n_n156  &  wire723 ) | ( n_n156  &  wire730 ) | ( n_n156  &  wire718 ) ;
 assign n_n4460 = ( n_n36  &  wire168 ) | ( n_n36  &  wire74 ) | ( n_n36  &  wire68 ) ;
 assign n_n4900 = ( n_n101  &  wire85 ) | ( n_n101  &  wire142 ) | ( n_n101  &  wire180 ) ;
 assign wire867 = ( wire155 ) | ( wire205 ) | ( wire215 ) | ( n_n155 ) ;
 assign n_n4518 = ( wire143  &  n_n212 ) | ( wire154  &  n_n212 ) | ( wire47  &  n_n212 ) ;
 assign wire1224 = ( wire168 ) | ( wire74 ) | ( wire68 ) | ( wire151 ) ;
 assign wire17100 = ( n_n212  &  wire181 ) | ( n_n212  &  wire151 ) ;
 assign wire532 = ( wire127  &  n_n212 ) | ( wire133  &  n_n212 ) ;
 assign wire4739 = ( n_n212  &  wire74 ) | ( n_n212  &  wire68 ) ;
 assign wire4740 = ( wire143  &  n_n197 ) | ( wire154  &  n_n197 ) ;
 assign wire17102 = ( wire47  &  n_n197 ) | ( n_n212  &  wire168 ) ;
 assign wire594 = ( wire55  &  n_n197 ) | ( n_n212  &  wire176 ) ;
 assign wire660 = ( n_n212  &  wire134 ) | ( n_n212  &  wire156 ) ;
 assign wire17521 = ( wire17518 ) | ( wire158  &  n_n197 ) | ( wire133  &  n_n197 ) ;
 assign wire17522 = ( wire532 ) | ( wire594 ) | ( wire660 ) | ( wire17516 ) ;
 assign n_n4116 = ( n_n4441 ) | ( wire575 ) | ( wire17521 ) | ( wire17522 ) ;
 assign wire104 = ( n_n177  &  wire720 ) | ( n_n177  &  wire715 ) ;
 assign n_n5111 = ( n_n47  &  n_n77 ) | ( n_n46  &  wire104 ) ;
 assign n_n5113 = ( n_n46  &  n_n89 ) | ( n_n47  &  wire104 ) ;
 assign wire868 = ( wire98 ) | ( wire93 ) | ( wire241 ) | ( wire273 ) ;
 assign n_n7254 = ( (~ i_7_)  &  i_6_  &  n_n162  &  n_n219 ) ;
 assign n_n7248 = ( (~ i_7_)  &  i_6_  &  n_n218  &  n_n19 ) ;
 assign n_n3562 = ( n_n47  &  wire168 ) | ( n_n47  &  wire74 ) | ( n_n47  &  wire68 ) ;
 assign wire3601 = ( wire143  &  n_n46 ) | ( wire154  &  n_n46 ) ;
 assign wire18168 = ( n_n47  &  wire48 ) | ( n_n46  &  wire181 ) ;
 assign wire18169 = ( n_n47  &  wire63 ) | ( wire47  &  n_n46 ) ;
 assign n_n3398 = ( n_n3562 ) | ( wire3601 ) | ( wire18168 ) | ( wire18169 ) ;
 assign wire481 = ( wire154  &  n_n47 ) | ( wire47  &  n_n47 ) ;
 assign wire3594 = ( n_n46  &  wire74 ) | ( n_n46  &  wire68 ) ;
 assign wire18172 = ( n_n46  &  wire168 ) | ( n_n47  &  wire181 ) ;
 assign wire18173 = ( n_n47  &  wire151 ) | ( n_n46  &  wire151 ) ;
 assign wire18174 = ( wire143  &  n_n47 ) | ( wire154  &  n_n47 ) | ( wire47  &  n_n47 ) ;
 assign n_n3050 = ( wire3594 ) | ( wire18172 ) | ( wire18173 ) | ( wire18174 ) ;
 assign wire124 = ( n_n184  &  wire720 ) | ( n_n184  &  wire722 ) | ( n_n184  &  wire715 ) ;
 assign wire128 = ( n_n184  &  wire723 ) | ( n_n184  &  wire730 ) | ( n_n184  &  wire727 ) ;
 assign wire875 = ( wire130 ) | ( wire139 ) | ( wire124 ) | ( wire128 ) ;
 assign wire18180 = ( wire3588 ) | ( wire18178 ) | ( n_n46  &  wire875 ) ;
 assign n_n3033 = ( n_n3398 ) | ( n_n3050 ) | ( wire18180 ) ;
 assign wire711 = ( (~ i_7_)  &  i_6_  &  n_n219  &  n_n218 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n219  &  n_n218 ) ;
 assign wire87 = ( wire730  &  n_n191 ) | ( wire717  &  n_n191 ) ;
 assign wire877 = ( n_n159  &  n_n124  &  n_n48 ) | ( n_n159  &  n_n48  &  n_n161 ) ;
 assign n_n2948 = ( i_7_  &  i_6_  &  n_n219  &  n_n48 ) | ( (~ i_7_)  &  i_6_  &  n_n219  &  n_n48 ) | ( i_7_  &  (~ i_6_)  &  n_n219  &  n_n48 ) ;
 assign wire16880 = ( (~ i_7_)  &  i_6_  &  n_n19  &  n_n111 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n19  &  n_n111 ) ;
 assign n_n231 = ( wire431 ) | ( wire389 ) | ( n_n7242 ) | ( wire16880 ) ;
 assign wire308 = ( i_15_  &  n_n156  &  n_n211 ) | ( (~ i_15_)  &  n_n156  &  n_n211 ) | ( i_15_  &  n_n156  &  n_n204 ) ;
 assign wire887 = ( i_9_  &  i_10_  &  i_11_  &  wire725 ) | ( i_9_  &  (~ i_10_)  &  i_11_  &  wire725 ) | ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire725 ) | ( (~ i_9_)  &  (~ i_10_)  &  (~ i_11_)  &  wire725 ) ;
 assign wire189 = ( i_8_  &  n_n48  &  n_n220  &  n_n18 ) | ( (~ i_8_)  &  n_n48  &  n_n220  &  n_n18 ) ;
 assign wire299 = ( i_15_  &  n_n211  &  n_n149 ) | ( (~ i_15_)  &  n_n211  &  n_n149 ) | ( i_15_  &  n_n149  &  n_n204 ) ;
 assign wire896 = ( i_8_  &  n_n162  &  n_n220  &  n_n18 ) | ( (~ i_8_)  &  n_n162  &  n_n220  &  n_n18 ) ;
 assign wire894 = ( (~ i_9_)  &  (~ i_10_)  &  i_11_  &  wire725 ) | ( (~ i_9_)  &  i_10_  &  (~ i_11_)  &  wire725 ) ;
 assign wire561 = ( n_n48  &  n_n220  &  wire131  &  n_n161 ) ;
 assign wire4658 = ( wire168  &  wire968 ) | ( wire968  &  wire193 ) | ( wire968  &  wire196 ) ;
 assign wire4659 = ( n_n33  &  n_n55 ) | ( n_n33  &  wire51 ) | ( n_n33  &  wire17215 ) ;
 assign wire17217 = ( n_n31  &  wire181 ) | ( n_n135  &  n_n32 ) ;
 assign wire899 = ( wire129 ) | ( wire130 ) | ( wire304 ) | ( wire306 ) ;
 assign wire200 = ( i_15_  &  n_n211  &  n_n177 ) | ( (~ i_15_)  &  n_n211  &  n_n177 ) | ( i_15_  &  n_n177  &  n_n204 ) ;
 assign wire201 = ( i_15_  &  n_n211  &  n_n170 ) | ( (~ i_15_)  &  n_n211  &  n_n170 ) | ( i_15_  &  n_n170  &  n_n204 ) ;
 assign wire902 = ( wire131 ) | ( wire308 ) | ( wire200 ) | ( wire201 ) ;
 assign wire376 = ( i_15_  &  n_n149  &  n_n213 ) | ( (~ i_15_)  &  n_n149  &  n_n213 ) ;
 assign n_n201 = ( (~ i_14_)  &  i_13_  &  (~ i_12_) ) ;
 assign wire904 = ( i_15_  &  n_n149  &  n_n213 ) | ( (~ i_15_)  &  n_n149  &  n_n213 ) | ( (~ i_15_)  &  n_n149  &  n_n201 ) ;
 assign wire2861 = ( n_n34  &  wire376 ) | ( wire729  &  n_n177  &  n_n34 ) ;
 assign wire18892 = ( n_n36  &  wire175 ) | ( wire729  &  n_n156  &  n_n36 ) ;
 assign n_n1862 = ( wire2861 ) | ( wire18892 ) | ( n_n36  &  wire123 ) ;
 assign wire911 = ( i_15_  &  n_n177  &  n_n213 ) | ( (~ i_15_)  &  n_n177  &  n_n213 ) | ( i_15_  &  n_n170  &  n_n213 ) | ( (~ i_15_)  &  n_n170  &  n_n213 ) ;
 assign wire18901 = ( wire18883 ) | ( wire18884 ) | ( wire18890 ) | ( wire18891 ) ;
 assign n_n1799 = ( n_n1862 ) | ( wire18901 ) | ( _31998 ) ;
 assign wire246 = ( i_15_  &  n_n184  &  n_n213 ) | ( (~ i_15_)  &  n_n184  &  n_n213 ) | ( (~ i_15_)  &  n_n184  &  n_n209 ) ;
 assign wire254 = ( n_n184  &  wire729 ) | ( n_n184  &  wire717 ) | ( n_n184  &  wire726 ) ;
 assign wire913 = ( n_n183 ) | ( wire184 ) | ( wire246 ) | ( wire254 ) ;
 assign n_n2881 = ( n_n218  &  n_n220  &  n_n126  &  wire147 ) ;
 assign wire69 = ( wire729  &  n_n170 ) | ( n_n170  &  wire726 ) ;
 assign n_n1708 = ( n_n123  &  n_n176 ) | ( n_n125  &  wire69 ) ;
 assign wire223 = ( i_15_  &  n_n177  &  n_n213 ) | ( (~ i_15_)  &  n_n177  &  n_n213 ) | ( (~ i_15_)  &  n_n177  &  n_n209 ) ;
 assign wire239 = ( wire729  &  n_n177 ) | ( n_n177  &  wire717 ) | ( n_n177  &  wire726 ) ;
 assign wire916 = ( wire118 ) | ( wire179 ) | ( wire223 ) | ( wire239 ) ;
 assign wire51 = ( wire729  &  n_n191 ) | ( n_n191  &  wire726 ) ;
 assign n_n1717 = ( n_n125  &  n_n176 ) | ( n_n123  &  wire51 ) ;
 assign wire564 = ( n_n33  &  wire127 ) | ( n_n33  &  wire133 ) ;
 assign wire924 = ( n_n183 ) | ( wire184 ) | ( wire246 ) | ( wire254 ) ;
 assign wire2610 = ( n_n33  &  wire349 ) | ( n_n33  &  wire210 ) | ( n_n33  &  wire357 ) ;
 assign wire19138 = ( n_n33  &  wire127 ) | ( n_n33  &  wire133 ) | ( n_n33  &  wire60 ) ;
 assign n_n1170 = ( wire2610 ) | ( wire19138 ) | ( n_n32  &  wire924 ) ;
 assign wire70 = ( wire729  &  n_n199 ) | ( n_n199  &  wire726 ) ;
 assign wire233 = ( wire720  &  n_n216 ) | ( wire715  &  n_n216 ) | ( wire727  &  n_n216 ) ;
 assign wire251 = ( i_15_  &  n_n205  &  n_n216 ) | ( (~ i_15_)  &  n_n205  &  n_n216 ) | ( i_15_  &  n_n216  &  n_n204 ) ;
 assign wire925 = ( wire142 ) | ( wire70 ) | ( wire233 ) | ( wire251 ) ;
 assign wire928 = ( wire721  &  n_n199 ) | ( wire728  &  n_n199 ) | ( wire721  &  n_n216 ) | ( wire728  &  n_n216 ) ;
 assign n_n4674 = ( n_n125  &  n_n198 ) | ( n_n123  &  wire70 ) ;
 assign n_n78 = ( (~ i_9_)  &  (~ i_10_)  &  i_11_  &  wire724 ) ;
 assign n_n974 = ( n_n39  &  wire53 ) | ( n_n38  &  n_n78 ) ;
 assign n_n215 = ( i_14_  &  (~ i_13_)  &  i_12_ ) ;
 assign wire933 = ( i_15_  &  n_n205  &  n_n170 ) | ( (~ i_15_)  &  n_n205  &  n_n170 ) | ( i_15_  &  n_n170  &  n_n215 ) ;
 assign n_n7260 = ( i_7_  &  i_6_  &  n_n219  &  n_n48 ) ;
 assign n_n7266 = ( (~ i_7_)  &  i_6_  &  n_n219  &  n_n218 ) ;
 assign wire19929 = ( i_7_  &  (~ i_6_)  &  n_n219  &  n_n48 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n219  &  n_n48 ) ;
 assign wire19933 = ( n_n7264 ) | ( n_n7262 ) | ( wire19930 ) ;
 assign wire551 = ( (~ i_7_)  &  i_6_  &  n_n218  &  n_n19 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n218  &  n_n19 ) ;
 assign n_n202 = ( i_9_  &  i_10_  &  i_11_  &  wire726 ) ;
 assign n_n72 = ( i_9_  &  i_10_  &  (~ i_11_)  &  wire724 ) ;
 assign n_n131 = ( (~ i_9_)  &  (~ i_10_)  &  i_11_  &  wire721 ) ;
 assign n_n182 = ( (~ i_9_)  &  (~ i_10_)  &  (~ i_11_)  &  wire722 ) ;
 assign n_n143 = ( (~ i_9_)  &  i_10_  &  (~ i_11_)  &  wire726 ) ;
 assign n_n137 = ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire721 ) ;
 assign n_n128 = ( (~ i_9_)  &  i_10_  &  (~ i_11_)  &  wire719 ) ;
 assign n_n190 = ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire720 ) ;
 assign n_n196 = ( (~ i_9_)  &  i_10_  &  i_11_  &  wire722 ) ;
 assign n_n64 = ( i_9_  &  i_10_  &  i_11_  &  wire728 ) ;
 assign n_n175 = ( i_9_  &  (~ i_10_)  &  i_11_  &  wire722 ) ;
 assign n_n171 = ( i_9_  &  (~ i_10_)  &  i_11_  &  wire726 ) ;
 assign n_n7264 = ( i_7_  &  i_6_  &  n_n219  &  n_n218 ) ;
 assign n_n74 = ( i_9_  &  i_10_  &  (~ i_11_)  &  wire730 ) ;
 assign wire566 = ( n_n33  &  wire55 ) | ( n_n33  &  wire149 ) ;
 assign wire670 = ( wire139  &  n_n32 ) | ( n_n32  &  wire128 ) ;
 assign n_n4808 = ( n_n162  &  n_n220  &  n_n161  &  wire128 ) ;
 assign wire683 = ( n_n43  &  wire124 ) | ( n_n43  &  wire128 ) ;
 assign wire524 = ( wire725  &  n_n191  &  n_n43 ) ;
 assign wire672 = ( n_n42  &  wire63 ) | ( n_n42  &  wire48 ) ;
 assign n_n4564 = ( n_n36  &  n_n140 ) | ( n_n34  &  wire153 ) ;
 assign wire709 = ( n_n36  &  n_n63 ) | ( n_n34  &  wire135 ) ;
 assign n_n4169 = ( n_n4564 ) | ( wire709 ) | ( n_n36  &  wire247 ) ;
 assign wire942 = ( wire80 ) | ( wire78 ) | ( n_n55 ) | ( wire252 ) ;
 assign wire359 = ( wire729  &  n_n41  &  n_n216 ) | ( n_n41  &  wire726  &  n_n216 ) ;
 assign n_n1514 = ( n_n38  &  n_n54 ) | ( n_n38  &  n_n52 ) | ( n_n39  &  n_n52 ) ;
 assign wire432 = ( wire154  &  n_n36 ) | ( wire47  &  n_n36 ) ;
 assign wire17034 = ( wire143  &  n_n36 ) | ( n_n34  &  wire68 ) ;
 assign wire17035 = ( n_n36  &  wire181 ) | ( n_n34  &  wire151 ) ;
 assign n_n4996 = ( n_n108  &  n_n148 ) | ( n_n101  &  wire60 ) ;
 assign n_n4994 = ( n_n162  &  n_n220  &  n_n126  &  wire234 ) ;
 assign wire511 = ( n_n108  &  wire60 ) | ( n_n101  &  n_n155 ) ;
 assign wire946 = ( wire155 ) | ( wire215 ) | ( wire234 ) | ( wire220 ) ;
 assign wire449 = ( n_n31  &  wire134 ) | ( n_n31  &  wire156 ) ;
 assign wire656 = ( n_n31  &  wire176 ) | ( n_n31  &  wire123 ) ;
 assign wire17410 = ( n_n30  &  wire55 ) | ( n_n30  &  wire181 ) ;
 assign wire443 = ( n_n31  &  wire154 ) | ( n_n31  &  wire47 ) ;
 assign n_n4240 = ( n_n31  &  wire122 ) | ( n_n30  &  n_n128 ) ;
 assign wire4965 = ( n_n30  &  wire153 ) | ( n_n30  &  wire135 ) ;
 assign wire4966 = ( n_n31  &  wire247 ) | ( wire719  &  n_n31  &  n_n199 ) ;
 assign n_n4154 = ( wire4965 ) | ( wire4966 ) | ( n_n31  &  n_n63 ) ;
 assign wire654 = ( n_n30  &  wire176 ) | ( n_n30  &  wire123 ) ;
 assign wire739 = ( n_n220  &  n_n156  &  n_n111 ) ;
 assign wire279 = ( n_n177  &  wire722 ) | ( n_n177  &  wire727 ) | ( n_n177  &  wire716 ) ;
 assign n_n4602 = ( n_n48  &  n_n220  &  n_n126  &  wire279 ) ;
 assign wire605 = ( n_n39  &  wire279 ) | ( n_n39  &  n_n177  &  wire724 ) ;
 assign wire59 = ( n_n156  &  wire720 ) | ( n_n156  &  wire715 ) ;
 assign n_n5075 = ( n_n65  &  n_n41 ) | ( n_n40  &  wire59 ) ;
 assign wire54 = ( n_n184  &  wire720 ) | ( n_n184  &  wire715 ) ;
 assign wire498 = ( n_n47  &  n_n89 ) | ( n_n46  &  wire54 ) ;
 assign wire951 = ( n_n117 ) | ( wire94 ) | ( wire184 ) | ( wire268 ) ;
 assign n_n6492 = ( n_n156  &  n_n41  &  wire726 ) ;
 assign n_n3413 = ( n_n71  &  n_n41 ) | ( n_n40  &  wire118 ) ;
 assign wire546 = ( wire137  &  n_n46 ) | ( wire146  &  n_n46 ) ;
 assign wire674 = ( n_n47  &  wire134 ) | ( n_n47  &  wire156 ) ;
 assign n_n3889 = ( wire137  &  n_n47 ) | ( wire146  &  n_n47 ) | ( wire131  &  n_n47 ) ;
 assign wire671 = ( wire63  &  n_n46 ) | ( wire48  &  n_n46 ) ;
 assign wire463 = ( i_7_  &  i_6_  &  n_n219  &  n_n48 ) | ( i_7_  &  (~ i_6_)  &  n_n219  &  n_n48 ) ;
 assign wire960 = ( wire55 ) | ( wire127 ) | ( wire158 ) | ( wire133 ) ;
 assign wire959 = ( wire158 ) | ( wire134 ) | ( wire156 ) | ( wire123 ) ;
 assign wire1730 = ( wire129 ) | ( wire139 ) | ( wire124 ) | ( wire128 ) ;
 assign wire18555 = ( n_n125  &  wire52 ) | ( n_n123  &  wire1729 ) ;
 assign wire4485 = ( n_n212  &  wire308 ) | ( n_n212  &  wire201 ) ;
 assign wire4486 = ( n_n197  &  wire299 ) | ( n_n197  &  wire200 ) | ( n_n197  &  wire201 ) ;
 assign wire17367 = ( wire149  &  n_n197 ) | ( n_n212  &  wire176 ) ;
 assign wire17368 = ( wire131  &  n_n197 ) | ( wire149  &  n_n212 ) ;
 assign wire968 = ( i_8_  &  n_n162  &  n_n220  &  n_n157 ) | ( (~ i_8_)  &  n_n162  &  n_n220  &  n_n157 ) ;
 assign wire115 = ( wire717  &  n_n149 ) | ( n_n149  &  wire726 ) | ( n_n149  &  wire724 ) ;
 assign wire116 = ( n_n156  &  wire717 ) | ( n_n156  &  wire726 ) | ( n_n156  &  wire724 ) ;
 assign wire371 = ( i_15_  &  n_n156  &  n_n211 ) | ( (~ i_15_)  &  n_n156  &  n_n211 ) ;
 assign wire17253 = ( i_15_  &  n_n211  &  n_n149 ) | ( (~ i_15_)  &  n_n211  &  n_n149 ) | ( (~ i_15_)  &  n_n149  &  n_n201 ) ;
 assign wire971 = ( wire115 ) | ( wire116 ) | ( wire371 ) | ( wire17253 ) ;
 assign n_n5739 = ( n_n220  &  n_n111  &  n_n161  &  n_n216 ) ;
 assign wire17258 = ( n_n57  &  n_n125 ) | ( n_n53  &  n_n123 ) ;
 assign wire17259 = ( n_n125  &  wire1115 ) | ( n_n123  &  wire1114 ) ;
 assign wire17260 = ( n_n55  &  wire255 ) | ( n_n113  &  n_n182 ) ;
 assign n_n2340 = ( wire17258 ) | ( wire17259 ) | ( wire17260 ) ;
 assign n_n5743 = ( n_n220  &  n_n177  &  n_n111  &  n_n161 ) ;
 assign wire440 = ( n_n220  &  n_n111  &  n_n161  &  n_n191 ) ;
 assign wire973 = ( wire725  &  n_n191 ) | ( wire729  &  n_n191 ) | ( n_n191  &  wire726 ) ;
 assign wire4619 = ( n_n113  &  wire62 ) | ( n_n113  &  wire202 ) ;
 assign wire17268 = ( wire17265 ) | ( wire17266 ) | ( n_n112  &  wire973 ) ;
 assign wire366 = ( i_15_  &  n_n211  &  n_n170 ) | ( (~ i_15_)  &  n_n211  &  n_n170 ) ;
 assign wire17272 = ( i_9_  &  (~ i_10_)  &  i_11_  &  wire729 ) | ( (~ i_9_)  &  (~ i_10_)  &  i_11_  &  wire729 ) ;
 assign wire975 = ( wire120 ) | ( wire117 ) | ( wire366 ) | ( wire17272 ) ;
 assign wire979 = ( i_8_  &  n_n218  &  n_n220  &  n_n157 ) | ( (~ i_8_)  &  n_n218  &  n_n220  &  n_n157 ) ;
 assign wire978 = ( i_15_  &  n_n211  &  n_n191 ) | ( (~ i_15_)  &  n_n211  &  n_n191 ) | ( i_15_  &  n_n211  &  n_n199 ) | ( (~ i_15_)  &  n_n211  &  n_n199 ) ;
 assign wire362 = ( i_15_  &  n_n211  &  n_n177 ) | ( (~ i_15_)  &  n_n211  &  n_n177 ) ;
 assign n_n2310 = ( wire524 ) | ( wire526 ) | ( wire4531 ) | ( wire17329 ) ;
 assign wire17333 = ( n_n41  &  n_n102 ) | ( n_n41  &  wire70 ) | ( n_n41  &  n_n202 ) ;
 assign wire397 = ( wire729  &  n_n177  &  n_n41 ) | ( n_n177  &  n_n41  &  wire726 ) ;
 assign wire229 = ( n_n170  &  wire730 ) | ( n_n170  &  wire717 ) | ( n_n170  &  wire724 ) ;
 assign wire265 = ( n_n177  &  wire730 ) | ( n_n177  &  wire717 ) | ( n_n177  &  wire724 ) ;
 assign wire989 = ( i_9_  &  (~ i_10_)  &  i_11_  &  wire721 ) | ( (~ i_9_)  &  (~ i_10_)  &  i_11_  &  wire721 ) | ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire721 ) ;
 assign wire988 = ( i_9_  &  (~ i_10_)  &  i_11_  &  wire721 ) | ( (~ i_9_)  &  (~ i_10_)  &  i_11_  &  wire721 ) | ( i_9_  &  i_10_  &  (~ i_11_)  &  wire721 ) | ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire721 ) ;
 assign wire302 = ( wire729  &  n_n149 ) | ( wire717  &  n_n149 ) | ( n_n149  &  wire718 ) ;
 assign wire303 = ( wire729  &  n_n156 ) | ( n_n156  &  wire717 ) | ( n_n156  &  wire718 ) ;
 assign wire316 = ( i_15_  &  n_n149  &  n_n213 ) | ( (~ i_15_)  &  n_n149  &  n_n213 ) | ( i_15_  &  n_n149  &  n_n207 ) ;
 assign wire18831 = ( i_9_  &  i_10_  &  i_11_  &  wire721 ) | ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire721 ) ;
 assign wire993 = ( wire302 ) | ( wire303 ) | ( wire316 ) | ( wire18831 ) ;
 assign wire18832 = ( _1992 ) | ( _1993 ) | ( wire213  &  _32114 ) ;
 assign wire685 = ( n_n108  &  wire156 ) | ( n_n108  &  wire123 ) ;
 assign n_n5011 = ( n_n108  &  n_n169 ) | ( n_n101  &  wire69 ) ;
 assign wire110 = ( n_n156  &  wire720 ) | ( n_n156  &  wire727 ) ;
 assign n_n1517 = ( n_n39  &  n_n143 ) | ( n_n38  &  wire110 ) ;
 assign wire457 = ( n_n39  &  wire207 ) | ( n_n38  &  n_n143 ) ;
 assign wire572 = ( n_n156  &  wire720  &  _32682 ) | ( n_n156  &  wire727  &  _32682 ) ;
 assign wire1003 = ( n_n170  &  wire715 ) | ( n_n170  &  wire727 ) | ( n_n170  &  wire716 ) ;
 assign wire1006 = ( wire179 ) | ( n_n176 ) | ( wire223 ) | ( wire239 ) ;
 assign n_n832 = ( _32818 ) | ( n_n43  &  wire340 ) | ( n_n43  &  _32815 ) ;
 assign wire1012 = ( i_9_  &  i_10_  &  i_11_  &  wire719 ) | ( (~ i_9_)  &  i_10_  &  i_11_  &  wire719 ) | ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire719 ) ;
 assign wire291 = ( wire722  &  n_n216 ) | ( wire727  &  n_n216 ) | ( n_n216  &  wire716 ) ;
 assign wire297 = ( wire722  &  n_n199 ) | ( wire727  &  n_n199 ) | ( n_n199  &  wire716 ) ;
 assign wire19621 = ( wire720  &  n_n199 ) | ( wire715  &  n_n199 ) | ( n_n199  &  wire724 ) ;
 assign wire1017 = ( wire111 ) | ( wire291 ) | ( wire297 ) | ( wire19621 ) ;
 assign n_n56 = ( (~ i_9_)  &  (~ i_10_)  &  i_11_  &  wire728 ) ;
 assign n_n133 = ( i_9_  &  (~ i_10_)  &  i_11_  &  wire721 ) ;
 assign wire198 = ( n_n156  &  wire730 ) | ( n_n156  &  wire716 ) | ( n_n156  &  wire718 ) ;
 assign wire18773 = ( wire729  &  n_n156 ) | ( wire719  &  n_n199 ) ;
 assign wire1021 = ( wire247 ) | ( wire116 ) | ( wire198 ) | ( wire18773 ) ;
 assign wire186 = ( wire725  &  n_n170 ) | ( n_n170  &  wire721 ) ;
 assign wire217 = ( n_n184  &  wire719 ) | ( n_n184  &  wire721 ) | ( n_n184  &  wire728 ) ;
 assign wire18780 = ( n_n184  &  wire725 ) | ( wire719  &  n_n191 ) ;
 assign wire1023 = ( wire182 ) | ( wire186 ) | ( wire217 ) | ( wire18780 ) ;
 assign wire256 = ( n_n184  &  wire725 ) | ( n_n184  &  wire721 ) ;
 assign wire216 = ( n_n184  &  wire719 ) | ( n_n184  &  wire728 ) ;
 assign wire1022 = ( n_n132 ) | ( wire150 ) | ( wire256 ) | ( wire216 ) ;
 assign wire224 = ( n_n177  &  wire717 ) | ( n_n177  &  wire724 ) | ( n_n177  &  wire718 ) ;
 assign n_n4981 = ( n_n108  &  wire80 ) | ( n_n101  &  n_n59 ) ;
 assign wire208 = ( n_n170  &  wire722 ) | ( n_n170  &  wire715 ) | ( n_n170  &  wire727 ) ;
 assign wire225 = ( n_n170  &  wire717 ) | ( n_n170  &  wire724 ) | ( n_n170  &  wire718 ) ;
 assign wire148 = ( n_n170  &  wire723 ) | ( n_n170  &  wire730 ) | ( n_n170  &  wire716 ) ;
 assign wire17083 = ( wire729  &  n_n170 ) | ( n_n170  &  wire720 ) | ( n_n170  &  wire726 ) ;
 assign wire1030 = ( wire208 ) | ( wire225 ) | ( wire148 ) | ( wire17083 ) ;
 assign n_n4620 = ( n_n41  &  n_n198 ) | ( n_n40  &  wire70 ) ;
 assign wire1173 = ( n_n148 ) | ( wire234 ) | ( wire84 ) | ( wire220 ) ;
 assign wire17528 = ( wire361 ) | ( wire363 ) | ( n_n40  &  wire180 ) ;
 assign n_n4131 = ( wire17528 ) | ( wire426 ) | ( _4657 ) | ( _30108 ) ;
 assign wire17534 = ( n_n3979 ) | ( n_n1542 ) | ( wire645 ) | ( wire664 ) ;
 assign n_n4109 = ( n_n4131 ) | ( wire17537 ) | ( _30119 ) | ( _30120 ) ;
 assign wire249 = ( wire723  &  n_n149 ) | ( wire730  &  n_n149 ) | ( n_n149  &  wire718 ) ;
 assign wire571 = ( wire157  &  n_n40 ) | ( wire725  &  n_n156  &  n_n40 ) ;
 assign wire17033 = ( wire143  &  n_n34 ) | ( wire154  &  n_n34 ) | ( wire47  &  n_n34 ) ;
 assign wire549 = ( n_n41  &  wire85 ) | ( n_n41  &  wire142 ) | ( n_n41  &  n_n214 ) ;
 assign n_n4476 = ( n_n41  &  wire219 ) | ( n_n41  &  wire108 ) | ( n_n41  &  wire258 ) ;
 assign wire537 = ( n_n40  &  wire85 ) | ( n_n40  &  wire142 ) ;
 assign wire4842 = ( n_n40  &  n_n214 ) | ( n_n40  &  wire108 ) | ( n_n40  &  wire258 ) ;
 assign wire17007 = ( n_n41  &  n_n198 ) | ( n_n41  &  wire70 ) | ( n_n40  &  wire70 ) ;
 assign wire621 = ( n_n4476 ) | ( wire537 ) | ( wire4842 ) | ( wire17007 ) ;
 assign wire17553 = ( wire597 ) | ( wire17543 ) | ( wire17548 ) | ( wire17549 ) ;
 assign n_n3417 = ( n_n40  &  wire98 ) | ( n_n41  &  n_n117 ) ;
 assign n_n6384 = ( n_n40  &  wire726  &  n_n216 ) ;
 assign n_n3419 = ( n_n41  &  wire98 ) | ( n_n40  &  n_n102 ) ;
 assign wire1036 = ( n_n89 ) | ( wire93 ) | ( wire241 ) | ( wire273 ) ;
 assign n_n3421 = ( n_n41  &  n_n102 ) | ( n_n40  &  wire81 ) ;
 assign wire391 = ( wire720  &  n_n41  &  n_n216 ) | ( wire715  &  n_n41  &  n_n216 ) ;
 assign wire1041 = ( (~ i_9_)  &  i_10_  &  (~ i_11_)  &  wire729 ) | ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire729 ) ;
 assign wire1044 = ( n_n159  &  n_n218  &  n_n35 ) | ( n_n159  &  n_n218  &  n_n124 ) ;
 assign wire1049 = ( wire131 ) | ( wire129 ) | ( wire304 ) | ( wire200 ) ;
 assign wire4481 = ( n_n197  &  wire130 ) | ( n_n197  &  wire304 ) | ( n_n197  &  wire306 ) ;
 assign wire17374 = ( n_n197  &  wire129 ) | ( n_n212  &  wire130 ) ;
 assign wire526 = ( n_n135  &  n_n43 ) | ( n_n42  &  n_n59 ) ;
 assign wire4531 = ( n_n42  &  wire93 ) | ( n_n184  &  wire725  &  n_n42 ) ;
 assign wire17329 = ( n_n42  &  n_n89 ) | ( n_n41  &  n_n210 ) ;
 assign wire374 = ( wire730  &  n_n199 ) | ( wire717  &  n_n199 ) | ( n_n199  &  wire724 ) ;
 assign wire1056 = ( i_9_  &  (~ i_10_)  &  i_11_  &  wire725 ) | ( i_9_  &  i_10_  &  (~ i_11_)  &  wire725 ) | ( (~ i_9_)  &  i_10_  &  (~ i_11_)  &  wire725 ) ;
 assign wire4505 = ( n_n101  &  wire202 ) | ( n_n101  &  wire17349 ) | ( n_n101  &  wire17350 ) ;
 assign wire4506 = ( n_n108  &  wire265 ) | ( n_n108  &  wire17352 ) | ( n_n108  &  wire17353 ) ;
 assign wire4508 = ( n_n101  &  wire307 ) | ( wire722  &  n_n191  &  n_n101 ) ;
 assign wire4509 = ( n_n108  &  wire62 ) | ( n_n108  &  wire202 ) ;
 assign n_n2257 = ( wire4505 ) | ( wire4506 ) | ( wire4508 ) | ( wire4509 ) ;
 assign wire1060 = ( wire69 ) | ( n_n175 ) | ( wire229 ) | ( wire265 ) ;
 assign wire263 = ( wire730  &  n_n216 ) | ( wire717  &  n_n216 ) | ( wire724  &  n_n216 ) ;
 assign wire17361 = ( wire729  &  n_n199 ) | ( wire722  &  n_n199 ) | ( n_n199  &  wire726 ) ;
 assign wire1064 = ( wire86 ) | ( wire374 ) | ( wire263 ) | ( wire17361 ) ;
 assign wire250 = ( n_n177  &  wire723 ) | ( n_n177  &  wire730 ) | ( n_n177  &  wire716 ) ;
 assign wire1069 = ( wire179 ) | ( n_n176 ) | ( wire223 ) | ( wire239 ) ;
 assign wire62 = ( n_n184  &  wire729 ) | ( n_n184  &  wire726 ) ;
 assign n_n5019 = ( n_n101  &  n_n190 ) | ( n_n108  &  wire62 ) ;
 assign wire19179 = ( wire729  &  n_n191 ) | ( wire717  &  n_n191 ) | ( n_n191  &  wire726 ) ;
 assign wire1070 = ( wire139 ) | ( wire128 ) | ( wire54 ) | ( wire19179 ) ;
 assign wire65 = ( wire721  &  n_n191 ) | ( wire728  &  n_n191 ) ;
 assign wire1902 = ( (~ i_9_)  &  i_10_  &  i_11_ ) | ( (~ i_9_)  &  (~ i_10_)  &  (~ i_11_) ) ;
 assign wire16987 = ( i_7_  &  i_8_  &  i_6_ ) ;
 assign wire760 = ( n_n220  &  n_n111  &  wire1902  &  wire16987 ) ;
 assign wire1072 = ( (~ i_9_)  &  (~ i_10_)  &  i_11_ ) | ( (~ i_9_)  &  i_10_  &  (~ i_11_) ) ;
 assign wire385 = ( i_15_  &  n_n205  &  n_n199 ) | ( (~ i_15_)  &  n_n205  &  n_n199 ) ;
 assign wire19196 = ( wire729  &  n_n199 ) | ( wire727  &  n_n199 ) ;
 assign wire19197 = ( wire720  &  n_n199 ) | ( wire715  &  n_n199 ) | ( wire717  &  n_n199 ) ;
 assign wire1075 = ( wire108 ) | ( wire385 ) | ( wire19196 ) | ( wire19197 ) ;
 assign wire277 = ( n_n170  &  wire720 ) | ( n_n170  &  wire715 ) | ( n_n170  &  wire727 ) ;
 assign wire1077 = ( wire98 ) | ( wire51 ) | ( wire148 ) | ( wire277 ) ;
 assign wire276 = ( n_n184  &  wire720 ) | ( n_n184  &  wire715 ) | ( n_n184  &  wire727 ) ;
 assign wire211 = ( n_n184  &  wire723 ) | ( n_n184  &  wire730 ) | ( n_n184  &  wire716 ) ;
 assign wire271 = ( i_15_  &  n_n184  &  n_n205 ) | ( (~ i_15_)  &  n_n184  &  n_n205 ) | ( i_15_  &  n_n184  &  n_n204 ) ;
 assign wire1079 = ( wire51 ) | ( wire276 ) | ( wire211 ) | ( wire271 ) ;
 assign n_n972 = ( n_n38  &  n_n84 ) | ( n_n39  &  wire110 ) ;
 assign wire1084 = ( i_15_  &  n_n191  &  n_n207 ) | ( (~ i_15_)  &  n_n191  &  n_n207 ) | ( i_15_  &  n_n191  &  n_n209 ) ;
 assign wire1089 = ( i_9_  &  (~ i_10_)  &  i_11_  &  wire719 ) | ( i_9_  &  i_10_  &  (~ i_11_)  &  wire719 ) | ( (~ i_9_)  &  i_10_  &  (~ i_11_)  &  wire719 ) ;
 assign wire1087 = ( i_9_  &  (~ i_10_)  &  i_11_  &  wire719 ) | ( i_9_  &  i_10_  &  (~ i_11_)  &  wire719 ) | ( (~ i_9_)  &  i_10_  &  (~ i_11_)  &  wire719 ) ;
 assign wire1090 = ( i_9_  &  i_10_  &  i_11_  &  wire728 ) | ( (~ i_9_)  &  i_10_  &  i_11_  &  wire728 ) | ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire728 ) ;
 assign wire3433 = ( n_n5  &  n_n144 ) | ( n_n5  &  n_n186 ) | ( n_n5  &  wire170 ) ;
 assign wire3434 = ( n_n4  &  wire95 ) | ( n_n4  &  wire729  &  n_n191 ) ;
 assign wire18316 = ( wire3435 ) | ( n_n4  &  wire729  &  n_n156 ) ;
 assign n_n164 = ( (~ i_9_)  &  (~ i_10_)  &  i_11_  &  wire726 ) ;
 assign n_n5103 = ( n_n132  &  n_n47 ) | ( n_n46  &  wire186 ) ;
 assign wire212 = ( wire719  &  n_n216 ) | ( wire728  &  n_n216 ) ;
 assign n_n5067 = ( n_n41  &  n_n61 ) | ( n_n40  &  wire212 ) ;
 assign wire221 = ( wire730  &  n_n149 ) | ( n_n149  &  wire716 ) | ( n_n149  &  wire718 ) ;
 assign wire298 = ( wire722  &  n_n149 ) | ( wire723  &  n_n149 ) | ( wire727  &  n_n149 ) ;
 assign wire1096 = ( n_n65 ) | ( wire115 ) | ( wire221 ) | ( wire298 ) ;
 assign wire591 = ( n_n108  &  wire208 ) | ( n_n108  &  wire148 ) ;
 assign wire515 = ( wire725  &  n_n177  &  n_n125 ) ;
 assign wire4948 = ( n_n220  &  n_n170  &  n_n111  &  wire16987 ) ;
 assign wire657 = ( n_n5743 ) | ( wire4948 ) ;
 assign wire1789 = ( n_n169 ) | ( wire208 ) | ( wire225 ) | ( wire148 ) ;
 assign wire17013 = ( wire397 ) | ( wire361 ) | ( n_n40  &  wire180 ) ;
 assign n_n4424 = ( wire17013 ) | ( wire696 ) | ( _5873 ) | ( _29156 ) ;
 assign wire518 = ( n_n40  &  n_n176 ) | ( n_n41  &  wire69 ) ;
 assign wire57 = ( wire729  &  n_n177 ) | ( n_n177  &  wire726 ) ;
 assign wire653 = ( n_n40  &  wire224 ) | ( n_n40  &  wire57 ) ;
 assign wire694 = ( n_n41  &  wire208 ) | ( n_n41  &  wire148 ) ;
 assign wire17018 = ( n_n5060 ) | ( n_n5059 ) | ( n_n5058 ) | ( wire4900 ) ;
 assign wire17019 = ( wire4904 ) | ( wire4905 ) | ( wire4908 ) | ( wire17016 ) ;
 assign n_n4404 = ( n_n4424 ) | ( _29191 ) | ( _29192 ) | ( _29193 ) ;
 assign wire666 = ( n_n47  &  wire150 ) | ( n_n46  &  wire182 ) ;
 assign wire17050 = ( wire597 ) | ( wire620 ) | ( wire17041 ) | ( wire17045 ) ;
 assign wire17064 = ( wire17060 ) | ( wire17061 ) | ( wire17063 ) ;
 assign n_n4312 = ( n_n48  &  wire714  &  wire157  &  n_n18 ) ;
 assign wire141 = ( wire725  &  n_n216 ) | ( wire721  &  n_n216 ) | ( wire728  &  n_n216 ) ;
 assign wire258 = ( wire717  &  n_n199 ) | ( n_n199  &  wire724 ) | ( n_n199  &  wire718 ) ;
 assign wire125 = ( wire719  &  n_n216 ) | ( wire721  &  n_n216 ) | ( wire728  &  n_n216 ) ;
 assign n_n4566 = ( n_n218  &  wire714  &  n_n157  &  wire125 ) ;
 assign wire46 = ( n_n177  &  wire720 ) | ( n_n177  &  wire722 ) | ( n_n177  &  wire715 ) ;
 assign n_n1553 = ( n_n41  &  n_n176 ) | ( n_n40  &  wire51 ) ;
 assign wire209 = ( wire719  &  n_n170 ) | ( n_n170  &  wire728 ) ;
 assign n_n5059 = ( n_n41  &  n_n57 ) | ( n_n40  &  wire209 ) ;
 assign n_n5058 = ( n_n132  &  n_n41 ) | ( n_n40  &  wire186 ) ;
 assign wire577 = ( wire143  &  n_n47 ) | ( n_n47  &  wire181 ) ;
 assign wire1115 = ( i_9_  &  i_10_  &  (~ i_11_)  &  wire725 ) | ( (~ i_9_)  &  i_10_  &  (~ i_11_)  &  wire725 ) ;
 assign wire1114 = ( i_9_  &  (~ i_10_)  &  i_11_  &  wire725 ) | ( (~ i_9_)  &  i_10_  &  (~ i_11_)  &  wire725 ) ;
 assign wire1116 = ( n_n177  &  wire722 ) | ( n_n170  &  wire722 ) | ( n_n177  &  wire724 ) ;
 assign wire1117 = ( (~ i_9_)  &  (~ i_10_)  &  i_11_  &  wire725 ) | ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire725 ) ;
 assign wire1120 = ( n_n156  &  wire730 ) | ( wire730  &  n_n149 ) | ( n_n149  &  wire726 ) ;
 assign wire358 = ( i_15_  &  n_n211  &  n_n216 ) | ( (~ i_15_)  &  n_n211  &  n_n216 ) ;
 assign wire17395 = ( i_15_  &  n_n211  &  n_n199 ) | ( (~ i_15_)  &  n_n211  &  n_n199 ) | ( (~ i_15_)  &  n_n199  &  n_n201 ) ;
 assign wire1124 = ( wire164 ) | ( wire243 ) | ( wire358 ) | ( wire17395 ) ;
 assign wire1126 = ( n_n156  &  wire723 ) | ( wire723  &  n_n149 ) | ( n_n156  &  wire718 ) | ( n_n149  &  wire718 ) ;
 assign wire292 = ( wire729  &  n_n191 ) | ( wire717  &  n_n191 ) | ( n_n191  &  wire718 ) ;
 assign wire311 = ( i_15_  &  n_n184  &  n_n213 ) | ( (~ i_15_)  &  n_n184  &  n_n213 ) | ( i_15_  &  n_n184  &  n_n207 ) ;
 assign wire317 = ( n_n184  &  wire729 ) | ( n_n184  &  wire717 ) | ( n_n184  &  wire718 ) ;
 assign wire319 = ( i_15_  &  n_n191  &  n_n213 ) | ( (~ i_15_)  &  n_n191  &  n_n213 ) | ( i_15_  &  n_n191  &  n_n207 ) ;
 assign wire1129 = ( wire292 ) | ( wire311 ) | ( wire317 ) | ( wire319 ) ;
 assign wire321 = ( i_15_  &  n_n156  &  n_n213 ) | ( (~ i_15_)  &  n_n156  &  n_n213 ) | ( i_15_  &  n_n156  &  n_n207 ) ;
 assign wire326 = ( i_15_  &  n_n170  &  n_n213 ) | ( (~ i_15_)  &  n_n170  &  n_n213 ) | ( i_15_  &  n_n170  &  n_n207 ) ;
 assign wire327 = ( wire729  &  n_n170 ) | ( n_n170  &  wire717 ) | ( n_n170  &  wire718 ) ;
 assign wire1132 = ( wire303 ) | ( wire321 ) | ( wire326 ) | ( wire327 ) ;
 assign wire197 = ( i_15_  &  n_n216  &  n_n213 ) | ( (~ i_15_)  &  n_n216  &  n_n213 ) | ( i_15_  &  n_n216  &  n_n207 ) ;
 assign wire203 = ( wire729  &  n_n199 ) | ( wire717  &  n_n199 ) | ( n_n199  &  wire718 ) ;
 assign wire309 = ( wire729  &  n_n216 ) | ( wire717  &  n_n216 ) | ( n_n216  &  wire718 ) ;
 assign wire323 = ( i_15_  &  n_n199  &  n_n213 ) | ( (~ i_15_)  &  n_n199  &  n_n213 ) | ( i_15_  &  n_n199  &  n_n207 ) ;
 assign wire1135 = ( wire197 ) | ( wire203 ) | ( wire309 ) | ( wire323 ) ;
 assign wire1136 = ( i_15_  &  n_n199  &  n_n213 ) | ( (~ i_15_)  &  n_n199  &  n_n213 ) | ( (~ i_15_)  &  n_n199  &  n_n201 ) ;
 assign wire83 = ( n_n156  &  wire721 ) | ( n_n156  &  wire728 ) ;
 assign wire384 = ( n_n177  &  wire720 ) | ( n_n177  &  wire715 ) | ( n_n177  &  wire727 ) ;
 assign wire1143 = ( n_n184  &  wire721 ) | ( n_n184  &  wire728 ) | ( wire721  &  n_n191 ) | ( wire728  &  n_n191 ) ;
 assign wire330 = ( wire729  &  n_n199 ) | ( wire717  &  n_n199 ) | ( n_n199  &  wire726 ) ;
 assign wire1145 = ( wire98 ) | ( wire52 ) | ( wire51 ) | ( wire330 ) ;
 assign wire19221 = ( n_n184  &  wire729 ) | ( n_n177  &  wire720 ) ;
 assign wire1147 = ( wire276 ) | ( wire211 ) | ( wire271 ) | ( wire19221 ) ;
 assign wire1150 = ( n_n102 ) | ( wire142 ) | ( wire233 ) | ( wire251 ) ;
 assign wire1152 = ( wire179 ) | ( n_n172 ) | ( wire223 ) | ( wire271 ) ;
 assign wire500 = ( wire729  &  n_n191  &  _30362 ) | ( n_n191  &  wire726  &  _30362 ) ;
 assign wire1154 = ( wire63 ) | ( wire52 ) | ( wire276 ) | ( wire211 ) ;
 assign wire1153 = ( n_n183 ) | ( wire184 ) | ( wire246 ) | ( wire254 ) ;
 assign n_n3415 = ( n_n41  &  wire53 ) | ( n_n40  &  n_n77 ) ;
 assign wire1160 = ( i_9_  &  (~ i_10_)  &  i_11_  &  wire719 ) | ( i_9_  &  i_10_  &  (~ i_11_)  &  wire719 ) ;
 assign wire1159 = ( (~ i_9_)  &  (~ i_10_)  &  i_11_  &  wire719 ) | ( (~ i_9_)  &  i_10_  &  (~ i_11_)  &  wire719 ) ;
 assign n_n7262 = ( (~ i_7_)  &  i_6_  &  n_n219  &  n_n48 ) ;
 assign n_n73 = ( i_9_  &  i_10_  &  (~ i_11_)  &  wire718 ) ;
 assign n_n1606 = ( n_n46  &  n_n169 ) | ( n_n47  &  wire57 ) ;
 assign wire100 = ( n_n177  &  wire722 ) | ( n_n177  &  wire715 ) | ( n_n177  &  wire727 ) ;
 assign wire1170 = ( n_n176 ) | ( wire224 ) | ( wire250 ) | ( wire100 ) ;
 assign n_n3979 = ( n_n40  &  wire90 ) | ( n_n41  &  n_n142 ) ;
 assign wire361 = ( wire729  &  n_n40  &  n_n216 ) | ( n_n40  &  wire726  &  n_n216 ) ;
 assign wire363 = ( wire729  &  n_n156  &  n_n41 ) | ( n_n156  &  n_n41  &  wire726 ) ;
 assign wire426 = ( n_n41  &  wire215 ) | ( n_n156  &  wire720  &  n_n41 ) ;
 assign wire442 = ( n_n41  &  wire155 ) | ( n_n41  &  wire205 ) ;
 assign wire1174 = ( wire94 ) | ( wire184 ) | ( wire268 ) | ( wire54 ) ;
 assign wire1177 = ( i_9_  &  i_10_  &  i_11_  &  wire725 ) | ( (~ i_9_)  &  i_10_  &  i_11_  &  wire725 ) | ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire725 ) ;
 assign wire1176 = ( wire1177 ) | ( wire729  &  n_n156 ) ;
 assign wire1179 = ( i_9_  &  (~ i_10_)  &  i_11_  &  wire725 ) | ( (~ i_9_)  &  (~ i_10_)  &  i_11_  &  wire725 ) | ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire725 ) ;
 assign wire1178 = ( i_9_  &  (~ i_10_)  &  i_11_  &  wire725 ) | ( (~ i_9_)  &  (~ i_10_)  &  i_11_  &  wire725 ) | ( i_9_  &  i_10_  &  (~ i_11_)  &  wire725 ) | ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire725 ) ;
 assign wire655 = ( wire725  &  n_n31  &  n_n216 ) ;
 assign wire1190 = ( i_9_  &  (~ i_10_)  &  i_11_  &  wire725 ) | ( i_9_  &  i_10_  &  (~ i_11_)  &  wire725 ) | ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire725 ) ;
 assign wire1189 = ( i_9_  &  (~ i_10_)  &  i_11_  &  wire725 ) | ( i_9_  &  i_10_  &  (~ i_11_)  &  wire725 ) | ( (~ i_9_)  &  (~ i_10_)  &  (~ i_11_)  &  wire725 ) ;
 assign wire1188 = ( (~ i_9_)  &  (~ i_10_)  &  i_11_  &  wire725 ) | ( (~ i_9_)  &  i_10_  &  (~ i_11_)  &  wire725 ) ;
 assign wire380 = ( n_n177  &  wire723 ) | ( n_n177  &  wire716 ) | ( n_n177  &  wire718 ) ;
 assign wire18986 = ( wire729  &  n_n177 ) | ( n_n177  &  wire715 ) | ( n_n177  &  wire717 ) ;
 assign wire1194 = ( wire380 ) | ( wire18986 ) ;
 assign wire364 = ( i_15_  &  n_n216  &  n_n213 ) | ( (~ i_15_)  &  n_n216  &  n_n213 ) ;
 assign wire1197 = ( i_9_  &  (~ i_10_)  &  i_11_  &  wire721 ) | ( i_9_  &  i_10_  &  (~ i_11_)  &  wire721 ) | ( (~ i_9_)  &  (~ i_10_)  &  (~ i_11_)  &  wire721 ) ;
 assign wire1196 = ( i_9_  &  (~ i_10_)  &  i_11_  &  wire721 ) | ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire721 ) ;
 assign wire1195 = ( (~ i_9_)  &  (~ i_10_)  &  i_11_  &  wire721 ) | ( (~ i_9_)  &  i_10_  &  (~ i_11_)  &  wire721 ) ;
 assign wire18834 = ( n_n30  &  wire1196 ) | ( n_n31  &  wire1195 ) | ( n_n30  &  wire1195 ) ;
 assign wire1401 = ( wire292 ) | ( wire311 ) | ( wire317 ) | ( wire319 ) ;
 assign wire331 = ( i_15_  &  n_n177  &  n_n213 ) | ( (~ i_15_)  &  n_n177  &  n_n213 ) | ( i_15_  &  n_n177  &  n_n207 ) ;
 assign n_n1826 = ( n_n47  &  wire1401 ) | ( n_n46  &  wire1401 ) | ( n_n47  &  wire331 ) ;
 assign wire1200 = ( wire197 ) | ( wire203 ) | ( wire309 ) | ( wire323 ) ;
 assign wire1199 = ( i_8_  &  n_n48  &  n_n220  &  n_n18 ) | ( (~ i_8_)  &  n_n48  &  n_n220  &  n_n18 ) ;
 assign wire18961 = ( wire2775 ) | ( wire721  &  n_n199  &  wire228 ) ;
 assign wire18962 = ( wire2776 ) | ( wire18955 ) | ( n_n108  &  wire1469 ) ;
 assign wire18966 = ( wire18965 ) | ( wire1200  &  wire1199 ) ;
 assign n_n1803 = ( n_n1826 ) | ( wire18961 ) | ( wire18962 ) | ( wire18966 ) ;
 assign wire18981 = ( n_n139  &  wire189 ) | ( n_n47  &  wire1766 ) ;
 assign wire312 = ( wire729  &  n_n177 ) | ( n_n177  &  wire717 ) | ( n_n177  &  wire718 ) ;
 assign wire1201 = ( wire326 ) | ( wire327 ) | ( wire331 ) | ( wire312 ) ;
 assign wire261 = ( wire723  &  n_n216 ) | ( n_n216  &  wire716 ) | ( n_n216  &  wire718 ) ;
 assign wire264 = ( wire723  &  n_n199 ) | ( n_n199  &  wire716 ) | ( n_n199  &  wire718 ) ;
 assign wire375 = ( wire729  &  n_n216 ) | ( wire717  &  n_n216 ) ;
 assign wire19001 = ( wire729  &  n_n199 ) | ( wire715  &  n_n199 ) | ( wire717  &  n_n199 ) ;
 assign wire1205 = ( wire261 ) | ( wire264 ) | ( wire375 ) | ( wire19001 ) ;
 assign wire1207 = ( n_n177  &  wire721 ) | ( n_n170  &  wire721 ) | ( n_n177  &  wire728 ) | ( n_n170  &  wire728 ) ;
 assign wire92 = ( wire721  &  n_n199 ) | ( wire728  &  n_n199 ) ;
 assign wire19413 = ( n_n201  &  _32515 ) | ( n_n201  &  _32516 ) ;
 assign wire19414 = ( n_n184  &  wire728 ) | ( wire721  &  n_n216 ) | ( wire728  &  n_n216 ) ;
 assign wire1211 = ( wire232 ) | ( wire92 ) | ( wire19413 ) | ( wire19414 ) ;
 assign n_n1542 = ( n_n41  &  n_n148 ) | ( n_n40  &  wire60 ) ;
 assign n_n4641 = ( n_n46  &  n_n214 ) | ( n_n47  &  wire70 ) ;
 assign wire693 = ( n_n47  &  wire74 ) | ( n_n47  &  wire68 ) ;
 assign wire169 = ( wire723  &  n_n216 ) | ( wire727  &  n_n216 ) ;
 assign wire19320 = ( wire715  &  n_n216 ) | ( wire717  &  n_n216 ) ;
 assign wire1214 = ( wire86 ) | ( wire162 ) | ( wire169 ) | ( wire19320 ) ;
 assign wire274 = ( i_15_  &  n_n205  &  n_n170 ) | ( (~ i_15_)  &  n_n205  &  n_n170 ) | ( i_15_  &  n_n170  &  n_n204 ) ;
 assign wire1216 = ( n_n155 ) | ( wire148 ) | ( wire277 ) | ( wire274 ) ;
 assign wire1218 = ( i_15_  &  n_n205  &  n_n216 ) | ( (~ i_15_)  &  n_n205  &  n_n216 ) | ( i_15_  &  n_n216  &  n_n215 ) ;
 assign wire2083 = ( n_n36  &  wire385 ) | ( wire720  &  n_n36  &  n_n191 ) ;
 assign n_n369 = ( wire2083 ) | ( wire154  &  n_n34 ) | ( n_n34  &  wire1218 ) ;
 assign wire335 = ( wire720  &  n_n216 ) | ( wire727  &  n_n216 ) ;
 assign wire652 = ( n_n46  &  wire218 ) | ( n_n47  &  wire141 ) ;
 assign wire1229 = ( n_n159  &  n_n124  &  n_n48 ) | ( n_n159  &  n_n48  &  n_n161 ) ;
 assign wire18706 = ( wire18703 ) | ( n_n14  &  wire730  &  n_n149 ) ;
 assign n_n3054 = ( wire18706 ) | ( wire18704 ) | ( wire18705 ) | ( _2661 ) ;
 assign n_n2770 = ( wire137  &  n_n197 ) | ( wire146  &  n_n197 ) | ( wire131  &  n_n197 ) ;
 assign wire1234 = ( wire116 ) | ( i_15_  &  n_n156  &  n_n211 ) | ( (~ i_15_)  &  n_n156  &  n_n211 ) ;
 assign wire412 = ( (~ i_9_)  &  (~ i_10_)  &  i_11_ ) | ( (~ i_9_)  &  i_10_  &  (~ i_11_) ) ;
 assign wire1239 = ( i_15_  &  n_n191  &  n_n204 ) | ( i_15_  &  n_n191  &  n_n201 ) | ( (~ i_15_)  &  n_n191  &  n_n201 ) ;
 assign wire18938 = ( n_n113  &  n_n115 ) | ( n_n108  &  n_n107 ) ;
 assign wire18939 = ( wire760 ) | ( wire2797 ) | ( n_n112  &  wire1239 ) ;
 assign n_n3638 = ( n_n218  &  wire714  &  n_n157  &  wire139 ) ;
 assign wire1242 = ( i_9_  &  i_10_  &  i_11_  &  wire721 ) | ( (~ i_9_)  &  i_10_  &  i_11_  &  wire721 ) | ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire721 ) ;
 assign wire1244 = ( i_9_  &  (~ i_10_)  &  i_11_  &  wire721 ) | ( i_9_  &  i_10_  &  (~ i_11_)  &  wire721 ) | ( (~ i_9_)  &  i_10_  &  (~ i_11_)  &  wire721 ) ;
 assign wire1243 = ( i_8_  &  n_n16  &  n_n218  &  n_n220 ) | ( (~ i_8_)  &  n_n16  &  n_n218  &  n_n220 ) ;
 assign wire1246 = ( wire292 ) | ( wire311 ) | ( wire317 ) | ( wire319 ) ;
 assign n_n1811 = ( n_n30  &  wire309 ) | ( n_n31  &  wire1246 ) | ( n_n30  &  wire1246 ) ;
 assign wire1247 = ( i_9_  &  i_10_  &  (~ i_11_)  &  wire721 ) | ( (~ i_9_)  &  i_10_  &  (~ i_11_)  &  wire721 ) ;
 assign wire1251 = ( n_n177  &  wire721 ) | ( n_n170  &  wire721 ) | ( n_n177  &  wire728 ) | ( n_n170  &  wire728 ) ;
 assign wire1255 = ( wire63 ) | ( wire98 ) | ( wire206 ) | ( wire330 ) ;
 assign wire1257 = ( n_n177  &  wire721 ) | ( n_n149  &  wire721 ) | ( n_n177  &  wire728 ) | ( n_n149  &  wire728 ) ;
 assign wire4869 = ( n_n39  &  wire237 ) | ( n_n39  &  n_n170  &  wire724 ) ;
 assign n_n817 = ( n_n974 ) | ( wire4869 ) | ( n_n38  &  wire104 ) ;
 assign wire167 = ( i_15_  &  n_n191  &  n_n207 ) | ( (~ i_15_)  &  n_n191  &  n_n207 ) | ( (~ i_15_)  &  n_n191  &  n_n209 ) ;
 assign wire2329 = ( n_n162  &  n_n220  &  n_n200  &  wire167 ) ;
 assign wire2331 = ( n_n184  &  wire719  &  n_n32 ) ;
 assign wire19480 = ( wire719  &  n_n149  &  n_n33 ) | ( wire719  &  n_n33  &  n_n191 ) ;
 assign wire19481 = ( n_n132  &  n_n33 ) | ( n_n31  &  wire111 ) ;
 assign wire320 = ( wire722  &  n_n191 ) | ( wire727  &  n_n191 ) | ( n_n191  &  wire716 ) ;
 assign wire19660 = ( wire720  &  n_n191 ) | ( wire715  &  n_n191 ) | ( n_n191  &  wire724 ) ;
 assign wire1259 = ( wire320 ) | ( wire19660 ) ;
 assign wire195 = ( n_n184  &  wire722 ) | ( n_n184  &  wire727 ) | ( n_n184  &  wire716 ) ;
 assign wire19663 = ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire724 ) | ( (~ i_9_)  &  (~ i_10_)  &  (~ i_11_)  &  wire724 ) ;
 assign wire1261 = ( wire98 ) | ( wire320 ) | ( wire195 ) | ( wire19663 ) ;
 assign wire1260 = ( n_n118 ) | ( wire104 ) | ( wire54 ) | ( wire195 ) ;
 assign wire1263 = ( wire182 ) | ( wire725  &  n_n177 ) ;
 assign wire686 = ( wire132  &  n_n47 ) | ( n_n47  &  wire126 ) ;
 assign wire1271 = ( wire132 ) | ( wire149 ) | ( wire126 ) | ( wire147 ) ;
 assign n_n4692 = ( n_n218  &  n_n220  &  n_n200  &  wire46 ) ;
 assign wire1277 = ( i_8_  &  n_n162  &  n_n220  &  n_n18 ) | ( (~ i_8_)  &  n_n162  &  n_n220  &  n_n18 ) ;
 assign wire175 = ( i_15_  &  n_n156  &  n_n213 ) | ( (~ i_15_)  &  n_n156  &  n_n213 ) ;
 assign wire383 = ( i_15_  &  n_n177  &  n_n213 ) | ( (~ i_15_)  &  n_n177  &  n_n213 ) ;
 assign wire1279 = ( i_15_  &  n_n191  &  n_n213 ) | ( (~ i_15_)  &  n_n191  &  n_n213 ) | ( (~ i_15_)  &  n_n191  &  n_n201 ) ;
 assign wire1285 = ( wire326 ) | ( wire327 ) | ( wire331 ) | ( wire312 ) ;
 assign wire1287 = ( n_n149  &  wire721 ) | ( n_n149  &  wire728 ) ;
 assign wire1286 = ( n_n156  &  wire721 ) | ( n_n149  &  wire721 ) | ( n_n156  &  wire728 ) | ( n_n149  &  wire728 ) ;
 assign wire473 = ( n_n115  &  n_n32 ) | ( n_n33  &  n_n137 ) ;
 assign wire19253 = ( n_n177  &  wire720 ) | ( wire720  &  n_n149 ) | ( wire715  &  n_n149 ) ;
 assign wire1290 = ( wire179 ) | ( wire223 ) | ( wire239 ) | ( wire19253 ) ;
 assign wire19250 = ( wire729  &  n_n156 ) | ( wire729  &  n_n170 ) | ( n_n170  &  wire726 ) ;
 assign wire1289 = ( wire155 ) | ( wire227 ) | ( wire232 ) | ( wire19250 ) ;
 assign wire19260 = ( wire729  &  n_n156 ) | ( wire729  &  n_n149 ) | ( n_n149  &  wire726 ) ;
 assign wire1292 = ( wire155 ) | ( wire227 ) | ( wire232 ) | ( wire19260 ) ;
 assign wire557 = ( wire126  &  n_n212 ) | ( wire147  &  n_n212 ) ;
 assign wire1294 = ( n_n77 ) | ( wire148 ) | ( wire277 ) | ( wire274 ) ;
 assign wire1293 = ( wire179 ) | ( wire53 ) | ( wire223 ) | ( wire239 ) ;
 assign n_n1566 = ( n_n43  &  n_n115 ) | ( n_n42  &  wire65 ) ;
 assign wire88 = ( n_n184  &  wire721 ) | ( n_n184  &  wire728 ) ;
 assign wire1295 = ( wire727  &  n_n216 ) | ( wire717  &  n_n216 ) | ( n_n216  &  wire718 ) ;
 assign n_n1575 = ( n_n43  &  n_n183 ) | ( n_n42  &  wire62 ) ;
 assign wire349 = ( i_15_  &  n_n205  &  n_n191 ) | ( (~ i_15_)  &  n_n205  &  n_n191 ) | ( i_15_  &  n_n191  &  n_n204 ) ;
 assign wire1297 = ( wire184 ) | ( wire246 ) | ( wire254 ) | ( wire349 ) ;
 assign wire19464 = ( wire720  &  n_n149 ) | ( wire715  &  n_n149 ) | ( n_n149  &  wire724 ) ;
 assign wire1302 = ( wire290 ) | ( wire199 ) | ( n_n72 ) | ( wire19464 ) ;
 assign wire19469 = ( n_n184  &  wire720 ) | ( n_n184  &  wire715 ) | ( n_n184  &  wire724 ) ;
 assign wire1305 = ( wire98 ) | ( wire320 ) | ( wire195 ) | ( wire19469 ) ;
 assign wire329 = ( n_n170  &  wire723 ) | ( n_n170  &  wire730 ) | ( n_n170  &  wire718 ) ;
 assign wire1311 = ( wire329 ) | ( n_n170  &  wire726 ) ;
 assign wire171 = ( wire719  &  n_n191 ) | ( wire728  &  n_n191 ) ;
 assign n_n2859 = ( n_n123  &  n_n63 ) | ( n_n125  &  wire171 ) ;
 assign n_n4657 = ( n_n218  &  n_n220  &  n_n126  &  wire182 ) ;
 assign wire160 = ( wire725  &  n_n191 ) | ( wire721  &  n_n191 ) ;
 assign wire174 = ( wire725  &  n_n177 ) | ( n_n177  &  wire721 ) | ( n_n177  &  wire728 ) ;
 assign wire651 = ( wire157  &  n_n47 ) | ( n_n46  &  wire174 ) ;
 assign n_n3570 = ( n_n108  &  wire156 ) | ( n_n108  &  wire176 ) | ( n_n108  &  wire123 ) ;
 assign n_n3573 = ( wire137  &  n_n108 ) | ( wire146  &  n_n108 ) | ( n_n108  &  wire46 ) ;
 assign wire1319 = ( wire137 ) | ( wire146 ) | ( wire131 ) | ( wire46 ) ;
 assign wire4182 = ( wire131  &  n_n108 ) | ( n_n108  &  wire134 ) ;
 assign n_n3823 = ( n_n3573 ) | ( wire4182 ) | ( n_n101  &  wire1319 ) ;
 assign wire222 = ( wire719  &  n_n191 ) | ( wire721  &  n_n191 ) | ( wire728  &  n_n191 ) ;
 assign wire1321 = ( n_n134 ) | ( wire214 ) | ( wire174 ) | ( wire222 ) ;
 assign wire1326 = ( n_n65 ) | ( wire115 ) | ( wire221 ) | ( wire298 ) ;
 assign n_n5070 = ( n_n41  &  wire214 ) | ( n_n40  &  n_n140 ) ;
 assign wire3496 = ( n_n41  &  wire172 ) | ( wire719  &  n_n41  &  n_n191 ) ;
 assign wire3497 = ( wire725  &  n_n40  &  n_n216 ) | ( wire721  &  n_n40  &  n_n216 ) ;
 assign wire18272 = ( wire3498 ) | ( wire18269 ) | ( n_n40  &  wire217 ) ;
 assign wire18273 = ( n_n5067 ) | ( n_n5059 ) | ( wire18270 ) ;
 assign n_n3037 = ( wire3496 ) | ( wire3497 ) | ( wire18272 ) | ( wire18273 ) ;
 assign wire469 = ( n_n177  &  wire717 ) | ( n_n177  &  wire724 ) ;
 assign wire1331 = ( wire53 ) | ( wire117 ) | ( wire281 ) | ( wire294 ) ;
 assign wire673 = ( n_n40  &  wire247 ) | ( n_n41  &  wire218 ) ;
 assign wire18283 = ( n_n6492 ) | ( n_n3413 ) | ( n_n40  &  wire1432 ) ;
 assign n_n3029 = ( n_n3037 ) | ( wire18287 ) | ( _30987 ) | ( _30988 ) ;
 assign wire1336 = ( wire157 ) | ( wire186 ) | ( wire209 ) | ( wire174 ) ;
 assign wire173 = ( wire725  &  n_n149 ) | ( n_n149  &  wire721 ) ;
 assign n_n2733 = ( n_n33  &  wire173 ) | ( wire719  &  n_n149  &  n_n33 ) ;
 assign wire1341 = ( i_15_  &  n_n216  &  n_n213 ) | ( (~ i_15_)  &  n_n216  &  n_n213 ) | ( (~ i_15_)  &  n_n216  &  n_n209 ) ;
 assign wire378 = ( n_n177  &  wire721 ) | ( n_n177  &  wire728 ) ;
 assign wire1345 = ( i_8_  &  n_n162  &  n_n16  &  n_n220 ) | ( (~ i_8_)  &  n_n162  &  n_n16  &  n_n220 ) ;
 assign wire1343 = ( wire720  &  n_n199 ) | ( wire715  &  n_n199 ) | ( wire727  &  n_n199 ) ;
 assign wire1342 = ( n_n149  &  wire721 ) | ( n_n156  &  wire728 ) | ( n_n149  &  wire728 ) ;
 assign wire165 = ( i_15_  &  n_n184  &  n_n207 ) | ( (~ i_15_)  &  n_n184  &  n_n207 ) | ( (~ i_15_)  &  n_n184  &  n_n209 ) ;
 assign wire1347 = ( wire48 ) | ( wire124 ) | ( wire167 ) | ( wire165 ) ;
 assign wire280 = ( i_15_  &  n_n177  &  n_n207 ) | ( (~ i_15_)  &  n_n177  &  n_n207 ) | ( (~ i_15_)  &  n_n177  &  n_n209 ) ;
 assign wire1346 = ( wire124 ) | ( wire167 ) | ( wire165 ) | ( wire280 ) ;
 assign wire2302 = ( n_n212  &  wire134 ) | ( n_n212  &  wire121 ) | ( n_n212  &  wire194 ) ;
 assign wire2303 = ( wire55  &  n_n197 ) | ( n_n197  &  wire280 ) | ( n_n197  &  wire121 ) ;
 assign wire19510 = ( wire132  &  n_n197 ) | ( wire132  &  n_n212 ) | ( n_n197  &  wire46 ) ;
 assign n_n784 = ( wire2302 ) | ( wire2303 ) | ( wire19510 ) ;
 assign wire629 = ( n_n218  &  n_n220  &  wire47  &  n_n200 ) ;
 assign wire2308 = ( n_n218  &  n_n220  &  n_n200  &  wire1347 ) ;
 assign wire19506 = ( n_n212  &  wire46 ) | ( n_n212  &  wire1346 ) ;
 assign wire19516 = ( wire629 ) | ( wire2295 ) | ( wire2296 ) | ( wire19513 ) ;
 assign n_n752 = ( n_n784 ) | ( wire2308 ) | ( wire19506 ) | ( wire19516 ) ;
 assign wire166 = ( wire720  &  n_n191 ) | ( wire723  &  n_n191 ) | ( wire727  &  n_n191 ) ;
 assign wire269 = ( n_n184  &  wire720 ) | ( n_n184  &  wire723 ) | ( n_n184  &  wire727 ) ;
 assign wire275 = ( i_15_  &  n_n184  &  n_n205 ) | ( (~ i_15_)  &  n_n184  &  n_n205 ) | ( (~ i_15_)  &  n_n184  &  n_n211 ) ;
 assign wire278 = ( i_15_  &  n_n205  &  n_n191 ) | ( (~ i_15_)  &  n_n205  &  n_n191 ) | ( (~ i_15_)  &  n_n211  &  n_n191 ) ;
 assign wire1354 = ( wire166 ) | ( wire269 ) | ( wire275 ) | ( wire278 ) ;
 assign wire1357 = ( i_9_  &  i_10_  &  i_11_  &  wire728 ) | ( (~ i_9_)  &  i_10_  &  i_11_  &  wire728 ) | ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire728 ) ;
 assign wire282 = ( i_15_  &  n_n205  &  n_n170 ) | ( (~ i_15_)  &  n_n205  &  n_n170 ) | ( (~ i_15_)  &  n_n211  &  n_n170 ) ;
 assign wire283 = ( n_n170  &  wire720 ) | ( n_n170  &  wire723 ) | ( n_n170  &  wire727 ) ;
 assign wire1363 = ( wire244 ) | ( wire140 ) | ( wire282 ) | ( wire283 ) ;
 assign wire296 = ( wire720  &  n_n199 ) | ( wire723  &  n_n199 ) | ( wire727  &  n_n199 ) ;
 assign wire262 = ( i_15_  &  n_n205  &  n_n216 ) | ( (~ i_15_)  &  n_n205  &  n_n216 ) | ( (~ i_15_)  &  n_n211  &  n_n216 ) ;
 assign wire332 = ( i_15_  &  n_n205  &  n_n199 ) | ( (~ i_15_)  &  n_n205  &  n_n199 ) | ( (~ i_15_)  &  n_n211  &  n_n199 ) ;
 assign wire342 = ( wire720  &  n_n216 ) | ( wire723  &  n_n216 ) | ( wire727  &  n_n216 ) ;
 assign wire1366 = ( wire296 ) | ( wire262 ) | ( wire332 ) | ( wire342 ) ;
 assign wire1367 = ( (~ i_9_)  &  i_10_  &  (~ i_11_)  &  wire725 ) | ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire725 ) ;
 assign wire479 = ( n_n125  &  wire155 ) | ( n_n125  &  wire215 ) | ( n_n125  &  n_n155 ) ;
 assign n_n3525 = ( wire137  &  n_n36 ) | ( wire146  &  n_n36 ) | ( wire131  &  n_n36 ) ;
 assign wire1375 = ( n_n220  &  n_n156  &  n_n111 ) | ( n_n220  &  n_n177  &  n_n111 ) ;
 assign n_n3561 = ( n_n47  &  wire63 ) | ( n_n47  &  wire48 ) | ( n_n47  &  wire52 ) ;
 assign n_n3578 = ( wire143  &  n_n108 ) | ( wire154  &  n_n108 ) | ( n_n108  &  wire181 ) ;
 assign wire4067 = ( wire143  &  n_n101 ) | ( wire154  &  n_n101 ) | ( wire47  &  n_n101 ) ;
 assign wire17716 = ( n_n5739 ) | ( wire440 ) | ( n_n112  &  wire160 ) ;
 assign wire17717 = ( wire447 ) | ( n_n5743 ) | ( wire47  &  n_n108 ) ;
 assign wire1378 = ( wire63 ) | ( wire48 ) | ( wire52 ) | ( wire129 ) ;
 assign wire18454 = ( wire3498 ) | ( wire18269 ) | ( n_n40  &  wire217 ) ;
 assign wire18455 = ( n_n5067 ) | ( wire673 ) | ( n_n40  &  wire172 ) ;
 assign n_n3180 = ( wire3496 ) | ( wire3497 ) | ( wire18454 ) | ( wire18455 ) ;
 assign wire1381 = ( wire132 ) | ( wire149 ) | ( wire126 ) | ( wire147 ) ;
 assign wire1383 = ( wire55 ) | ( wire127 ) | ( wire158 ) | ( wire133 ) ;
 assign wire18461 = ( n_n5075 ) | ( wire3479 ) | ( _31229 ) ;
 assign n_n3170 = ( n_n3180 ) | ( wire3275 ) | ( _31237 ) | ( _31238 ) ;
 assign wire1386 = ( wire168 ) | ( wire74 ) | ( wire68 ) | ( wire151 ) ;
 assign wire1390 = ( i_9_  &  i_10_  &  (~ i_11_)  &  wire730 ) | ( (~ i_9_)  &  i_10_  &  (~ i_11_)  &  wire730 ) ;
 assign wire1389 = ( (~ i_9_)  &  i_10_  &  (~ i_11_)  &  wire730 ) | ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire730 ) ;
 assign wire170 = ( wire729  &  n_n149 ) | ( wire730  &  n_n149 ) ;
 assign wire18534 = ( wire719  &  n_n199 ) | ( wire725  &  n_n216 ) ;
 assign wire1395 = ( wire247 ) | ( wire125 ) | ( wire160 ) | ( wire18534 ) ;
 assign wire1404 = ( n_n156  &  wire721 ) | ( n_n149  &  wire721 ) | ( n_n156  &  wire728 ) | ( n_n149  &  wire728 ) ;
 assign wire1405 = ( n_n170  &  wire721 ) | ( n_n170  &  wire728 ) | ( wire721  &  n_n191 ) | ( wire728  &  n_n191 ) ;
 assign wire2080 = ( wire154  &  n_n36 ) | ( n_n36  &  wire19714 ) ;
 assign n_n371 = ( wire712 ) | ( wire2080 ) | ( n_n34  &  n_n198 ) ;
 assign wire1416 = ( i_9_  &  (~ i_10_)  &  i_11_  &  wire728 ) | ( i_9_  &  i_10_  &  (~ i_11_)  &  wire728 ) ;
 assign wire1415 = ( i_9_  &  (~ i_10_)  &  i_11_  &  wire728 ) | ( (~ i_9_)  &  i_10_  &  (~ i_11_)  &  wire728 ) | ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire728 ) ;
 assign wire1414 = ( (~ i_9_)  &  (~ i_10_)  &  i_11_  &  wire728 ) | ( (~ i_9_)  &  (~ i_10_)  &  (~ i_11_)  &  wire728 ) ;
 assign wire759 = ( n_n220  &  n_n111  &  n_n149 ) ;
 assign wire645 = ( n_n40  &  wire155 ) | ( n_n40  &  wire205 ) ;
 assign wire664 = ( n_n41  &  wire234 ) | ( n_n41  &  wire84 ) ;
 assign wire394 = ( n_n125  &  wire224 ) | ( n_n125  &  wire250 ) | ( n_n125  &  wire57 ) ;
 assign wire240 = ( wire717  &  n_n191 ) | ( n_n191  &  wire724 ) | ( n_n191  &  wire718 ) ;
 assign wire187 = ( wire722  &  n_n191 ) | ( wire715  &  n_n191 ) | ( wire727  &  n_n191 ) ;
 assign wire210 = ( wire723  &  n_n191 ) | ( wire730  &  n_n191 ) | ( n_n191  &  wire716 ) ;
 assign wire17741 = ( i_9_  &  (~ i_10_)  &  i_11_  &  wire720 ) | ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire720 ) ;
 assign wire1420 = ( wire240 ) | ( wire187 ) | ( wire210 ) | ( wire17741 ) ;
 assign n_n3592 = ( n_n125  &  wire240 ) | ( n_n125  &  wire187 ) | ( n_n125  &  wire210 ) ;
 assign wire648 = ( wire137  &  n_n212 ) | ( n_n212  &  wire46 ) ;
 assign wire681 = ( n_n197  &  wire63 ) | ( n_n197  &  wire48 ) ;
 assign wire17766 = ( n_n197  &  wire52 ) | ( n_n197  &  wire129 ) ;
 assign wire17767 = ( n_n212  &  wire63 ) | ( n_n212  &  wire52 ) | ( n_n212  &  wire129 ) ;
 assign n_n3834 = ( wire648 ) | ( wire681 ) | ( wire17766 ) | ( wire17767 ) ;
 assign n_n3601 = ( n_n212  &  wire134 ) | ( n_n212  &  wire156 ) | ( n_n212  &  wire123 ) ;
 assign wire504 = ( wire146  &  n_n212 ) | ( wire131  &  n_n212 ) ;
 assign n_n3833 = ( n_n2770 ) | ( n_n4692 ) | ( n_n3601 ) | ( wire504 ) ;
 assign wire1425 = ( n_n51 ) | ( wire245 ) | ( wire144 ) | ( wire122 ) ;
 assign wire1427 = ( n_n159  &  n_n35  &  n_n48 ) | ( n_n159  &  n_n124  &  n_n48 ) ;
 assign wire1432 = ( n_n65 ) | ( wire115 ) | ( wire221 ) | ( wire298 ) ;
 assign wire19099 = ( n_n156  &  wire727 ) | ( n_n156  &  wire717 ) ;
 assign wire1436 = ( wire90 ) | ( wire198 ) | ( wire175 ) | ( wire19099 ) ;
 assign wire1437 = ( wire48 ) | ( wire124 ) | ( wire167 ) | ( wire165 ) ;
 assign wire19599 = ( n_n47  &  wire48 ) | ( n_n47  &  wire124 ) ;
 assign wire19600 = ( n_n47  &  wire46 ) | ( n_n47  &  wire167 ) | ( n_n47  &  wire165 ) ;
 assign n_n772 = ( wire19599 ) | ( wire19600 ) | ( n_n46  &  wire1437 ) ;
 assign wire235 = ( i_15_  &  n_n205  &  n_n149 ) | ( (~ i_15_)  &  n_n205  &  n_n149 ) | ( (~ i_15_)  &  n_n211  &  n_n149 ) ;
 assign wire236 = ( wire720  &  n_n149 ) | ( wire723  &  n_n149 ) | ( wire727  &  n_n149 ) ;
 assign wire1444 = ( wire166 ) | ( wire269 ) | ( wire275 ) | ( wire278 ) ;
 assign wire325 = ( n_n177  &  wire720 ) | ( n_n177  &  wire723 ) | ( n_n177  &  wire727 ) ;
 assign n_n326 = ( n_n47  &  wire1444 ) | ( n_n46  &  wire1444 ) | ( n_n47  &  wire325 ) ;
 assign wire19701 = ( n_n156  &  wire730 ) | ( n_n156  &  wire718 ) ;
 assign wire1446 = ( wire244 ) | ( wire235 ) | ( wire236 ) | ( wire19701 ) ;
 assign wire497 = ( n_n41  &  n_n190 ) | ( n_n41  &  wire187 ) | ( n_n41  &  wire210 ) ;
 assign wire1450 = ( n_n190 ) | ( wire240 ) | ( wire187 ) | ( wire210 ) ;
 assign wire636 = ( wire157  &  n_n36 ) | ( n_n34  &  wire174 ) ;
 assign wire18253 = ( wire729  &  n_n177 ) | ( n_n177  &  wire720 ) | ( n_n177  &  wire715 ) ;
 assign wire1459 = ( wire120 ) | ( wire179 ) | ( wire324 ) | ( wire18253 ) ;
 assign wire1463 = ( (~ i_7_)  &  i_6_ ) | ( (~ i_7_)  &  (~ i_6_) ) ;
 assign wire4223 = ( n_n162  &  n_n19  &  wire1463 ) | ( n_n48  &  n_n19  &  wire1463 ) ;
 assign wire17588 = ( (~ i_7_)  &  i_6_  &  n_n19  &  n_n111 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n19  &  n_n111 ) ;
 assign n_n2956 = ( n_n7254 ) | ( wire551 ) | ( wire4223 ) | ( wire17588 ) ;
 assign wire1465 = ( wire134 ) | ( wire156 ) | ( wire176 ) | ( wire123 ) ;
 assign wire1470 = ( i_9_  &  (~ i_10_)  &  i_11_  &  wire721 ) | ( (~ i_9_)  &  (~ i_10_)  &  i_11_  &  wire721 ) | ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire721 ) ;
 assign wire1469 = ( i_9_  &  (~ i_10_)  &  i_11_  &  wire721 ) | ( (~ i_9_)  &  (~ i_10_)  &  i_11_  &  wire721 ) | ( i_9_  &  i_10_  &  (~ i_11_)  &  wire721 ) | ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire721 ) ;
 assign wire401 = ( (~ i_9_)  &  i_10_  &  i_11_  &  wire719 ) | ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire719 ) ;
 assign wire1477 = ( i_9_  &  i_10_  &  i_11_  &  wire728 ) | ( i_9_  &  (~ i_10_)  &  i_11_  &  wire728 ) | ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire728 ) | ( (~ i_9_)  &  (~ i_10_)  &  (~ i_11_)  &  wire728 ) ;
 assign wire1476 = ( i_9_  &  i_10_  &  i_11_  &  wire728 ) | ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire728 ) | ( (~ i_9_)  &  (~ i_10_)  &  (~ i_11_)  &  wire728 ) ;
 assign wire1480 = ( i_8_  &  n_n17  &  n_n48  &  n_n220 ) | ( (~ i_8_)  &  n_n17  &  n_n48  &  n_n220 ) ;
 assign wire1479 = ( n_n177  &  wire720 ) | ( n_n170  &  wire720 ) | ( n_n177  &  wire727 ) | ( n_n170  &  wire727 ) ;
 assign wire1478 = ( (~ i_9_)  &  (~ i_10_)  &  i_11_  &  wire728 ) | ( (~ i_9_)  &  i_10_  &  (~ i_11_)  &  wire728 ) ;
 assign wire336 = ( n_n177  &  wire723 ) | ( n_n177  &  wire730 ) | ( n_n177  &  wire718 ) ;
 assign wire19895 = ( n_n177  &  wire720 ) | ( n_n177  &  wire727 ) | ( n_n177  &  wire726 ) ;
 assign wire1483 = ( wire110 ) | ( n_n164 ) | ( wire336 ) | ( wire19895 ) ;
 assign wire161 = ( n_n170  &  wire720 ) | ( n_n170  &  wire727 ) ;
 assign wire1482 = ( n_n185 ) | ( wire336 ) | ( wire19895 ) | ( wire161 ) ;
 assign wire16886 = ( n_n3276 ) | ( wire462 ) | ( wire16884 ) | ( wire16885 ) ;
 assign n_n5021 = ( n_n101  &  wire86 ) | ( n_n108  &  n_n190 ) ;
 assign wire565 = ( n_n197  &  wire134 ) | ( n_n197  &  wire156 ) ;
 assign wire1488 = ( _30471 ) | ( n_n156  &  wire719 ) | ( n_n156  &  wire728 ) ;
 assign wire579 = ( n_n212  &  wire52 ) | ( n_n212  &  wire129 ) ;
 assign wire1489 = ( wire137 ) | ( wire146 ) | ( wire46 ) ;
 assign wire3985 = ( n_n30  &  wire134 ) | ( n_n30  &  wire156 ) ;
 assign wire17787 = ( n_n30  &  wire131 ) | ( n_n30  &  wire176 ) | ( n_n30  &  wire123 ) ;
 assign n_n3514 = ( n_n31  &  wire63 ) | ( n_n31  &  wire48 ) | ( n_n31  &  wire52 ) ;
 assign wire1491 = ( wire143 ) | ( wire154 ) | ( wire63 ) | ( wire48 ) ;
 assign wire17793 = ( n_n30  &  wire181 ) | ( n_n31  &  wire129 ) ;
 assign n_n3511 = ( n_n31  &  wire137 ) | ( n_n31  &  wire146 ) | ( n_n31  &  wire131 ) ;
 assign wire690 = ( n_n30  &  wire137 ) | ( n_n30  &  wire46 ) ;
 assign wire1493 = ( wire63 ) | ( wire48 ) | ( wire52 ) | ( wire129 ) ;
 assign wire1496 = ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire725 ) | ( (~ i_9_)  &  (~ i_10_)  &  (~ i_11_)  &  wire725 ) ;
 assign wire230 = ( n_n170  &  wire723 ) | ( n_n170  &  wire716 ) | ( n_n170  &  wire718 ) ;
 assign wire1498 = ( n_n82 ) | ( wire260 ) | ( wire373 ) | ( wire230 ) ;
 assign wire347 = ( wire723  &  n_n149 ) | ( n_n149  &  wire716 ) | ( n_n149  &  wire718 ) ;
 assign wire352 = ( wire729  &  n_n170 ) | ( n_n170  &  wire717 ) ;
 assign wire1497 = ( n_n70 ) | ( wire230 ) | ( wire347 ) | ( wire352 ) ;
 assign wire1500 = ( n_n156  &  wire721 ) | ( n_n149  &  wire721 ) | ( n_n156  &  wire728 ) | ( n_n149  &  wire728 ) ;
 assign wire1499 = ( n_n156  &  wire721 ) | ( n_n149  &  wire721 ) | ( n_n156  &  wire728 ) | ( n_n149  &  wire728 ) ;
 assign wire1503 = ( n_n177  &  wire721 ) | ( n_n170  &  wire721 ) | ( n_n177  &  wire728 ) | ( n_n170  &  wire728 ) ;
 assign wire1504 = ( wire127 ) | ( wire133 ) | ( wire60 ) | ( wire227 ) ;
 assign wire357 = ( wire720  &  n_n191 ) | ( wire715  &  n_n191 ) | ( wire727  &  n_n191 ) ;
 assign wire19328 = ( i_15_  &  n_n170  &  n_n213 ) | ( (~ i_15_)  &  n_n170  &  n_n213 ) | ( (~ i_15_)  &  n_n170  &  n_n209 ) ;
 assign wire1507 = ( wire349 ) | ( wire210 ) | ( wire357 ) | ( wire19328 ) ;
 assign wire314 = ( n_n184  &  wire723 ) | ( n_n184  &  wire730 ) | ( n_n184  &  wire718 ) ;
 assign wire1510 = ( wire314 ) | ( n_n184  &  wire726 ) ;
 assign wire259 = ( n_n177  &  wire720 ) | ( n_n177  &  wire727 ) ;
 assign wire337 = ( wire723  &  n_n191 ) | ( wire730  &  n_n191 ) | ( n_n191  &  wire718 ) ;
 assign wire19831 = ( wire720  &  n_n191 ) | ( wire727  &  n_n191 ) | ( n_n191  &  wire726 ) ;
 assign wire1513 = ( n_n178 ) | ( wire259 ) | ( wire337 ) | ( wire19831 ) ;
 assign wire338 = ( n_n184  &  wire720 ) | ( n_n184  &  wire727 ) ;
 assign wire1512 = ( n_n202 ) | ( wire337 ) | ( wire19831 ) | ( wire338 ) ;
 assign wire689 = ( wire157  &  n_n212 ) | ( n_n197  &  wire174 ) ;
 assign wire1519 = ( wire172 ) | ( wire51 ) | ( wire240 ) | ( wire210 ) ;
 assign wire1520 = ( wire130 ) | ( wire139 ) | ( wire124 ) | ( wire128 ) ;
 assign wire370 = ( wire729  &  n_n156 ) | ( n_n156  &  wire730 ) ;
 assign wire18367 = ( n_n7346 ) | ( n_n5319 ) | ( wire185  &  n_n3 ) ;
 assign n_n3176 = ( wire707 ) | ( wire18367 ) | ( _3127 ) ;
 assign wire1524 = ( i_5_  &  (~ i_3_)  &  i_4_  &  n_n19 ) | ( (~ i_5_)  &  (~ i_3_)  &  i_4_  &  n_n19 ) | ( i_5_  &  (~ i_3_)  &  (~ i_4_)  &  n_n19 ) | ( (~ i_5_)  &  (~ i_3_)  &  (~ i_4_)  &  n_n19 ) ;
 assign wire1527 = ( n_n159  &  n_n218  &  n_n35 ) | ( n_n159  &  n_n218  &  n_n124 ) ;
 assign wire315 = ( wire729  &  n_n149 ) | ( wire717  &  n_n149 ) | ( n_n149  &  wire726 ) ;
 assign wire1537 = ( n_n184  &  wire721 ) | ( n_n177  &  wire721 ) | ( n_n184  &  wire728 ) | ( n_n177  &  wire728 ) ;
 assign wire19442 = ( wire729  &  n_n156 ) | ( n_n184  &  wire728 ) ;
 assign wire19443 = ( wire721  &  n_n199 ) | ( wire728  &  n_n199 ) | ( wire721  &  n_n216 ) | ( wire728  &  n_n216 ) ;
 assign wire1539 = ( wire155 ) | ( wire232 ) | ( wire19442 ) | ( wire19443 ) ;
 assign n_n1163 = ( wire2359 ) | ( _32495 ) | ( n_n30  &  wire1539 ) ;
 assign wire348 = ( i_15_  &  n_n205  &  n_n191 ) | ( (~ i_15_)  &  n_n205  &  n_n191 ) ;
 assign wire1544 = ( wire137 ) | ( wire146 ) | ( n_n84 ) | ( wire46 ) ;
 assign wire1553 = ( wire721  &  n_n199 ) | ( wire728  &  n_n199 ) | ( wire721  &  n_n216 ) | ( wire728  &  n_n216 ) ;
 assign wire1556 = ( n_n177  &  wire721 ) | ( n_n170  &  wire721 ) | ( n_n177  &  wire728 ) | ( n_n170  &  wire728 ) ;
 assign wire1558 = ( n_n184  &  wire721 ) | ( n_n177  &  wire721 ) | ( n_n184  &  wire728 ) | ( n_n177  &  wire728 ) ;
 assign wire1560 = ( wire721  &  n_n191 ) | ( wire728  &  n_n191 ) | ( wire721  &  n_n199 ) | ( wire728  &  n_n199 ) ;
 assign wire1562 = ( n_n184  &  wire721 ) | ( n_n184  &  wire728 ) | ( wire721  &  n_n191 ) | ( wire728  &  n_n191 ) ;
 assign wire295 = ( wire723  &  n_n199 ) | ( wire730  &  n_n199 ) | ( n_n199  &  wire718 ) ;
 assign wire333 = ( wire723  &  n_n216 ) | ( wire730  &  n_n216 ) | ( n_n216  &  wire718 ) ;
 assign wire19882 = ( wire720  &  n_n199 ) | ( wire727  &  n_n199 ) | ( n_n199  &  wire726 ) ;
 assign wire1568 = ( n_n202 ) | ( wire295 ) | ( wire333 ) | ( wire19882 ) ;
 assign wire1570 = ( i_15_  &  n_n156  &  n_n205 ) | ( (~ i_15_)  &  n_n156  &  n_n205 ) | ( i_15_  &  n_n156  &  n_n215 ) ;
 assign wire560 = ( n_n47  &  wire176 ) | ( n_n47  &  wire123 ) ;
 assign wire688 = ( n_n46  &  wire156 ) | ( n_n46  &  wire123 ) ;
 assign wire289 = ( n_n156  &  wire722 ) | ( n_n156  &  wire723 ) | ( n_n156  &  wire727 ) ;
 assign wire18426 = ( wire729  &  n_n156 ) | ( n_n156  &  wire720 ) | ( n_n156  &  wire715 ) ;
 assign wire1576 = ( wire116 ) | ( wire198 ) | ( wire289 ) | ( wire18426 ) ;
 assign n_n3555 = ( n_n47  &  wire127 ) | ( n_n47  &  wire158 ) | ( n_n47  &  wire133 ) ;
 assign wire1580 = ( (~ i_9_)  &  i_10_  &  i_11_  &  wire721 ) | ( i_9_  &  (~ i_10_)  &  i_11_  &  wire721 ) | ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire721 ) ;
 assign wire1579 = ( i_9_  &  i_10_  &  i_11_  &  wire721 ) | ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire721 ) ;
 assign wire1578 = ( (~ i_9_)  &  (~ i_10_)  &  i_11_  &  wire721 ) | ( (~ i_9_)  &  (~ i_10_)  &  (~ i_11_)  &  wire721 ) ;
 assign wire19318 = ( wire729  &  n_n199 ) | ( wire717  &  n_n199 ) ;
 assign wire1581 = ( wire108 ) | ( wire385 ) | ( wire19318 ) ;
 assign wire1582 = ( n_n184  &  wire721 ) | ( n_n184  &  wire728 ) | ( wire721  &  n_n191 ) | ( wire728  &  n_n191 ) ;
 assign wire19835 = ( wire720  &  n_n199 ) | ( wire727  &  n_n199 ) | ( n_n199  &  wire726 ) ;
 assign wire1587 = ( wire335 ) | ( wire295 ) | ( wire333 ) | ( wire19835 ) ;
 assign wire19901 = ( i_9_  &  i_10_  &  i_11_  &  wire726 ) | ( (~ i_9_)  &  (~ i_10_)  &  (~ i_11_)  &  wire726 ) ;
 assign wire1590 = ( wire314 ) | ( wire338 ) | ( wire333 ) | ( wire19901 ) ;
 assign wire19905 = ( wire720  &  n_n149 ) | ( wire727  &  n_n149 ) | ( n_n149  &  wire726 ) ;
 assign wire1592 = ( n_n150 ) | ( wire248 ) | ( wire249 ) | ( wire19905 ) ;
 assign wire121 = ( i_15_  &  n_n170  &  n_n207 ) | ( (~ i_15_)  &  n_n170  &  n_n207 ) | ( (~ i_15_)  &  n_n170  &  n_n209 ) ;
 assign wire434 = ( n_n39  &  n_n156  &  wire728 ) | ( n_n39  &  n_n149  &  wire728 ) ;
 assign wire538 = ( n_n125  &  wire108 ) | ( n_n125  &  wire258 ) ;
 assign wire539 = ( n_n125  &  wire86 ) | ( n_n125  &  wire180 ) ;
 assign wire17918 = ( wire152 ) | ( wire150 ) ;
 assign wire17919 = ( wire153 ) | ( wire217 ) | ( wire719  &  n_n191 ) ;
 assign wire17920 = ( wire80 ) | ( wire78 ) | ( _30833 ) ;
 assign wire17921 = ( wire157 ) | ( n_n63 ) | ( wire135 ) | ( wire17916 ) ;
 assign wire1601 = ( wire17918 ) | ( wire17919 ) | ( wire17920 ) | ( wire17921 ) ;
 assign n_n2777 = ( n_n212  &  wire139 ) | ( n_n212  &  wire124 ) | ( n_n212  &  wire128 ) ;
 assign wire1602 = ( wire130 ) | ( wire139 ) | ( wire124 ) | ( wire128 ) ;
 assign wire607 = ( wire146  &  n_n34 ) | ( wire131  &  n_n34 ) ;
 assign wire640 = ( n_n34  &  wire63 ) | ( n_n34  &  wire48 ) ;
 assign wire584 = ( wire132  &  n_n36 ) | ( n_n36  &  wire126 ) ;
 assign wire107 = ( n_n184  &  wire722 ) | ( n_n184  &  wire715 ) | ( n_n184  &  wire727 ) ;
 assign wire339 = ( i_15_  &  n_n191  &  n_n207 ) | ( (~ i_15_)  &  n_n191  &  n_n207 ) ;
 assign wire19523 = ( i_15_  &  n_n184  &  n_n207 ) | ( (~ i_15_)  &  n_n184  &  n_n207 ) | ( i_15_  &  n_n184  &  n_n215 ) ;
 assign wire1605 = ( wire187 ) | ( wire107 ) | ( wire339 ) | ( wire19523 ) ;
 assign wire19767 = ( wire720  &  n_n199 ) | ( wire727  &  n_n199 ) | ( n_n199  &  wire726 ) ;
 assign wire1613 = ( wire335 ) | ( wire295 ) | ( wire333 ) | ( wire19767 ) ;
 assign wire99 = ( n_n177  &  wire730 ) | ( n_n177  &  wire718 ) ;
 assign wire1617 = ( wire282 ) | ( wire283 ) | ( wire325 ) | ( wire99 ) ;
 assign wire18028 = ( n_n47  &  wire149 ) | ( n_n47  &  wire147 ) ;
 assign n_n3485 = ( wire674 ) | ( n_n3889 ) | ( wire686 ) | ( wire18028 ) ;
 assign wire698 = ( n_n125  &  wire208 ) | ( n_n125  &  wire148 ) ;
 assign wire3820 = ( n_n31  &  wire55 ) | ( n_n31  &  wire127 ) | ( n_n31  &  wire133 ) ;
 assign wire17926 = ( n_n31  &  wire149 ) | ( n_n31  &  wire158 ) ;
 assign n_n3510 = ( n_n31  &  wire132 ) | ( n_n31  &  wire126 ) | ( n_n31  &  wire147 ) ;
 assign wire1625 = ( wire130 ) | ( wire139 ) | ( wire124 ) | ( wire128 ) ;
 assign wire578 = ( wire126  &  n_n197 ) | ( wire147  &  n_n197 ) ;
 assign wire3177 = ( wire126  &  n_n212 ) | ( wire147  &  n_n212 ) ;
 assign wire18581 = ( wire149  &  n_n197 ) | ( wire132  &  n_n212 ) ;
 assign wire18582 = ( wire132  &  n_n197 ) | ( wire149  &  n_n212 ) ;
 assign wire18583 = ( wire126  &  n_n197 ) | ( wire147  &  n_n197 ) | ( n_n197  &  wire46 ) ;
 assign wire1627 = ( wire130 ) | ( wire139 ) | ( wire124 ) | ( wire128 ) ;
 assign wire17880 = ( n_n36  &  wire52 ) | ( n_n36  &  wire129 ) ;
 assign wire17881 = ( n_n36  &  wire139 ) | ( n_n36  &  wire124 ) | ( n_n36  &  wire128 ) ;
 assign wire642 = ( n_n36  &  wire63 ) | ( n_n36  &  wire48 ) ;
 assign wire322 = ( i_15_  &  n_n216  &  n_n207 ) | ( (~ i_15_)  &  n_n216  &  n_n207 ) | ( (~ i_15_)  &  n_n216  &  n_n209 ) ;
 assign wire1628 = ( wire47 ) | ( wire124 ) | ( wire165 ) | ( wire322 ) ;
 assign wire407 = ( i_9_  &  i_10_  &  i_11_  &  wire719 ) | ( (~ i_9_)  &  (~ i_10_)  &  (~ i_11_)  &  wire719 ) ;
 assign wire1630 = ( i_9_  &  (~ i_10_)  &  i_11_  &  wire719 ) | ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire719 ) | ( (~ i_9_)  &  (~ i_10_)  &  (~ i_11_)  &  wire719 ) ;
 assign wire163 = ( i_15_  &  n_n149  &  n_n207 ) | ( (~ i_15_)  &  n_n149  &  n_n207 ) | ( (~ i_15_)  &  n_n149  &  n_n209 ) ;
 assign wire194 = ( i_15_  &  n_n156  &  n_n207 ) | ( (~ i_15_)  &  n_n156  &  n_n207 ) | ( (~ i_15_)  &  n_n156  &  n_n209 ) ;
 assign wire1632 = ( wire55 ) | ( wire134 ) | ( wire163 ) | ( wire194 ) ;
 assign n_n765 = ( n_n40  &  wire280 ) | ( n_n41  &  wire1632 ) | ( n_n40  &  wire1632 ) ;
 assign wire635 = ( n_n39  &  n_n134 ) | ( n_n38  &  n_n132 ) ;
 assign wire1633 = ( wire720  &  n_n149 ) | ( wire727  &  n_n149 ) ;
 assign wire19556 = ( wire635 ) | ( wire19552 ) | ( n_n39  &  wire1633 ) ;
 assign wire19557 = ( n_n969 ) | ( n_n972 ) | ( _32772 ) ;
 assign wire19560 = ( n_n765 ) | ( wire19548 ) | ( wire19549 ) ;
 assign wire346 = ( i_15_  &  n_n184  &  n_n205 ) | ( (~ i_15_)  &  n_n184  &  n_n205 ) ;
 assign wire19796 = ( i_9_  &  i_10_  &  i_11_  &  wire728 ) | ( i_9_  &  (~ i_10_)  &  i_11_  &  wire728 ) | ( (~ i_9_)  &  (~ i_10_)  &  (~ i_11_)  &  wire728 ) ;
 assign wire1636 = ( n_n60 ) | ( wire235 ) | ( wire236 ) | ( wire19796 ) ;
 assign wire1640 = ( wire296 ) | ( wire262 ) | ( wire332 ) | ( wire342 ) ;
 assign wire1639 = ( i_8_  &  n_n48  &  n_n220  &  n_n18 ) | ( (~ i_8_)  &  n_n48  &  n_n220  &  n_n18 ) ;
 assign wire19786 = ( wire419 ) | ( wire2027 ) | ( wire228  &  n_n56 ) ;
 assign wire19787 = ( wire2026 ) | ( wire2032 ) | ( wire19779 ) ;
 assign wire19793 = ( wire19792 ) | ( wire1640  &  wire1639 ) ;
 assign n_n302 = ( n_n326 ) | ( wire19786 ) | ( wire19787 ) | ( wire19793 ) ;
 assign wire354 = ( i_15_  &  n_n205  &  n_n177 ) | ( (~ i_15_)  &  n_n205  &  n_n177 ) | ( (~ i_15_)  &  n_n211  &  n_n177 ) ;
 assign wire1641 = ( wire282 ) | ( wire283 ) | ( wire325 ) | ( wire354 ) ;
 assign wire19799 = ( n_n62  &  wire189 ) | ( n_n47  &  wire1636 ) ;
 assign wire19812 = ( wire1999 ) | ( wire2000 ) | ( wire19807 ) | ( wire19808 ) ;
 assign wire17960 = ( n_n36  &  wire149 ) | ( n_n36  &  wire147 ) ;
 assign wire242 = ( n_n184  &  wire725 ) | ( n_n184  &  wire721 ) | ( n_n184  &  wire728 ) ;
 assign wire272 = ( n_n184  &  wire717 ) | ( n_n184  &  wire724 ) | ( n_n184  &  wire718 ) ;
 assign wire17944 = ( n_n184  &  wire729 ) | ( n_n184  &  wire719 ) | ( n_n184  &  wire726 ) ;
 assign wire1648 = ( wire211 ) | ( wire242 ) | ( wire272 ) | ( wire17944 ) ;
 assign wire17947 = ( n_n31  &  wire143 ) | ( n_n31  &  wire181 ) ;
 assign wire17948 = ( n_n31  &  wire154 ) | ( n_n31  &  wire47 ) | ( n_n31  &  wire151 ) ;
 assign n_n3470 = ( wire17947 ) | ( wire17948 ) | ( n_n32  &  wire1648 ) ;
 assign n_n2642 = ( n_n36  &  wire127 ) | ( n_n36  &  wire158 ) | ( n_n36  &  wire133 ) ;
 assign wire18611 = ( n_n184  &  wire725 ) | ( n_n177  &  wire719 ) ;
 assign wire1655 = ( wire217 ) | ( wire209 ) | ( wire174 ) | ( wire18611 ) ;
 assign wire1658 = ( i_8_  &  n_n162  &  n_n220  &  n_n18 ) | ( (~ i_8_)  &  n_n162  &  n_n220  &  n_n18 ) ;
 assign wire2232 = ( n_n40  &  wire151 ) | ( n_n40  &  wire192 ) ;
 assign wire19569 = ( wire391 ) | ( wire19567 ) | ( n_n116  &  wire1658 ) ;
 assign wire1659 = ( wire132 ) | ( wire46 ) | ( wire280 ) | ( wire121 ) ;
 assign wire19574 = ( _1018 ) | ( _32841 ) | ( n_n41  &  wire1659 ) ;
 assign wire1668 = ( i_8_  &  n_n48  &  n_n220  &  n_n18 ) | ( (~ i_8_)  &  n_n48  &  n_n220  &  n_n18 ) ;
 assign wire1666 = ( (~ i_9_)  &  (~ i_10_)  &  i_11_  &  wire728 ) | ( (~ i_9_)  &  i_10_  &  (~ i_11_)  &  wire728 ) ;
 assign wire19846 = ( wire1951 ) | ( n_n113  &  wire128 ) | ( n_n113  &  wire19843 ) ;
 assign wire18122 = ( n_n212  &  wire63 ) | ( n_n212  &  wire130 ) ;
 assign n_n3501 = ( wire648 ) | ( wire579 ) | ( n_n2777 ) | ( wire18122 ) ;
 assign wire18125 = ( wire132  &  n_n212 ) | ( wire149  &  n_n212 ) ;
 assign n_n3500 = ( wire557 ) | ( n_n3601 ) | ( wire504 ) | ( wire18125 ) ;
 assign wire19577 = ( i_9_  &  i_10_  &  i_11_  &  wire719 ) | ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire719 ) | ( (~ i_9_)  &  (~ i_10_)  &  (~ i_11_)  &  wire719 ) ;
 assign wire1674 = ( wire55 ) | ( wire163 ) | ( wire194 ) | ( wire19577 ) ;
 assign wire2218 = ( n_n43  &  wire187 ) | ( n_n43  &  wire339 ) ;
 assign wire19584 = ( n_n6271 ) | ( n_n6270 ) | ( n_n42  &  n_n183 ) ;
 assign n_n834 = ( wire2218 ) | ( wire19584 ) | ( n_n43  &  n_n190 ) ;
 assign wire1675 = ( (~ i_9_)  &  (~ i_10_)  &  i_11_  &  wire719 ) | ( (~ i_9_)  &  i_10_  &  (~ i_11_)  &  wire719 ) ;
 assign wire19587 = ( n_n134  &  n_n46 ) | ( n_n43  &  n_n183 ) ;
 assign wire19588 = ( n_n47  &  n_n130 ) | ( n_n46  &  n_n130 ) | ( n_n47  &  wire1675 ) | ( n_n46  &  wire1675 ) ;
 assign wire19591 = ( wire19589 ) | ( n_n42  &  wire107 ) | ( n_n42  &  wire340 ) ;
 assign wire19582 = ( wire19580 ) | ( n_n47  &  wire163 ) | ( n_n47  &  wire19576 ) ;
 assign wire19596 = ( wire2205 ) | ( _969 ) | ( _976 ) | ( _32877 ) ;
 assign wire415 = ( wire730  &  n_n216 ) | ( n_n216  &  wire718 ) ;
 assign wire1684 = ( wire269 ) | ( wire275 ) | ( wire342 ) | ( wire415 ) ;
 assign wire1689 = ( wire51 ) | ( wire240 ) | ( wire187 ) | ( wire210 ) ;
 assign wire696 = ( n_n41  &  wire224 ) | ( n_n41  &  wire250 ) ;
 assign n_n3542 = ( n_n41  &  wire224 ) | ( n_n41  &  wire250 ) | ( n_n41  &  wire100 ) ;
 assign wire3767 = ( n_n43  &  wire130 ) | ( n_n43  &  wire222 ) ;
 assign wire17979 = ( n_n43  &  wire52 ) | ( n_n43  &  wire139 ) ;
 assign wire17980 = ( n_n43  &  wire63 ) | ( n_n43  &  wire48 ) | ( n_n43  &  wire129 ) ;
 assign n_n3482 = ( wire683 ) | ( wire3767 ) | ( wire17979 ) | ( wire17980 ) ;
 assign wire18032 = ( wire419 ) | ( wire3710 ) | ( n_n47  &  wire151 ) ;
 assign n_n3487 = ( n_n3562 ) | ( wire481 ) | ( wire577 ) | ( wire18032 ) ;
 assign wire18039 = ( n_n3561 ) | ( wire3702 ) | ( wire18035 ) | ( wire18036 ) ;
 assign n_n3460 = ( n_n3485 ) | ( n_n3487 ) | ( wire18039 ) ;
 assign wire1695 = ( wire143 ) | ( wire154 ) | ( wire47 ) | ( wire181 ) ;
 assign wire1704 = ( i_8_  &  n_n17  &  n_n48  &  n_n220 ) | ( (~ i_8_)  &  n_n17  &  n_n48  &  n_n220 ) ;
 assign wire19624 = ( wire720  &  n_n191 ) | ( wire715  &  n_n191 ) | ( n_n191  &  wire724 ) ;
 assign wire1706 = ( wire320 ) | ( wire19624 ) ;
 assign wire1709 = ( i_9_  &  i_10_  &  i_11_  &  wire719 ) | ( (~ i_9_)  &  (~ i_10_)  &  i_11_  &  wire719 ) | ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire719 ) ;
 assign wire1708 = ( i_9_  &  (~ i_10_)  &  i_11_  &  wire719 ) | ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire719 ) ;
 assign wire1707 = ( (~ i_9_)  &  i_10_  &  i_11_  &  wire719 ) | ( (~ i_9_)  &  (~ i_10_)  &  (~ i_11_)  &  wire719 ) ;
 assign wire2182 = ( n_n46  &  wire322 ) | ( n_n46  &  wire192 ) ;
 assign wire19614 = ( wire47  &  n_n46 ) | ( n_n47  &  wire151 ) ;
 assign wire19617 = ( wire2181 ) | ( wire19613 ) | ( n_n46  &  wire151 ) ;
 assign wire19619 = ( n_n772 ) | ( wire2191 ) | ( wire19610 ) | ( wire19612 ) ;
 assign wire1717 = ( i_9_  &  (~ i_10_)  &  i_11_  &  wire728 ) | ( i_9_  &  i_10_  &  (~ i_11_)  &  wire728 ) | ( (~ i_9_)  &  i_10_  &  (~ i_11_)  &  wire728 ) ;
 assign wire1716 = ( i_9_  &  (~ i_10_)  &  i_11_  &  wire728 ) | ( i_9_  &  i_10_  &  (~ i_11_)  &  wire728 ) | ( (~ i_9_)  &  i_10_  &  (~ i_11_)  &  wire728 ) ;
 assign wire1720 = ( i_15_  &  n_n205  &  n_n191 ) | ( (~ i_15_)  &  n_n205  &  n_n191 ) | ( i_15_  &  n_n191  &  n_n215 ) | ( (~ i_15_)  &  n_n191  &  n_n215 ) ;
 assign wire18657 = ( n_n184  &  wire729 ) | ( n_n184  &  wire720 ) | ( n_n184  &  wire726 ) ;
 assign wire1723 = ( wire211 ) | ( wire107 ) | ( wire272 ) | ( wire18657 ) ;
 assign wire606 = ( wire137  &  n_n34 ) | ( n_n34  &  wire46 ) ;
 assign wire1729 = ( wire130 ) | ( wire139 ) | ( wire124 ) | ( wire128 ) ;
 assign wire17896 = ( n_n34  &  wire133 ) | ( n_n34  &  wire134 ) ;
 assign wire17897 = ( n_n34  &  wire156 ) | ( n_n34  &  wire123 ) ;
 assign wire17898 = ( n_n36  &  wire55 ) | ( n_n34  &  wire158 ) ;
 assign n_n2626 = ( n_n2642 ) | ( wire17896 ) | ( wire17897 ) | ( wire17898 ) ;
 assign wire19013 = ( wire729  &  n_n199 ) | ( wire715  &  n_n199 ) | ( wire717  &  n_n199 ) ;
 assign wire1735 = ( wire261 ) | ( wire264 ) | ( wire375 ) | ( wire19013 ) ;
 assign wire1739 = ( wire132 ) | ( wire55 ) | ( wire121 ) | ( wire163 ) ;
 assign wire1738 = ( (~ i_9_)  &  (~ i_10_)  &  i_11_  &  wire719 ) | ( i_9_  &  i_10_  &  (~ i_11_)  &  wire719 ) ;
 assign wire1741 = ( n_n84 ) | ( wire279 ) | ( wire54 ) | ( wire195 ) ;
 assign wire237 = ( n_n170  &  wire722 ) | ( n_n170  &  wire727 ) | ( n_n170  &  wire716 ) ;
 assign wire1740 = ( wire53 ) | ( n_n118 ) | ( wire195 ) | ( wire237 ) ;
 assign wire19633 = ( i_9_  &  (~ i_10_)  &  i_11_  &  wire724 ) | ( (~ i_9_)  &  i_10_  &  (~ i_11_)  &  wire724 ) ;
 assign wire1743 = ( wire118 ) | ( wire199 ) | ( wire279 ) | ( wire19633 ) ;
 assign wire1742 = ( wire118 ) | ( wire290 ) | ( n_n72 ) | ( wire59 ) ;
 assign wire1949 = ( n_n123  &  wire248 ) | ( n_n123  &  wire110 ) ;
 assign wire1748 = ( wire47 ) | ( wire74 ) | ( wire68 ) | ( wire151 ) ;
 assign wire1747 = ( (~ i_9_)  &  i_10_  &  i_11_ ) | ( (~ i_9_)  &  (~ i_10_)  &  i_11_ ) | ( (~ i_9_)  &  i_10_  &  (~ i_11_) ) | ( (~ i_9_)  &  (~ i_10_)  &  (~ i_11_) ) ;
 assign wire18044 = ( wire3696 ) | ( n_n113  &  wire256 ) ;
 assign n_n3492 = ( n_n3578 ) | ( wire18044 ) | ( n_n108  &  wire1748 ) ;
 assign wire18049 = ( wire48 ) | ( wire124 ) ;
 assign wire18050 = ( wire168 ) | ( wire52 ) | ( wire128 ) ;
 assign wire18051 = ( wire63 ) | ( wire129 ) | ( wire130 ) | ( wire139 ) ;
 assign n_n3491 = ( n_n108  &  wire18049 ) | ( n_n108  &  wire18050 ) | ( n_n108  &  wire18051 ) ;
 assign wire1751 = ( wire381 ) | ( n_n130 ) | ( wire186 ) | ( wire209 ) ;
 assign wire18057 = ( wire3700 ) | ( wire3701 ) | ( n_n57  &  n_n125 ) ;
 assign wire18058 = ( wire3690 ) | ( n_n125  &  wire1751 ) ;
 assign n_n3462 = ( n_n3492 ) | ( n_n3491 ) | ( wire18057 ) | ( wire18058 ) ;
 assign wire18063 = ( wire135 ) | ( wire125 ) | ( wire725  &  n_n216 ) ;
 assign wire18064 = ( wire55 ) | ( wire127 ) | ( wire158 ) | ( wire133 ) ;
 assign n_n3489 = ( n_n3570 ) | ( n_n108  &  wire18063 ) | ( n_n108  &  wire18064 ) ;
 assign wire18078 = ( n_n3489 ) | ( wire3685 ) | ( wire18071 ) | ( wire18076 ) ;
 assign n_n3451 = ( n_n3460 ) | ( n_n3462 ) | ( wire18078 ) ;
 assign wire1754 = ( i_9_  &  (~ i_10_)  &  i_11_  &  wire721 ) | ( i_9_  &  i_10_  &  (~ i_11_)  &  wire721 ) ;
 assign wire1753 = ( (~ i_9_)  &  (~ i_10_)  &  i_11_  &  wire721 ) | ( (~ i_9_)  &  i_10_  &  (~ i_11_)  &  wire721 ) ;
 assign wire19630 = ( n_n170  &  wire720 ) | ( n_n170  &  wire715 ) | ( n_n170  &  wire724 ) ;
 assign wire1756 = ( wire237 ) | ( wire19630 ) ;
 assign wire19654 = ( n_n170  &  wire720 ) | ( n_n170  &  wire715 ) | ( n_n170  &  wire724 ) ;
 assign wire1758 = ( n_n84 ) | ( wire279 ) | ( wire237 ) | ( wire19654 ) ;
 assign wire19856 = ( n_n170  &  wire720 ) | ( n_n170  &  wire727 ) | ( n_n170  &  wire726 ) ;
 assign wire1761 = ( n_n171 ) | ( wire329 ) | ( wire336 ) | ( wire19856 ) ;
 assign wire18978 = ( i_9_  &  i_10_  &  i_11_  &  wire721 ) | ( i_9_  &  (~ i_10_)  &  i_11_  &  wire721 ) | ( (~ i_9_)  &  (~ i_10_)  &  (~ i_11_)  &  wire721 ) ;
 assign wire1766 = ( n_n137 ) | ( wire302 ) | ( wire316 ) | ( wire18978 ) ;
 assign wire19672 = ( wire720  &  n_n199 ) | ( wire715  &  n_n199 ) | ( n_n199  &  wire724 ) ;
 assign wire1775 = ( wire111 ) | ( wire291 ) | ( wire297 ) | ( wire19672 ) ;
 assign wire1779 = ( i_9_  &  i_10_  &  i_11_  &  wire728 ) | ( (~ i_9_)  &  (~ i_10_)  &  i_11_  &  wire728 ) | ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire728 ) ;
 assign wire1778 = ( i_9_  &  (~ i_10_)  &  i_11_  &  wire728 ) | ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire728 ) ;
 assign wire1777 = ( (~ i_9_)  &  i_10_  &  i_11_  &  wire728 ) | ( (~ i_9_)  &  (~ i_10_)  &  (~ i_11_)  &  wire728 ) ;
 assign wire1780 = ( i_15_  &  n_n205  &  n_n149 ) | ( (~ i_15_)  &  n_n205  &  n_n149 ) ;
 assign wire3403 = ( n_n112  &  wire222 ) | ( wire725  &  n_n191  &  n_n112 ) ;
 assign wire18342 = ( n_n113  &  n_n115 ) | ( n_n42  &  n_n183 ) ;
 assign wire18345 = ( wire3404 ) | ( n_n43  &  wire1786 ) ;
 assign wire1782 = ( wire51 ) | ( wire240 ) | ( wire187 ) | ( wire210 ) ;
 assign wire1786 = ( wire51 ) | ( wire240 ) | ( wire187 ) | ( wire210 ) ;
 assign wire19021 = ( n_n6445 ) | ( wire2712 ) | ( wire2730 ) | ( wire2731 ) ;
 assign wire19023 = ( wire19010 ) | ( wire19015 ) | ( _32040 ) ;
 assign n_n1801 = ( wire19021 ) | ( wire19023 ) | ( _2123 ) | ( _32003 ) ;
 assign wire4974 = ( wire132  &  n_n34 ) | ( n_n34  &  wire149 ) ;
 assign wire16952 = ( n_n34  &  wire147 ) | ( n_n34  &  wire181 ) ;
 assign wire16953 = ( wire137  &  n_n36 ) | ( n_n34  &  wire126 ) ;
 assign wire16954 = ( wire146  &  n_n36 ) | ( wire131  &  n_n36 ) | ( n_n36  &  wire46 ) ;
 assign n_n4419 = ( wire4974 ) | ( wire16952 ) | ( wire16953 ) | ( wire16954 ) ;
 assign wire202 = ( n_n184  &  wire730 ) | ( n_n184  &  wire717 ) | ( n_n184  &  wire724 ) ;
 assign wire307 = ( wire730  &  n_n191 ) | ( wire717  &  n_n191 ) | ( n_n191  &  wire724 ) ;
 assign wire17339 = ( n_n184  &  wire729 ) | ( n_n184  &  wire722 ) | ( n_n184  &  wire726 ) ;
 assign wire1794 = ( n_n189 ) | ( wire202 ) | ( wire307 ) | ( wire17339 ) ;
 assign wire17149 = ( n_n4441 ) | ( wire575 ) | ( wire17145 ) | ( wire17146 ) ;
 assign wire18004 = ( n_n184  &  wire719 ) | ( wire725  &  n_n199 ) ;
 assign wire1807 = ( wire171 ) | ( wire160 ) | ( wire242 ) | ( wire18004 ) ;
 assign wire19500 = ( wire720  &  n_n199 ) | ( wire715  &  n_n199 ) | ( n_n199  &  wire724 ) ;
 assign wire1809 = ( n_n103 ) | ( wire291 ) | ( wire297 ) | ( wire19500 ) ;
 assign wire18007 = ( n_n156  &  wire719 ) | ( wire725  &  n_n149 ) ;
 assign wire1811 = ( wire381 ) | ( wire186 ) | ( wire209 ) | ( wire18007 ) ;
 assign wire18014 = ( wire720  &  n_n149 ) | ( wire719  &  n_n216 ) ;
 assign wire1812 = ( wire60 ) | ( wire220 ) | ( wire218 ) | ( wire18014 ) ;
 assign wire17903 = ( n_n184  &  wire725 ) | ( n_n177  &  wire719 ) ;
 assign wire1814 = ( wire217 ) | ( wire209 ) | ( wire174 ) | ( wire17903 ) ;
 assign wire49 = ( wire721  &  n_n216 ) | ( wire728  &  n_n216 ) ;
 assign wire50 = ( n_n156  &  wire717 ) | ( n_n156  &  wire718 ) ;
 assign wire56 = ( wire717  &  n_n216 ) | ( n_n216  &  wire718 ) ;
 assign wire72 = ( n_n170  &  wire721 ) | ( n_n170  &  wire728 ) ;
 assign wire79 = ( n_n177  &  wire717 ) | ( n_n177  &  wire718 ) ;
 assign wire82 = ( n_n149  &  wire721 ) | ( n_n149  &  wire728 ) ;
 assign wire438 = ( i_15_  &  n_n149  &  n_n207 ) | ( (~ i_15_)  &  n_n149  &  n_n207 ) ;
 assign wire399 = ( wire717  &  n_n216 ) | ( wire724  &  n_n216 ) ;
 assign wire340 = ( i_15_  &  n_n184  &  n_n207 ) | ( (~ i_15_)  &  n_n184  &  n_n207 ) ;
 assign wire284 = ( wire720  &  n_n191 ) | ( wire727  &  n_n191 ) ;
 assign wire177 = ( i_15_  &  n_n184  &  n_n211 ) | ( (~ i_15_)  &  n_n184  &  n_n211 ) ;
 assign wire183 = ( i_15_  &  n_n170  &  n_n213 ) | ( (~ i_15_)  &  n_n170  &  n_n213 ) ;
 assign wire425 = ( i_15_  &  n_n199  &  n_n207 ) | ( (~ i_15_)  &  n_n199  &  n_n207 ) ;
 assign wire192 = ( i_15_  &  n_n199  &  n_n207 ) | ( (~ i_15_)  &  n_n199  &  n_n207 ) | ( (~ i_15_)  &  n_n199  &  n_n209 ) ;
 assign wire193 = ( i_15_  &  n_n211  &  n_n199 ) | ( (~ i_15_)  &  n_n211  &  n_n199 ) | ( i_15_  &  n_n199  &  n_n204 ) ;
 assign wire424 = ( i_15_  &  n_n156  &  n_n207 ) | ( (~ i_15_)  &  n_n156  &  n_n207 ) ;
 assign wire196 = ( i_15_  &  n_n211  &  n_n216 ) | ( (~ i_15_)  &  n_n211  &  n_n216 ) | ( i_15_  &  n_n216  &  n_n204 ) ;
 assign wire204 = ( wire719  &  n_n149 ) | ( n_n149  &  wire728 ) ;
 assign wire293 = ( wire729  &  n_n191 ) | ( wire717  &  n_n191 ) ;
 assign wire300 = ( i_15_  &  n_n149  &  n_n213 ) | ( (~ i_15_)  &  n_n149  &  n_n213 ) | ( (~ i_15_)  &  n_n149  &  n_n209 ) ;
 assign wire301 = ( i_15_  &  n_n211  &  n_n191 ) | ( (~ i_15_)  &  n_n211  &  n_n191 ) ;
 assign wire305 = ( n_n184  &  wire729 ) | ( n_n184  &  wire717 ) ;
 assign wire310 = ( n_n184  &  wire723 ) | ( n_n184  &  wire716 ) | ( n_n184  &  wire718 ) ;
 assign wire318 = ( wire723  &  n_n191 ) | ( n_n191  &  wire716 ) | ( n_n191  &  wire718 ) ;
 assign wire328 = ( i_15_  &  n_n199  &  n_n213 ) | ( (~ i_15_)  &  n_n199  &  n_n213 ) | ( (~ i_15_)  &  n_n199  &  n_n209 ) ;
 assign wire345 = ( wire729  &  n_n149 ) | ( wire717  &  n_n149 ) ;
 assign wire369 = ( i_15_  &  n_n211  &  n_n149 ) | ( (~ i_15_)  &  n_n211  &  n_n149 ) ;
 assign wire372 = ( wire729  &  n_n156 ) | ( n_n156  &  wire730 ) | ( n_n156  &  wire717 ) ;
 assign wire398 = ( n_n159  &  n_n218  &  n_n35 ) | ( n_n159  &  n_n218  &  n_n124 ) ;
 assign wire400 = ( wire729  &  n_n177 ) | ( n_n177  &  wire717 ) ;
 assign wire405 = ( i_9_  &  (~ i_10_)  &  i_11_  &  wire719 ) | ( (~ i_9_)  &  (~ i_10_)  &  (~ i_11_)  &  wire719 ) ;
 assign wire406 = ( i_9_  &  (~ i_10_)  &  i_11_  &  wire719 ) | ( (~ i_9_)  &  i_10_  &  (~ i_11_)  &  wire719 ) ;
 assign wire408 = ( wire728  &  n_n199 ) | ( n_n156  &  wire726 ) ;
 assign wire409 = ( i_9_  &  (~ i_10_)  &  i_11_  &  wire728 ) | ( (~ i_9_)  &  i_10_  &  (~ i_11_)  &  wire728 ) ;
 assign wire410 = ( i_9_  &  i_10_  &  i_11_  &  wire721 ) | ( (~ i_9_)  &  (~ i_10_)  &  (~ i_11_)  &  wire721 ) ;
 assign wire414 = ( i_9_  &  i_10_  &  i_11_  &  wire728 ) | ( (~ i_9_)  &  (~ i_10_)  &  (~ i_11_)  &  wire728 ) ;
 assign wire416 = ( (~ i_9_)  &  i_10_  &  i_11_  &  wire728 ) | ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire728 ) ;
 assign wire418 = ( i_9_  &  i_10_  &  i_11_  &  wire725 ) | ( (~ i_9_)  &  (~ i_10_)  &  (~ i_11_)  &  wire725 ) ;
 assign wire1840 = ( wire219 ) | ( wire108 ) | ( n_n198 ) | ( wire258 ) ;
 assign wire16980 = ( wire729  &  n_n199 ) | ( wire720  &  n_n199 ) | ( n_n199  &  wire726 ) ;
 assign wire1853 = ( wire219 ) | ( wire108 ) | ( n_n198 ) | ( wire258 ) ;
 assign wire1862 = ( wire725  &  n_n199 ) | ( wire719  &  n_n216 ) ;
 assign wire815 = ( n_n159  &  n_n35  &  n_n111 ) | ( n_n159  &  n_n124  &  n_n111 ) ;
 assign wire1128 = ( n_n156  &  wire723 ) | ( wire723  &  n_n149 ) | ( n_n149  &  wire718 ) ;
 assign wire1209 = ( n_n177  &  wire721 ) | ( n_n170  &  wire721 ) | ( n_n170  &  wire728 ) ;
 assign wire1253 = ( n_n177  &  wire721 ) | ( n_n170  &  wire721 ) | ( n_n170  &  wire728 ) ;
 assign wire1409 = ( wire721  &  n_n199 ) | ( wire728  &  n_n199 ) | ( wire721  &  n_n216 ) | ( wire728  &  n_n216 ) ;
 assign wire1550 = ( n_n159  &  n_n35  &  n_n111 ) | ( n_n159  &  n_n124  &  n_n111 ) ;
 assign wire1557 = ( n_n170  &  wire721 ) | ( n_n177  &  wire728 ) | ( n_n170  &  wire728 ) ;
 assign wire138 = ( wire270  &  n_n2 ) | ( n_n2  &  wire372 ) ;
 assign wire439 = ( (~ i_7_)  &  i_6_  &  n_n48  &  n_n19 ) | ( i_7_  &  (~ i_6_)  &  n_n48  &  n_n19 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n48  &  n_n19 ) ;
 assign wire467 = ( n_n5  &  wire145 ) | ( n_n5  &  n_n151 ) | ( n_n5  &  wire370 ) ;
 assign wire499 = ( n_n30  &  wire110 ) | ( n_n30  &  wire249 ) | ( n_n30  &  wire19905 ) ;
 assign wire19899 = ( wire720  &  n_n191 ) | ( wire727  &  n_n191 ) | ( n_n191  &  wire726 ) ;
 assign wire507 = ( n_n31  &  wire337 ) | ( n_n31  &  wire338 ) | ( n_n31  &  wire19899 ) ;
 assign wire510 = ( n_n30  &  wire337 ) | ( n_n30  &  wire284 ) ;
 assign wire513 = ( n_n31  &  wire314 ) | ( n_n184  &  n_n31  &  wire726 ) ;
 assign wire520 = ( n_n31  &  wire329 ) | ( n_n31  &  wire161 ) ;
 assign wire552 = ( n_n30  &  wire248 ) | ( n_n30  &  n_n64 ) | ( n_n30  &  wire408 ) ;
 assign wire19888 = ( n_n149  &  wire726 ) | ( wire728  &  n_n216 ) ;
 assign wire556 = ( n_n36  &  wire19888 ) | ( n_n149  &  n_n36  &  wire718 ) ;
 assign wire1906 = ( n_n218  &  n_n35  &  n_n220  &  wire1779 ) ;
 assign wire1907 = ( n_n30  &  wire335 ) | ( n_n30  &  wire295 ) | ( n_n30  &  wire19882 ) ;
 assign wire19879 = ( (~ i_9_)  &  (~ i_10_)  &  i_11_  &  wire728 ) | ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire728 ) ;
 assign wire1910 = ( n_n33  &  wire278 ) | ( n_n33  &  wire19879 ) ;
 assign wire1912 = ( n_n184  &  wire728  &  n_n32 ) ;
 assign wire1914 = ( n_n32  &  wire269 ) | ( n_n32  &  wire275 ) ;
 assign wire1940 = ( n_n123  &  wire329 ) | ( n_n123  &  wire259 ) | ( n_n123  &  wire19856 ) ;
 assign wire19848 = ( n_n156  &  wire726 ) | ( wire728  &  n_n216 ) ;
 assign wire1945 = ( n_n125  &  wire207 ) | ( n_n125  &  wire416 ) | ( n_n125  &  wire19848 ) ;
 assign wire19850 = ( wire728  &  n_n191 ) | ( n_n149  &  wire726 ) ;
 assign wire1951 = ( n_n108  &  wire335 ) | ( n_n108  &  wire333 ) ;
 assign wire1960 = ( n_n123  &  wire336 ) | ( n_n177  &  wire726  &  n_n123 ) ;
 assign wire1961 = ( n_n125  &  wire248 ) | ( n_n125  &  wire110 ) ;
 assign wire1962 = ( n_n125  &  n_n202 ) | ( n_n125  &  wire295 ) | ( n_n125  &  wire19835 ) ;
 assign wire1968 = ( n_n218  &  n_n220  &  n_n126  &  wire1513 ) ;
 assign wire1971 = ( n_n125  &  wire314 ) | ( n_n125  &  wire338 ) ;
 assign wire1972 = ( n_n125  &  wire335 ) | ( n_n125  &  wire333 ) ;
 assign wire19827 = ( i_9_  &  i_10_  &  i_11_  &  wire728 ) | ( i_9_  &  (~ i_10_)  &  i_11_  &  wire728 ) | ( (~ i_9_)  &  (~ i_10_)  &  (~ i_11_)  &  wire728 ) ;
 assign wire1976 = ( n_n197  &  n_n60 ) | ( n_n197  &  wire235 ) | ( n_n197  &  wire19827 ) ;
 assign wire1979 = ( wire244  &  n_n197 ) | ( wire140  &  n_n197 ) ;
 assign wire19770 = ( i_9_  &  (~ i_10_)  &  i_11_  &  wire726 ) | ( (~ i_9_)  &  (~ i_10_)  &  i_11_  &  wire726 ) ;
 assign wire1982 = ( n_n101  &  wire336 ) | ( n_n101  &  wire259 ) | ( n_n101  &  wire19770 ) ;
 assign wire1983 = ( _314 ) | ( n_n108  &  wire248 ) | ( n_n108  &  wire161 ) ;
 assign wire1987 = ( n_n108  &  n_n202 ) | ( n_n108  &  wire295 ) | ( n_n108  &  wire19767 ) ;
 assign wire1990 = ( n_n101  &  wire338 ) | ( n_n101  &  wire726  &  n_n216 ) ;
 assign wire19766 = ( wire720  &  n_n191 ) | ( wire727  &  n_n191 ) | ( n_n191  &  wire726 ) ;
 assign wire1991 = ( n_n108  &  wire337 ) | ( n_n108  &  wire19766 ) ;
 assign wire19760 = ( i_9_  &  (~ i_10_)  &  i_11_  &  wire726 ) | ( (~ i_9_)  &  (~ i_10_)  &  (~ i_11_)  &  wire726 ) ;
 assign wire1992 = ( n_n108  &  wire336 ) | ( n_n108  &  wire259 ) | ( n_n108  &  wire19760 ) ;
 assign wire1995 = ( n_n101  &  wire314 ) | ( n_n184  &  n_n101  &  wire726 ) ;
 assign wire1996 = ( n_n108  &  wire314 ) | ( n_n108  &  wire338 ) ;
 assign wire1997 = ( n_n108  &  wire207 ) | ( n_n156  &  wire726  &  n_n108 ) ;
 assign wire19759 = ( wire720  &  n_n149 ) | ( wire727  &  n_n149 ) | ( n_n149  &  wire726 ) ;
 assign wire1998 = ( n_n101  &  wire249 ) | ( n_n101  &  wire19759 ) ;
 assign wire1999 = ( n_n48  &  n_n220  &  n_n161  &  wire1641 ) ;
 assign wire2000 = ( _453 ) | ( wire244  &  n_n47 ) | ( wire140  &  n_n47 ) ;
 assign wire2004 = ( n_n43  &  wire63 ) | ( n_n43  &  wire348 ) ;
 assign wire19780 = ( (~ i_15_)  &  n_n156  &  n_n209 ) | ( i_15_  &  n_n156  &  n_n215 ) | ( (~ i_15_)  &  n_n156  &  n_n215 ) ;
 assign wire2026 = ( n_n101  &  wire248 ) | ( n_n101  &  wire409 ) | ( n_n101  &  wire19780 ) ;
 assign wire19782 = ( i_9_  &  i_10_  &  (~ i_11_)  &  wire728 ) | ( (~ i_9_)  &  i_10_  &  (~ i_11_)  &  wire728 ) ;
 assign wire19783 = ( n_n177  &  wire728 ) | ( n_n149  &  wire726 ) ;
 assign wire2027 = ( n_n108  &  wire249 ) | ( n_n108  &  wire19782 ) | ( n_n108  &  wire19783 ) ;
 assign wire19778 = ( i_9_  &  i_10_  &  i_11_  &  wire728 ) | ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire728 ) ;
 assign wire2032 = ( n_n101  &  wire408 ) | ( n_n101  &  wire19778 ) ;
 assign wire2041 = ( n_n43  &  wire346 ) | ( wire728  &  n_n191  &  n_n43 ) ;
 assign wire2045 = ( n_n41  &  wire169 ) | ( n_n41  &  wire415 ) ;
 assign wire19727 = ( n_n156  &  wire720 ) | ( n_n170  &  wire718 ) ;
 assign wire19728 = ( i_15_  &  n_n156  &  n_n205 ) | ( (~ i_15_)  &  n_n156  &  n_n205 ) | ( (~ i_15_)  &  n_n205  &  n_n170 ) ;
 assign wire2062 = ( n_n36  &  wire156 ) | ( n_n36  &  wire19727 ) | ( n_n36  &  wire19728 ) ;
 assign wire19724 = ( n_n170  &  wire720 ) | ( n_n177  &  wire718 ) ;
 assign wire2068 = ( n_n36  &  wire19724 ) | ( n_n177  &  n_n36  &  wire726 ) ;
 assign wire2070 = ( n_n34  &  wire128 ) | ( n_n34  &  wire348 ) ;
 assign wire2078 = ( n_n34  &  wire346 ) | ( wire720  &  n_n34  &  n_n191 ) ;
 assign wire19716 = ( i_15_  &  n_n184  &  n_n205 ) | ( (~ i_15_)  &  n_n184  &  n_n205 ) | ( i_15_  &  n_n184  &  n_n215 ) ;
 assign wire2079 = ( n_n36  &  wire128 ) | ( n_n36  &  wire19716 ) ;
 assign wire19714 = ( i_15_  &  n_n205  &  n_n216 ) | ( (~ i_15_)  &  n_n205  &  n_n216 ) | ( i_15_  &  n_n216  &  n_n215 ) ;
 assign wire2099 = ( wire270  &  n_n3 ) | ( n_n3  &  wire372 ) ;
 assign wire2108 = ( n_n162  &  n_n35  &  n_n220  &  wire1415 ) ;
 assign wire2119 = ( n_n125  &  n_n103 ) | ( n_n125  &  wire297 ) | ( n_n125  &  wire19672 ) ;
 assign wire2124 = ( n_n212  &  n_n138 ) | ( n_n212  &  wire163 ) | ( n_n212  &  wire405 ) ;
 assign wire2125 = ( n_n197  &  n_n138 ) | ( n_n197  &  wire407 ) | ( n_n197  &  wire163 ) ;
 assign wire2130 = ( n_n197  &  wire134 ) | ( n_n197  &  wire194 ) ;
 assign wire2134 = ( n_n218  &  n_n124  &  n_n220  &  wire1261 ) ;
 assign wire2136 = ( n_n123  &  wire54 ) | ( wire724  &  n_n216  &  n_n123 ) ;
 assign wire2139 = ( n_n125  &  wire111 ) | ( n_n125  &  wire291 ) ;
 assign wire2141 = ( n_n123  &  wire104 ) | ( n_n123  &  wire237 ) | ( n_n123  &  wire19654 ) ;
 assign wire2146 = ( n_n112  &  wire187 ) | ( wire720  &  n_n191  &  n_n112 ) ;
 assign wire2149 = ( n_n218  &  n_n220  &  n_n126  &  wire1089 ) ;
 assign wire2153 = ( n_n108  &  wire111 ) | ( n_n108  &  wire291 ) ;
 assign wire2155 = ( n_n123  &  wire279 ) | ( n_n177  &  wire724  &  n_n123 ) ;
 assign wire2156 = ( n_n125  &  wire290 ) | ( n_n125  &  wire59 ) ;
 assign wire2157 = ( wire118  &  n_n125 ) | ( n_n125  &  n_n72 ) | ( n_n125  &  wire401 ) ;
 assign wire2163 = ( n_n125  &  wire199 ) | ( n_n149  &  wire724  &  n_n125 ) ;
 assign wire2169 = ( n_n101  &  wire104 ) | ( n_n170  &  n_n101  &  wire724 ) ;
 assign wire2174 = ( n_n108  &  wire104 ) | ( n_n184  &  wire724  &  n_n108 ) ;
 assign wire2176 = ( n_n108  &  n_n103 ) | ( n_n108  &  wire297 ) | ( n_n108  &  wire19621 ) ;
 assign wire2179 = ( n_n101  &  wire54 ) | ( n_n101  &  wire724  &  n_n216 ) ;
 assign wire19620 = ( wire720  &  n_n191 ) | ( wire715  &  n_n191 ) | ( n_n191  &  wire724 ) ;
 assign wire2180 = ( n_n108  &  wire320 ) | ( n_n108  &  wire19620 ) ;
 assign wire2181 = ( wire47  &  n_n47 ) | ( n_n47  &  wire322 ) | ( n_n47  &  wire192 ) ;
 assign wire19605 = ( n_n156  &  wire719 ) | ( n_n156  &  wire720 ) | ( n_n156  &  wire715 ) ;
 assign wire2190 = ( n_n101  &  wire290 ) | ( n_n101  &  wire406 ) | ( n_n101  &  wire19605 ) ;
 assign wire19607 = ( n_n156  &  wire719 ) | ( n_n149  &  wire724 ) ;
 assign wire19608 = ( i_9_  &  (~ i_10_)  &  i_11_  &  wire719 ) | ( (~ i_9_)  &  i_10_  &  (~ i_11_)  &  wire719 ) ;
 assign wire2191 = ( n_n108  &  wire199 ) | ( n_n108  &  wire19607 ) | ( n_n108  &  wire19608 ) ;
 assign wire19602 = ( i_9_  &  i_10_  &  i_11_  &  wire719 ) | ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire719 ) ;
 assign wire2195 = ( n_n101  &  wire402 ) | ( n_n101  &  wire19602 ) ;
 assign wire2197 = ( n_n184  &  wire719  &  wire228 ) ;
 assign wire2205 = ( wire132  &  n_n46 ) | ( n_n46  &  wire280 ) | ( n_n46  &  wire121 ) ;
 assign wire19535 = ( i_15_  &  n_n216  &  n_n207 ) | ( (~ i_15_)  &  n_n216  &  n_n207 ) | ( i_15_  &  n_n216  &  n_n215 ) ;
 assign wire2269 = ( n_n36  &  wire85 ) | ( n_n36  &  wire19535 ) ;
 assign wire19530 = ( i_15_  &  n_n170  &  n_n207 ) | ( (~ i_15_)  &  n_n170  &  n_n207 ) | ( i_15_  &  n_n170  &  n_n215 ) ;
 assign wire2277 = ( n_n34  &  wire208 ) | ( n_n34  &  wire100 ) | ( n_n34  &  wire19530 ) ;
 assign wire19531 = ( i_15_  &  n_n177  &  n_n207 ) | ( (~ i_15_)  &  n_n177  &  n_n207 ) ;
 assign wire2278 = ( n_n36  &  wire208 ) | ( n_n36  &  wire19530 ) | ( n_n36  &  wire19531 ) ;
 assign wire19528 = ( wire720  &  n_n149 ) | ( n_n177  &  wire716 ) ;
 assign wire19529 = ( i_15_  &  n_n156  &  n_n207 ) | ( (~ i_15_)  &  n_n156  &  n_n207 ) | ( i_15_  &  n_n156  &  n_n215 ) ;
 assign wire2282 = ( n_n36  &  wire215 ) | ( n_n36  &  wire19529 ) ;
 assign wire2283 = ( n_n34  &  n_n190 ) | ( n_n34  &  wire107 ) | ( n_n34  &  wire340 ) ;
 assign wire2287 = ( n_n34  &  wire187 ) | ( n_n34  &  wire339 ) ;
 assign wire2290 = ( n_n34  &  wire219 ) | ( n_n34  &  wire425 ) ;
 assign wire2293 = ( n_n36  &  wire425 ) | ( wire720  &  n_n36  &  n_n191 ) ;
 assign wire19519 = ( i_15_  &  n_n216  &  n_n207 ) | ( (~ i_15_)  &  n_n216  &  n_n207 ) | ( i_15_  &  n_n216  &  n_n215 ) ;
 assign wire2294 = ( n_n34  &  wire85 ) | ( n_n34  &  wire19519 ) ;
 assign wire2295 = ( wire47  &  n_n212 ) | ( n_n212  &  wire322 ) | ( n_n212  &  wire192 ) ;
 assign wire2296 = ( n_n197  &  wire151 ) | ( n_n197  &  wire322 ) | ( n_n197  &  wire192 ) ;
 assign wire19486 = ( wire720  &  n_n149 ) | ( wire719  &  n_n216 ) ;
 assign wire2323 = ( n_n36  &  wire84 ) | ( n_n36  &  wire438 ) | ( n_n36  &  wire19486 ) ;
 assign wire2324 = ( _1126 ) | ( n_n34  &  wire84 ) | ( n_n34  &  wire424 ) ;
 assign wire19472 = ( (~ i_9_)  &  (~ i_10_)  &  i_11_  &  wire724 ) | ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire724 ) ;
 assign wire2335 = ( n_n30  &  wire53 ) | ( n_n30  &  wire237 ) | ( n_n30  &  wire19472 ) ;
 assign wire2340 = ( n_n31  &  n_n90 ) | ( n_n31  &  wire195 ) | ( n_n31  &  wire19469 ) ;
 assign wire2343 = ( n_n30  &  wire291 ) | ( n_n30  &  wire724  &  n_n216 ) ;
 assign wire2344 = ( n_n31  &  wire98 ) | ( n_n31  &  wire320 ) ;
 assign wire2345 = ( n_n30  &  wire199 ) | ( n_n30  &  wire59 ) | ( n_n30  &  wire19464 ) ;
 assign wire2349 = ( n_n30  &  n_n142 ) | ( n_n30  &  wire290 ) | ( n_n30  &  wire402 ) ;
 assign wire2350 = ( n_n31  &  wire59 ) | ( n_n31  &  n_n170  &  wire724 ) ;
 assign wire19461 = ( n_n177  &  wire720 ) | ( n_n177  &  wire715 ) | ( n_n177  &  wire724 ) ;
 assign wire2351 = ( n_n30  &  wire279 ) | ( n_n30  &  wire19461 ) ;
 assign wire19447 = ( n_n177  &  wire721 ) | ( n_n177  &  wire728 ) ;
 assign wire19448 = ( n_n156  &  wire721 ) | ( n_n149  &  wire721 ) | ( n_n156  &  wire728 ) | ( n_n149  &  wire728 ) ;
 assign wire2352 = ( n_n30  &  wire19447 ) | ( n_n30  &  wire19448 ) ;
 assign wire19449 = ( n_n149  &  wire721 ) | ( n_n149  &  wire728 ) ;
 assign wire19450 = ( n_n156  &  wire721 ) | ( n_n170  &  wire721 ) | ( n_n156  &  wire728 ) | ( n_n170  &  wire728 ) ;
 assign wire2353 = ( n_n31  &  wire19449 ) | ( n_n31  &  wire19450 ) ;
 assign wire19440 = ( wire721  &  n_n199 ) | ( wire728  &  n_n199 ) ;
 assign wire19441 = ( wire721  &  n_n191 ) | ( wire728  &  n_n191 ) | ( wire721  &  n_n216 ) | ( wire728  &  n_n216 ) ;
 assign wire19438 = ( n_n184  &  wire721 ) | ( wire721  &  n_n191 ) | ( wire728  &  n_n191 ) ;
 assign wire2359 = ( n_n30  &  wire72 ) | ( n_n30  &  wire19438 ) ;
 assign wire19426 = ( n_n170  &  wire727 ) | ( n_n170  &  wire716 ) ;
 assign wire2364 = ( n_n38  &  wire53 ) | ( n_n38  &  wire19426 ) ;
 assign wire19427 = ( n_n170  &  wire720 ) | ( n_n177  &  wire716 ) ;
 assign wire2365 = ( n_n39  &  wire384 ) | ( n_n39  &  wire19427 ) ;
 assign wire2370 = ( n_n40  &  wire65 ) | ( n_n40  &  wire1557 ) ;
 assign wire19424 = ( n_n156  &  wire721 ) | ( n_n177  &  wire721 ) | ( n_n156  &  wire728 ) ;
 assign wire2372 = ( n_n40  &  wire82 ) | ( n_n40  &  wire19424 ) ;
 assign wire2374 = ( n_n40  &  wire127 ) | ( n_n40  &  wire133 ) ;
 assign wire19411 = ( n_n184  &  wire721 ) | ( n_n184  &  wire728 ) | ( wire721  &  n_n191 ) | ( wire728  &  n_n191 ) ;
 assign wire19412 = ( wire721  &  n_n199 ) | ( wire728  &  n_n199 ) | ( wire721  &  n_n216 ) | ( wire728  &  n_n216 ) ;
 assign wire2382 = ( n_n40  &  wire155 ) | ( n_n40  &  wire227 ) ;
 assign wire2384 = ( n_n34  &  wire223 ) | ( n_n34  &  wire274 ) ;
 assign wire2393 = ( n_n34  &  wire184 ) | ( n_n34  &  wire246 ) | ( n_n34  &  wire254 ) ;
 assign wire2398 = ( n_n36  &  wire179 ) | ( n_n36  &  wire223 ) | ( n_n36  &  wire239 ) ;
 assign wire2404 = ( n_n34  &  wire179 ) | ( n_n34  &  wire239 ) ;
 assign wire19387 = ( wire63 ) | ( wire52 ) | ( wire51 ) | ( wire148 ) ;
 assign wire2407 = ( n_n30  &  wire277 ) | ( n_n30  &  wire274 ) | ( n_n30  &  wire19387 ) ;
 assign wire2410 = ( n_n31  &  wire155 ) | ( n_n31  &  wire227 ) | ( n_n31  &  wire69 ) ;
 assign wire2415 = ( _1401 ) | ( n_n31  &  wire276 ) | ( n_n31  &  wire211 ) ;
 assign wire2417 = ( n_n34  &  wire70 ) | ( n_n34  &  wire233 ) ;
 assign wire2418 = ( n_n36  &  wire206 ) | ( n_n36  &  wire330 ) | ( n_n36  &  wire328 ) ;
 assign wire2424 = ( n_n34  &  wire142 ) | ( n_n34  &  wire251 ) ;
 assign wire2427 = ( n_n38  &  n_n173 ) | ( n_n38  &  wire249 ) | ( n_n38  &  wire384 ) ;
 assign wire2428 = ( n_n48  &  n_n220  &  n_n126  &  wire1003 ) ;
 assign wire2435 = ( n_n36  &  wire142 ) | ( n_n36  &  wire233 ) | ( n_n36  &  wire251 ) ;
 assign wire19339 = ( wire729  &  n_n170 ) | ( n_n170  &  wire717 ) | ( n_n170  &  wire726 ) ;
 assign wire2442 = ( n_n46  &  wire281 ) | ( n_n46  &  wire57 ) | ( n_n46  &  wire19339 ) ;
 assign wire2448 = ( n_n46  &  wire139 ) | ( n_n46  &  wire128 ) | ( n_n46  &  wire62 ) ;
 assign wire19337 = ( n_n183 ) | ( wire184 ) | ( wire246 ) | ( wire210 ) ;
 assign wire2449 = ( n_n47  &  wire349 ) | ( n_n47  &  wire357 ) | ( n_n47  &  wire19337 ) ;
 assign wire2451 = ( wire137  &  n_n47 ) | ( wire146  &  n_n47 ) | ( n_n47  &  wire254 ) ;
 assign wire2452 = ( n_n48  &  n_n220  &  n_n161  &  wire1507 ) ;
 assign wire2462 = ( wire720  &  n_n199  &  _32250 ) | ( wire715  &  n_n199  &  _32250 ) ;
 assign wire2463 = ( n_n101  &  wire123 ) | ( n_n101  &  wire88 ) | ( n_n101  &  wire1409 ) ;
 assign wire19315 = ( n_n184  &  wire728 ) | ( wire721  &  n_n191 ) | ( wire728  &  n_n191 ) ;
 assign wire2464 = ( n_n108  &  wire1409 ) | ( n_n108  &  wire19315 ) ;
 assign wire19312 = ( n_n184  &  wire721 ) | ( n_n177  &  wire721 ) | ( n_n177  &  wire728 ) ;
 assign wire2468 = ( n_n108  &  wire72 ) | ( n_n108  &  wire19312 ) ;
 assign wire2475 = ( n_n48  &  wire714  &  n_n18  &  wire1341 ) ;
 assign wire2480 = ( wire126  &  n_n101 ) | ( wire147  &  n_n101 ) | ( n_n101  &  wire53 ) ;
 assign wire19297 = ( wire729  &  n_n177 ) | ( n_n177  &  wire726 ) ;
 assign wire2481 = ( n_n108  &  wire79 ) | ( n_n108  &  wire19297 ) ;
 assign wire19295 = ( wire729  &  n_n191 ) | ( wire717  &  n_n191 ) | ( n_n191  &  wire726 ) ;
 assign wire2487 = ( n_n101  &  wire241 ) | ( n_n101  &  wire19295 ) ;
 assign wire2489 = ( _1862 ) | ( n_n101  &  wire221 ) | ( n_n101  &  wire315 ) ;
 assign wire19290 = ( wire729  &  n_n149 ) | ( wire727  &  n_n149 ) ;
 assign wire19291 = ( wire720  &  n_n149 ) | ( wire715  &  n_n149 ) | ( n_n149  &  wire726 ) ;
 assign wire2490 = ( n_n108  &  wire75 ) | ( n_n108  &  wire19290 ) | ( n_n108  &  wire19291 ) ;
 assign wire19279 = ( wire729  &  n_n177 ) | ( n_n177  &  wire726 ) ;
 assign wire2493 = ( n_n101  &  wire384 ) | ( n_n101  &  wire79 ) | ( n_n101  &  wire19279 ) ;
 assign wire2498 = ( n_n125  &  wire251 ) | ( n_n125  &  wire328 ) ;
 assign wire19246 = ( n_n156  &  wire721 ) | ( n_n156  &  wire728 ) | ( n_n149  &  wire728 ) ;
 assign wire2518 = ( n_n212  &  wire72 ) | ( n_n212  &  wire19246 ) ;
 assign wire19245 = ( n_n184  &  wire728 ) | ( wire721  &  n_n216 ) | ( wire728  &  n_n216 ) ;
 assign wire2523 = ( n_n197  &  wire92 ) | ( n_n197  &  wire19245 ) ;
 assign wire19243 = ( n_n184  &  wire721 ) | ( wire721  &  n_n191 ) | ( wire728  &  n_n191 ) ;
 assign wire2525 = ( n_n197  &  wire72 ) | ( n_n197  &  wire19243 ) ;
 assign wire2526 = ( n_n123  &  n_n183 ) | ( n_n123  &  wire233 ) | ( n_n123  &  wire251 ) ;
 assign wire2532 = ( n_n197  &  wire74 ) | ( n_n197  &  wire68 ) | ( n_n197  &  wire81 ) ;
 assign wire2537 = ( n_n212  &  n_n198 ) | ( n_n212  &  wire206 ) | ( n_n212  &  wire328 ) ;
 assign wire2545 = ( n_n125  &  wire142 ) | ( n_n125  &  wire233 ) ;
 assign wire2548 = ( n_n71  &  n_n123 ) | ( n_n123  &  wire92 ) | ( n_n123  &  wire49 ) ;
 assign wire19204 = ( n_n177  &  wire728 ) | ( wire721  &  n_n191 ) | ( wire728  &  n_n191 ) ;
 assign wire2557 = ( n_n125  &  wire88 ) | ( n_n125  &  wire19204 ) ;
 assign wire2559 = ( n_n125  &  wire83 ) | ( n_n125  &  wire1253 ) ;
 assign wire2560 = ( wire143  &  n_n101 ) | ( wire154  &  n_n101 ) | ( n_n101  &  wire111 ) ;
 assign wire19194 = ( i_15_  &  n_n191  &  n_n213 ) | ( (~ i_15_)  &  n_n191  &  n_n213 ) | ( (~ i_15_)  &  n_n191  &  n_n209 ) ;
 assign wire2565 = ( n_n108  &  wire241 ) | ( n_n108  &  wire19194 ) ;
 assign wire2567 = ( n_n220  &  n_n111  &  wire16987  &  wire1072 ) ;
 assign wire2568 = ( n_n101  &  wire206 ) | ( n_n101  &  wire330 ) | ( n_n101  &  wire328 ) ;
 assign wire2578 = ( n_n123  &  wire148 ) | ( n_n123  &  wire277 ) | ( n_n123  &  wire274 ) ;
 assign wire2579 = ( _1679 ) | ( wire179  &  n_n125 ) | ( n_n125  &  wire223 ) ;
 assign wire2584 = ( n_n125  &  wire276 ) | ( n_n125  &  wire211 ) | ( n_n125  &  wire271 ) ;
 assign wire2588 = ( n_n125  &  wire227 ) | ( n_n125  &  wire232 ) ;
 assign wire2594 = ( n_n125  &  wire221 ) | ( n_n125  &  wire315 ) | ( n_n125  &  wire300 ) ;
 assign wire2598 = ( wire98  &  n_n112 ) | ( wire52  &  n_n112 ) | ( n_n112  &  wire51 ) ;
 assign wire19150 = ( n_n184  &  wire729 ) | ( n_n184  &  wire728 ) ;
 assign wire2599 = ( n_n113  &  wire211 ) | ( n_n113  &  wire271 ) | ( n_n113  &  wire19150 ) ;
 assign wire2614 = ( n_n30  &  wire74 ) | ( n_n30  &  wire68 ) ;
 assign wire2615 = ( n_n31  &  wire142 ) | ( n_n31  &  wire233 ) | ( n_n31  &  wire251 ) ;
 assign wire19128 = ( n_n201  &  _32665 ) | ( n_n201  &  _32666 ) ;
 assign wire19129 = ( n_n170  &  wire721 ) | ( n_n170  &  wire728 ) | ( wire728  &  n_n191 ) ;
 assign wire2618 = ( n_n33  &  wire19128 ) | ( n_n33  &  wire19129 ) ;
 assign wire2630 = ( n_n48  &  wire714  &  n_n18  &  wire1582 ) ;
 assign wire19113 = ( n_n156  &  wire727 ) | ( wire728  &  n_n191 ) ;
 assign wire2634 = ( n_n48  &  wire714  &  n_n18  &  wire1553 ) ;
 assign wire19110 = ( n_n156  &  wire717 ) | ( wire721  &  n_n199 ) ;
 assign wire2635 = ( n_n46  &  wire90 ) | ( n_n46  &  n_n62 ) | ( n_n46  &  wire19110 ) ;
 assign wire2636 = ( n_n43  &  wire210 ) | ( n_n43  &  wire357 ) ;
 assign wire2645 = ( n_n41  &  wire206 ) | ( n_n41  &  wire330 ) | ( n_n41  &  wire328 ) ;
 assign wire2646 = ( _1289 ) | ( n_n40  &  wire74 ) | ( n_n40  &  wire68 ) ;
 assign wire2657 = ( n_n17  &  n_n48  &  wire714  &  wire1295 ) ;
 assign wire2666 = ( n_n42  &  wire349 ) | ( n_n42  &  wire210 ) ;
 assign wire2669 = ( n_n41  &  wire126 ) | ( n_n41  &  wire147 ) ;
 assign wire2676 = ( n_n17  &  n_n48  &  wire714  &  wire1154 ) ;
 assign wire2679 = ( n_n40  &  wire63 ) | ( n_n40  &  wire52 ) | ( n_n40  &  wire277 ) ;
 assign wire2691 = ( n_n36  &  wire83 ) | ( n_n36  &  wire1209 ) ;
 assign wire2692 = ( n_n34  &  wire118 ) | ( n_n34  &  wire60 ) ;
 assign wire19043 = ( n_n71 ) | ( wire155 ) | ( wire92 ) | ( wire49 ) ;
 assign wire2700 = ( n_n34  &  wire227 ) | ( n_n34  &  wire232 ) | ( n_n34  &  wire19043 ) ;
 assign wire19038 = ( n_n177  &  wire728 ) | ( wire721  &  n_n191 ) | ( wire728  &  n_n191 ) ;
 assign wire2703 = ( n_n36  &  wire88 ) | ( n_n36  &  wire19038 ) ;
 assign wire2704 = ( n_n30  &  wire197 ) | ( n_n30  &  wire203 ) | ( n_n30  &  wire323 ) ;
 assign wire2705 = ( n_n31  &  wire203 ) | ( n_n31  &  wire309 ) | ( n_n31  &  wire323 ) ;
 assign wire19016 = ( (~ i_9_)  &  (~ i_10_)  &  i_11_  &  wire715 ) | ( i_9_  &  i_10_  &  (~ i_11_)  &  wire715 ) ;
 assign wire2712 = ( n_n41  &  wire230 ) | ( n_n41  &  wire352 ) | ( n_n41  &  wire19016 ) ;
 assign wire2717 = ( n_n40  &  n_n107 ) | ( n_n40  &  wire264 ) | ( n_n40  &  wire19013 ) ;
 assign wire2720 = ( n_n184  &  wire721  &  wire1277 ) | ( wire721  &  n_n191  &  wire1277 ) ;
 assign wire2721 = ( n_n162  &  n_n220  &  n_n161  &  wire52 ) ;
 assign wire2724 = ( wire1704  &  wire318 ) | ( wire715  &  n_n191  &  wire1704 ) ;
 assign wire2726 = ( n_n41  &  wire305 ) | ( n_n41  &  wire310 ) ;
 assign wire2728 = ( n_n41  &  wire293 ) | ( n_n184  &  wire715  &  n_n41 ) ;
 assign wire19008 = ( n_n184  &  wire729 ) | ( n_n184  &  wire715 ) | ( n_n184  &  wire717 ) ;
 assign wire2729 = ( n_n40  &  wire310 ) | ( n_n40  &  wire19008 ) ;
 assign wire2730 = ( n_n40  &  wire293 ) | ( n_n170  &  wire715  &  n_n40 ) ;
 assign wire19006 = ( n_n177  &  wire715 ) | ( n_n177  &  wire717 ) ;
 assign wire2731 = ( n_n41  &  wire380 ) | ( n_n41  &  wire19006 ) ;
 assign wire2733 = ( n_n101  &  n_n107 ) | ( n_n101  &  wire264 ) | ( n_n101  &  wire19001 ) ;
 assign wire2738 = ( n_n101  &  wire261 ) | ( n_n101  &  wire375 ) ;
 assign wire2739 = ( n_n108  &  wire318 ) | ( wire715  &  n_n191  &  n_n108 ) ;
 assign wire18993 = ( (~ i_9_)  &  (~ i_10_)  &  i_11_  &  wire715 ) | ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire715 ) ;
 assign wire2740 = ( n_n101  &  wire293 ) | ( n_n101  &  wire318 ) | ( n_n101  &  wire18993 ) ;
 assign wire2743 = ( n_n108  &  wire293 ) | ( n_n184  &  wire715  &  n_n108 ) ;
 assign wire18992 = ( n_n184  &  wire729 ) | ( n_n184  &  wire715 ) | ( n_n184  &  wire717 ) ;
 assign wire2744 = ( n_n101  &  wire310 ) | ( n_n101  &  wire18992 ) ;
 assign wire2748 = ( n_n108  &  wire352 ) | ( n_n156  &  wire715  &  n_n108 ) ;
 assign wire18956 = ( wire715  &  n_n149 ) | ( wire721  &  n_n216 ) ;
 assign wire2775 = ( n_n108  &  wire347 ) | ( n_n108  &  wire345 ) | ( n_n108  &  wire18956 ) ;
 assign wire18958 = ( n_n156  &  wire715 ) | ( wire721  &  n_n216 ) ;
 assign wire18959 = ( wire729  &  n_n156 ) | ( n_n156  &  wire717 ) | ( wire729  &  n_n149 ) | ( wire717  &  n_n149 ) ;
 assign wire2776 = ( n_n101  &  wire260 ) | ( n_n101  &  wire18958 ) | ( n_n101  &  wire18959 ) ;
 assign wire18944 = ( i_15_  &  n_n177  &  n_n213 ) | ( (~ i_15_)  &  n_n177  &  n_n213 ) | ( i_15_  &  n_n170  &  n_n213 ) | ( (~ i_15_)  &  n_n170  &  n_n213 ) ;
 assign wire18945 = ( i_9_  &  (~ i_10_)  &  i_11_  &  wire729 ) | ( (~ i_9_)  &  (~ i_10_)  &  i_11_  &  wire729 ) ;
 assign wire2785 = ( wire146  &  n_n125 ) | ( n_n125  &  wire183 ) | ( n_n125  &  wire18945 ) ;
 assign wire2791 = ( wire1244  &  wire1243 ) ;
 assign wire2797 = ( n_n220  &  n_n111  &  wire16987  &  wire412 ) ;
 assign wire2801 = ( n_n113  &  wire305 ) | ( n_n113  &  wire310 ) ;
 assign wire2802 = ( n_n112  &  wire318 ) | ( wire715  &  n_n191  &  n_n112 ) ;
 assign wire2808 = ( wire123  &  n_n123 ) | ( n_n123  &  wire175 ) ;
 assign wire2809 = ( wire133  &  n_n125 ) | ( wire729  &  n_n149  &  n_n125 ) ;
 assign wire2814 = ( wire146  &  n_n123 ) | ( wire729  &  n_n177  &  n_n123 ) ;
 assign wire2815 = ( n_n125  &  wire123 ) | ( n_n125  &  wire175 ) ;
 assign wire2817 = ( wire143  &  n_n123 ) | ( n_n123  &  wire364 ) ;
 assign wire2825 = ( wire143  &  n_n125 ) | ( n_n125  &  wire364 ) ;
 assign wire18921 = ( i_9_  &  i_10_  &  i_11_  &  wire721 ) | ( i_9_  &  (~ i_10_)  &  i_11_  &  wire721 ) | ( (~ i_9_)  &  (~ i_10_)  &  (~ i_11_)  &  wire721 ) ;
 assign wire2828 = ( n_n197  &  n_n137 ) | ( n_n197  &  wire302 ) | ( n_n197  &  wire18921 ) ;
 assign wire2831 = ( n_n197  &  wire303 ) | ( n_n197  &  wire321 ) ;
 assign wire2842 = ( n_n123  &  wire139 ) | ( n_n184  &  wire729  &  n_n123 ) ;
 assign wire2843 = ( n_n125  &  wire139 ) | ( n_n125  &  wire313 ) ;
 assign wire18894 = ( i_9_  &  (~ i_10_)  &  i_11_  &  wire729 ) | ( (~ i_9_)  &  (~ i_10_)  &  i_11_  &  wire729 ) ;
 assign wire2853 = ( n_n36  &  wire183 ) | ( n_n36  &  wire18894 ) ;
 assign wire2865 = ( n_n34  &  n_n89 ) | ( n_n34  &  wire139 ) | ( n_n34  &  wire313 ) ;
 assign wire2866 = ( wire146  &  n_n36 ) | ( n_n36  &  n_n89 ) | ( n_n36  &  wire383 ) ;
 assign wire2870 = ( n_n34  &  wire257 ) | ( n_n184  &  wire729  &  n_n34 ) ;
 assign wire18879 = ( i_9_  &  i_10_  &  (~ i_11_)  &  wire729 ) | ( (~ i_9_)  &  i_10_  &  (~ i_11_)  &  wire729 ) ;
 assign wire2875 = ( n_n34  &  n_n139 ) | ( n_n34  &  wire175 ) | ( n_n34  &  wire18879 ) ;
 assign wire2897 = ( n_n41  &  wire260 ) | ( n_n41  &  wire373 ) | ( n_n41  &  n_n141 ) ;
 assign wire18859 = ( wire729  &  n_n149 ) | ( wire715  &  n_n149 ) | ( wire717  &  n_n149 ) ;
 assign wire18852 = ( n_n177  &  wire715 ) | ( n_n177  &  wire716 ) ;
 assign wire2910 = ( n_n38  &  wire1128 ) | ( n_n38  &  wire18852 ) ;
 assign wire18847 = ( (~ i_9_)  &  (~ i_10_)  &  i_11_  &  wire721 ) | ( (~ i_9_)  &  i_10_  &  (~ i_11_)  &  wire721 ) ;
 assign wire2914 = ( n_n33  &  wire293 ) | ( n_n33  &  wire18847 ) ;
 assign wire2915 = ( n_n162  &  wire714  &  n_n157  &  wire197 ) ;
 assign wire2939 = ( n_n32  &  wire305 ) | ( n_n32  &  wire310 ) ;
 assign wire18824 = ( (~ i_9_)  &  (~ i_10_)  &  i_11_  &  wire715 ) | ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire715 ) ;
 assign wire2940 = ( n_n33  &  wire230 ) | ( n_n33  &  wire318 ) | ( n_n33  &  wire18824 ) ;
 assign wire18821 = ( wire729  &  n_n149 ) | ( wire715  &  n_n149 ) | ( wire717  &  n_n149 ) ;
 assign wire2943 = ( n_n33  &  wire347 ) | ( n_n33  &  wire352 ) | ( n_n33  &  wire18821 ) ;
 assign wire2944 = ( n_n184  &  wire715  &  n_n32 ) ;
 assign wire18810 = ( n_n159  &  n_n35  &  n_n111 ) | ( n_n159  &  n_n124  &  n_n111 ) ;
 assign wire2952 = ( n_n3  &  wire95 ) | ( wire95  &  wire18810 ) ;
 assign wire18811 = ( n_n159  &  n_n218  &  n_n35 ) | ( n_n159  &  n_n218  &  n_n124 ) ;
 assign wire2953 = ( wire729  &  n_n156  &  n_n12 ) | ( wire729  &  n_n156  &  wire18811 ) ;
 assign wire2958 = ( n_n9  &  wire95 ) | ( n_n6  &  wire95 ) | ( wire95  &  n_n12 ) ;
 assign wire2959 = ( n_n5  &  n_n71 ) | ( n_n71  &  n_n9 ) | ( n_n71  &  n_n6 ) ;
 assign wire2964 = ( n_n31  &  wire118 ) | ( n_n31  &  wire221 ) | ( n_n31  &  wire298 ) ;
 assign wire18784 = ( wire725  &  n_n156 ) | ( wire725  &  n_n177 ) | ( n_n156  &  wire721 ) ;
 assign wire2970 = ( n_n30  &  wire152 ) | ( n_n30  &  wire18784 ) ;
 assign wire2974 = ( n_n30  &  wire59 ) | ( n_n30  &  wire289 ) ;
 assign wire2975 = ( n_n31  &  wire115 ) | ( wire729  &  n_n31  &  n_n149 ) ;
 assign wire2979 = ( n_n30  &  wire172 ) | ( n_n30  &  wire209 ) ;
 assign wire18771 = ( wire725  &  n_n199 ) | ( wire725  &  n_n216 ) | ( wire721  &  n_n216 ) ;
 assign wire2981 = ( n_n31  &  wire218 ) | ( n_n31  &  wire212 ) | ( n_n31  &  wire18771 ) ;
 assign wire2995 = ( n_n33  &  wire63 ) | ( n_n33  &  wire52 ) | ( n_n33  &  wire222 ) ;
 assign wire3001 = ( n_n30  &  n_n95 ) | ( n_n30  &  wire111 ) | ( n_n30  &  wire341 ) ;
 assign wire3006 = ( n_n30  &  wire206 ) | ( n_n30  &  wire243 ) | ( n_n30  &  wire368 ) ;
 assign wire3013 = ( n_n162  &  n_n35  &  n_n220  &  wire860 ) ;
 assign wire18744 = ( n_n89 ) | ( wire93 ) | ( wire241 ) | ( wire54 ) ;
 assign wire3014 = ( n_n31  &  wire273 ) | ( n_n31  &  wire268 ) | ( n_n31  &  wire18744 ) ;
 assign wire3015 = ( n_n30  &  wire162 ) | ( n_n30  &  wire164 ) ;
 assign wire3044 = ( i_7_  &  i_6_  &  n_n162  &  n_n19 ) ;
 assign wire3059 = ( n_n162  &  n_n16  &  n_n19 ) | ( n_n16  &  n_n48  &  n_n19 ) ;
 assign wire3060 = ( n_n218  &  n_n19  &  n_n18 ) | ( n_n19  &  n_n111  &  n_n18 ) ;
 assign wire18696 = ( n_n159  &  n_n218  &  n_n35 ) | ( n_n159  &  n_n218  &  n_n124 ) ;
 assign wire3066 = ( wire344  &  wire815 ) | ( wire344  &  wire18696 ) ;
 assign wire3067 = ( n_n6  &  n_n68 ) | ( n_n68  &  wire398 ) | ( n_n68  &  wire815 ) ;
 assign wire3068 = ( n_n162  &  n_n124  &  n_n220  &  wire381 ) ;
 assign wire3069 = ( n_n162  &  n_n220  &  n_n161  &  wire172 ) ;
 assign wire3078 = ( n_n101  &  wire80 ) | ( n_n101  &  wire78 ) ;
 assign wire18687 = ( n_n156  &  wire719 ) | ( wire725  &  n_n170 ) ;
 assign wire3079 = ( wire381  &  n_n108 ) | ( n_n108  &  wire18687 ) ;
 assign wire3080 = ( n_n108  &  wire173 ) | ( n_n108  &  wire204 ) ;
 assign wire18686 = ( n_n156  &  wire719 ) | ( wire725  &  n_n149 ) ;
 assign wire3081 = ( wire245  &  n_n101 ) | ( n_n101  &  wire18686 ) ;
 assign wire3102 = ( n_n101  &  wire234 ) | ( n_n101  &  wire220 ) ;
 assign wire3111 = ( _2752 ) | ( n_n108  &  wire222 ) | ( n_n108  &  wire242 ) ;
 assign wire3113 = ( n_n101  &  wire155 ) | ( n_n101  &  wire205 ) | ( n_n101  &  wire215 ) ;
 assign wire3123 = ( n_n42  &  wire256 ) | ( n_n42  &  wire216 ) ;
 assign wire3124 = ( n_n43  &  wire130 ) | ( n_n43  &  n_n116 ) | ( n_n43  &  wire242 ) ;
 assign wire3135 = ( wire152  &  n_n212 ) | ( wire719  &  n_n149  &  n_n212 ) ;
 assign wire18617 = ( wire725  &  n_n156 ) | ( wire725  &  n_n149 ) | ( n_n149  &  wire721 ) ;
 assign wire3136 = ( wire157  &  n_n197 ) | ( n_n197  &  wire204 ) | ( n_n197  &  wire18617 ) ;
 assign wire18609 = ( wire725  &  n_n170 ) | ( wire725  &  n_n191 ) | ( wire721  &  n_n191 ) ;
 assign wire3142 = ( n_n197  &  wire252 ) | ( n_n197  &  wire171 ) | ( n_n197  &  wire18609 ) ;
 assign wire3143 = ( n_n17  &  n_n218  &  wire714  &  wire1655 ) ;
 assign wire3154 = ( n_n197  &  wire242 ) | ( n_n184  &  wire719  &  n_n197 ) ;
 assign wire3155 = ( n_n212  &  wire247 ) | ( n_n212  &  wire171 ) | ( n_n212  &  wire160 ) ;
 assign wire3195 = ( i_7_  &  i_6_  &  n_n159  &  n_n111 ) | ( i_7_  &  (~ i_6_)  &  n_n159  &  n_n111 ) ;
 assign wire3201 = ( wire168  &  n_n123 ) | ( n_n123  &  wire68 ) | ( n_n123  &  wire151 ) ;
 assign wire18529 = ( n_n177  &  wire719 ) | ( wire725  &  n_n170 ) ;
 assign wire3219 = ( wire252  &  n_n123 ) | ( n_n123  &  wire174 ) | ( n_n123  &  wire18529 ) ;
 assign wire3222 = ( n_n123  &  wire171 ) | ( n_n123  &  wire160 ) ;
 assign wire18528 = ( n_n184  &  wire725 ) | ( n_n177  &  wire719 ) ;
 assign wire3223 = ( n_n125  &  wire217 ) | ( n_n125  &  wire18528 ) ;
 assign wire3225 = ( wire132  &  n_n125 ) | ( wire149  &  n_n125 ) | ( wire126  &  n_n125 ) ;
 assign wire3229 = ( wire63  &  n_n123 ) | ( wire48  &  n_n123 ) | ( n_n123  &  wire129 ) ;
 assign wire3234 = ( n_n65  &  n_n2 ) | ( n_n2  &  n_n89 ) | ( n_n2  &  wire87 ) ;
 assign wire3244 = ( wire145  &  n_n3 ) | ( n_n3  &  n_n186 ) | ( n_n3  &  wire170 ) ;
 assign wire3245 = ( n_n4  &  wire185 ) | ( n_n4  &  wire270 ) ;
 assign wire3256 = ( n_n65  &  n_n9 ) | ( n_n9  &  n_n89 ) | ( n_n9  &  wire87 ) ;
 assign wire3257 = ( n_n10  &  n_n65 ) | ( n_n10  &  wire77 ) | ( n_n10  &  wire87 ) ;
 assign wire3258 = ( n_n41  &  wire1386 ) | ( n_n41  &  wire724  &  n_n216 ) ;
 assign wire3264 = ( _2990 ) | ( wire154  &  n_n40 ) | ( n_n40  &  wire124 ) ;
 assign wire3271 = ( wire143  &  n_n41 ) | ( wire154  &  n_n41 ) ;
 assign wire3275 = ( _3004 ) | ( n_n41  &  wire134 ) | ( n_n41  &  wire123 ) ;
 assign wire3279 = ( n_n40  &  wire198 ) | ( n_n40  &  wire289 ) ;
 assign wire18457 = ( n_n149  &  wire726 ) | ( n_n149  &  wire724 ) ;
 assign wire3280 = ( n_n41  &  wire127 ) | ( n_n41  &  wire133 ) | ( n_n41  &  wire18457 ) ;
 assign wire3312 = ( n_n46  &  wire111 ) | ( n_n46  &  wire341 ) ;
 assign wire18416 = ( wire729  &  n_n199 ) | ( wire723  &  n_n199 ) | ( wire727  &  n_n199 ) ;
 assign wire3313 = ( n_n47  &  wire206 ) | ( n_n47  &  wire243 ) | ( n_n47  &  wire18416 ) ;
 assign wire3325 = ( n_n46  &  n_n102 ) | ( n_n46  &  wire162 ) | ( n_n46  &  wire164 ) ;
 assign wire3337 = ( n_n47  &  wire256 ) | ( n_n47  &  wire216 ) ;
 assign wire18394 = ( n_n184  &  wire725 ) | ( wire719  &  n_n191 ) ;
 assign wire3338 = ( wire172  &  n_n46 ) | ( n_n46  &  wire217 ) | ( n_n46  &  wire18394 ) ;
 assign wire18386 = ( wire725  &  n_n199 ) | ( wire725  &  n_n216 ) | ( wire721  &  n_n216 ) ;
 assign wire3342 = ( n_n47  &  wire218 ) | ( n_n47  &  wire212 ) | ( n_n47  &  wire18386 ) ;
 assign wire3353 = ( n_n46  &  n_n77 ) | ( n_n46  &  wire117 ) | ( n_n46  &  wire281 ) ;
 assign wire3374 = ( wire185  &  wire1427 ) | ( wire270  &  wire1427 ) | ( wire1427  &  wire372 ) ;
 assign wire3375 = ( wire270  &  n_n3 ) | ( n_n3  &  wire372 ) ;
 assign wire3385 = ( n_n43  &  n_n138 ) | ( n_n43  &  wire62 ) | ( n_n43  &  wire272 ) ;
 assign wire3392 = ( n_n43  &  wire211 ) | ( n_n43  &  wire107 ) ;
 assign wire3397 = ( wire172  &  n_n43 ) | ( n_n43  &  wire216 ) ;
 assign wire3404 = ( n_n42  &  wire211 ) | ( n_n42  &  wire107 ) | ( n_n42  &  wire272 ) ;
 assign wire3409 = ( wire48  &  n_n112 ) | ( wire52  &  n_n112 ) | ( wire129  &  n_n112 ) ;
 assign wire3415 = ( n_n5  &  wire145 ) | ( n_n5  &  n_n151 ) | ( n_n5  &  wire370 ) ;
 assign wire3425 = ( n_n4  &  wire185 ) | ( n_n4  &  wire87 ) ;
 assign wire3435 = ( i_7_  &  i_6_  &  n_n159  &  n_n111 ) ;
 assign wire3437 = ( n_n9  &  wire145 ) | ( n_n9  &  n_n186 ) | ( n_n9  &  wire170 ) ;
 assign wire3438 = ( n_n10  &  n_n144 ) | ( n_n10  &  n_n186 ) | ( n_n10  &  wire170 ) ;
 assign wire3471 = ( n_n40  &  wire198 ) | ( n_n40  &  wire289 ) ;
 assign wire3479 = ( n_n40  &  wire116 ) | ( wire729  &  n_n156  &  n_n40 ) ;
 assign wire3498 = ( n_n41  &  wire256 ) | ( n_n41  &  wire216 ) ;
 assign wire3515 = ( n_n48  &  n_n220  &  n_n200  &  wire1459 ) ;
 assign wire18260 = ( n_n77 ) | ( wire117 ) | ( wire281 ) | ( wire59 ) ;
 assign wire3516 = ( n_n41  &  wire294 ) | ( n_n41  &  wire289 ) | ( n_n41  &  wire18260 ) ;
 assign wire3520 = ( _3332 ) | ( n_n40  &  wire241 ) | ( n_n40  &  wire94 ) ;
 assign wire3524 = ( n_n41  &  wire179 ) | ( n_n41  &  wire324 ) | ( n_n41  &  wire104 ) ;
 assign wire3526 = ( n_n41  &  wire243 ) | ( wire729  &  n_n41  &  n_n199 ) ;
 assign wire3531 = ( n_n41  &  wire81 ) | ( n_n41  &  wire206 ) | ( n_n41  &  wire368 ) ;
 assign wire3533 = ( n_n41  &  wire162 ) | ( n_n41  &  wire341 ) | ( n_n41  &  wire399 ) ;
 assign wire3550 = ( n_n40  &  wire144 ) | ( n_n40  &  wire122 ) ;
 assign wire3551 = ( wire725  &  n_n149  &  n_n41 ) ;
 assign wire3563 = ( wire158  &  n_n46 ) | ( wire133  &  n_n46 ) ;
 assign wire18194 = ( wire725  &  n_n170 ) | ( wire725  &  n_n191 ) | ( wire721  &  n_n191 ) ;
 assign wire3570 = ( n_n46  &  wire252 ) | ( n_n46  &  wire171 ) | ( n_n46  &  wire18194 ) ;
 assign wire3575 = ( n_n46  &  wire153 ) | ( n_n46  &  wire135 ) | ( n_n46  &  wire125 ) ;
 assign wire3580 = ( n_n47  &  wire171 ) | ( n_n47  &  wire160 ) ;
 assign wire18188 = ( n_n184  &  wire719 ) | ( wire725  &  n_n216 ) ;
 assign wire3581 = ( n_n46  &  wire242 ) | ( n_n46  &  wire18188 ) ;
 assign wire3588 = ( n_n47  &  wire52 ) | ( n_n47  &  wire139 ) | ( n_n47  &  wire128 ) ;
 assign wire3607 = ( n_n48  &  wire714  &  wire152  &  n_n18 ) ;
 assign wire3621 = ( wire253  &  n_n6 ) | ( wire253  &  wire398 ) | ( wire253  &  wire1550 ) ;
 assign wire18157 = ( n_n159  &  n_n218  &  n_n35 ) | ( n_n159  &  n_n218  &  n_n124 ) ;
 assign wire3622 = ( n_n156  &  wire717  &  wire1550 ) | ( n_n156  &  wire717  &  wire18157 ) ;
 assign wire3624 = ( n_n162  &  n_n19  &  n_n157 ) | ( n_n48  &  n_n19  &  n_n157 ) ;
 assign wire3643 = ( n_n212  &  wire74 ) | ( n_n212  &  wire68 ) ;
 assign wire18117 = ( n_n148 ) | ( wire90 ) | ( wire69 ) | ( wire225 ) ;
 assign wire3653 = ( n_n125  &  wire205 ) | ( n_n125  &  wire84 ) | ( n_n125  &  wire18117 ) ;
 assign wire18111 = ( n_n176 ) | ( wire62 ) | ( wire107 ) | ( wire18107 ) ;
 assign wire18102 = ( wire234 ) | ( wire220 ) ;
 assign wire18103 = ( wire60 ) | ( wire242 ) | ( n_n184  &  wire719 ) ;
 assign wire18104 = ( wire218 ) | ( wire171 ) | ( wire160 ) | ( wire18098 ) ;
 assign wire3662 = ( n_n125  &  wire18102 ) | ( n_n125  &  wire18103 ) | ( n_n125  &  wire18104 ) ;
 assign wire18092 = ( (~ i_9_)  &  i_10_  &  i_11_  &  wire720 ) | ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire720 ) ;
 assign wire3665 = ( n_n125  &  wire219 ) | ( n_n125  &  wire70 ) | ( n_n125  &  wire18092 ) ;
 assign wire18087 = ( wire127 ) | ( wire153 ) | ( wire719  &  n_n191 ) ;
 assign wire18088 = ( wire172 ) | ( wire133 ) | ( n_n63 ) | ( wire135 ) ;
 assign wire3671 = ( n_n212  &  wire18087 ) | ( n_n212  &  wire18088 ) ;
 assign wire3676 = ( _3637 ) | ( _3638 ) | ( _3639 ) ;
 assign wire18067 = ( _30765 ) | ( wire719  &  _29117 ) | ( wire719  &  _30347 ) ;
 assign wire18068 = ( _30763 ) | ( wire725  &  _28911 ) | ( wire725  &  _29613 ) ;
 assign wire18069 = ( wire172 ) | ( wire150 ) | ( wire217 ) | ( wire173 ) ;
 assign wire3685 = ( n_n108  &  wire18067 ) | ( n_n108  &  wire18068 ) | ( n_n108  &  wire18069 ) ;
 assign wire18053 = ( n_n184  &  wire729 ) | ( n_n184  &  wire719 ) | ( n_n184  &  wire728 ) ;
 assign wire3690 = ( n_n113  &  wire94 ) | ( n_n113  &  wire184 ) | ( n_n113  &  wire18053 ) ;
 assign wire3696 = ( n_n220  &  n_n111  &  wire16987  &  wire1747 ) ;
 assign wire3700 = ( n_n113  &  wire268 ) | ( n_n113  &  wire54 ) ;
 assign wire3701 = ( wire245  &  n_n125 ) | ( wire725  &  n_n149  &  n_n125 ) ;
 assign wire3702 = ( n_n47  &  wire139 ) | ( n_n47  &  wire128 ) ;
 assign wire3710 = ( n_n220  &  n_n111  &  wire17072  &  wire412 ) ;
 assign wire3723 = ( n_n39  &  wire53 ) | ( n_n39  &  n_n143 ) | ( n_n39  &  wire237 ) ;
 assign wire3747 = ( n_n41  &  wire225 ) | ( n_n170  &  wire720  &  n_n41 ) ;
 assign wire17993 = ( wire62 ) | ( wire240 ) | ( wire107 ) | ( wire17989 ) ;
 assign wire3755 = ( n_n41  &  wire211 ) | ( n_n41  &  wire272 ) | ( n_n41  &  wire17993 ) ;
 assign wire3759 = ( n_n43  &  wire256 ) | ( n_n43  &  wire216 ) ;
 assign wire3773 = ( _3809 ) | ( _3810 ) | ( _3811 ) ;
 assign wire3774 = ( n_n220  &  n_n111  &  n_n149  &  n_n126 ) ;
 assign wire3810 = ( n_n32  &  wire107 ) | ( n_n184  &  wire720  &  n_n32 ) ;
 assign wire17940 = ( wire78 ) | ( wire217 ) | ( wire719  &  n_n170 ) ;
 assign wire17941 = ( _30861 ) | ( wire725  &  _28911 ) | ( wire725  &  _29613 ) ;
 assign wire17942 = ( wire157 ) | ( wire172 ) | ( wire150 ) | ( wire173 ) ;
 assign wire3811 = ( n_n36  &  wire17940 ) | ( n_n36  &  wire17941 ) | ( n_n36  &  wire17942 ) ;
 assign wire3828 = ( n_n36  &  wire152 ) | ( wire719  &  n_n149  &  n_n36 ) ;
 assign wire17909 = ( wire725  &  n_n156 ) | ( wire725  &  n_n149 ) | ( n_n149  &  wire721 ) ;
 assign wire3829 = ( wire157  &  n_n34 ) | ( n_n34  &  wire204 ) | ( n_n34  &  wire17909 ) ;
 assign wire17901 = ( wire725  &  n_n170 ) | ( wire725  &  n_n191 ) | ( wire721  &  n_n191 ) ;
 assign wire3835 = ( n_n34  &  wire252 ) | ( n_n34  &  wire171 ) | ( n_n34  &  wire17901 ) ;
 assign wire3836 = ( n_n218  &  wire714  &  n_n157  &  wire1814 ) ;
 assign wire3850 = ( n_n34  &  wire242 ) | ( n_n184  &  wire719  &  n_n34 ) ;
 assign wire3851 = ( n_n36  &  wire247 ) | ( n_n36  &  wire171 ) | ( n_n36  &  wire160 ) ;
 assign wire3866 = ( wire132  &  n_n34 ) | ( n_n34  &  wire149 ) | ( n_n34  &  wire46 ) ;
 assign wire3886 = ( _3948 ) | ( n_n111  &  _30568  &  _30569 ) ;
 assign wire3887 = ( i_7_  &  i_6_  &  n_n162  &  n_n19 ) | ( i_7_  &  (~ i_6_)  &  n_n162  &  n_n19 ) ;
 assign wire3895 = ( n_n4  &  wire145 ) | ( n_n5  &  wire145 ) | ( n_n6  &  wire145 ) ;
 assign wire3896 = ( n_n5  &  n_n186 ) | ( n_n9  &  n_n186 ) | ( n_n6  &  n_n186 ) ;
 assign wire3897 = ( n_n4  &  wire717  &  n_n191 ) | ( wire717  &  n_n191  &  wire1044 ) ;
 assign wire3899 = ( (~ i_7_)  &  i_6_  &  n_n159  &  _30595 ) | ( i_7_  &  (~ i_6_)  &  n_n159  &  _30595 ) ;
 assign wire3900 = ( n_n10  &  wire145 ) | ( n_n9  &  wire145 ) | ( wire145  &  n_n12 ) ;
 assign wire3901 = ( n_n10  &  n_n186 ) | ( n_n14  &  n_n186 ) | ( n_n186  &  n_n12 ) ;
 assign wire3957 = ( n_n36  &  wire172 ) | ( n_n36  &  wire80 ) | ( n_n36  &  wire78 ) ;
 assign wire17808 = ( wire725  &  n_n156 ) | ( n_n156  &  wire721 ) | ( wire725  &  n_n191 ) ;
 assign wire3958 = ( n_n34  &  wire144 ) | ( n_n34  &  wire222 ) | ( n_n34  &  wire17808 ) ;
 assign wire3964 = ( n_n34  &  wire214 ) | ( n_n34  &  wire212 ) ;
 assign wire3973 = ( n_n30  &  wire146 ) | ( n_n30  &  wire52 ) | ( n_n30  &  wire129 ) ;
 assign wire3990 = ( n_n31  &  wire157 ) | ( n_n31  &  wire80 ) | ( n_n31  &  wire78 ) ;
 assign wire17781 = ( n_n177  &  wire719 ) | ( wire725  &  n_n191 ) ;
 assign wire3991 = ( n_n30  &  wire174 ) | ( n_n30  &  wire222 ) | ( n_n30  &  wire17781 ) ;
 assign wire3996 = ( n_n30  &  wire214 ) | ( n_n30  &  wire212 ) ;
 assign wire3998 = ( wire143  &  n_n197 ) | ( wire154  &  n_n197 ) ;
 assign wire4013 = ( n_n125  &  wire86 ) | ( n_n125  &  wire180 ) | ( n_n125  &  n_n190 ) ;
 assign wire4020 = ( wire172  &  n_n212 ) | ( wire719  &  n_n191  &  n_n212 ) ;
 assign wire4021 = ( n_n197  &  wire214 ) | ( n_n197  &  wire212 ) ;
 assign wire4026 = ( n_n212  &  wire80 ) | ( n_n212  &  wire78 ) ;
 assign wire4027 = ( wire144  &  n_n197 ) | ( n_n197  &  n_n59 ) | ( n_n197  &  wire222 ) ;
 assign wire17739 = ( n_n155 ) | ( wire224 ) | ( wire250 ) | ( wire57 ) ;
 assign wire4043 = ( wire215  &  n_n123 ) | ( n_n123  &  wire100 ) | ( n_n123  &  wire17739 ) ;
 assign wire4048 = ( wire172  &  n_n123 ) | ( n_n138  &  n_n123 ) | ( n_n123  &  wire125 ) ;
 assign wire4064 = ( wire80  &  n_n123 ) | ( wire78  &  n_n123 ) ;
 assign wire4065 = ( wire381  &  n_n125 ) | ( n_n156  &  wire719  &  n_n125 ) ;
 assign wire4080 = ( wire143  &  n_n46 ) | ( wire154  &  n_n46 ) ;
 assign wire4088 = ( n_n46  &  wire52 ) | ( n_n46  &  wire129 ) ;
 assign wire4102 = ( n_n42  &  wire52 ) | ( n_n42  &  wire129 ) ;
 assign wire4103 = ( n_n162  &  wire714  &  n_n18  &  wire222 ) ;
 assign wire4104 = ( n_n41  &  wire381 ) | ( n_n41  &  wire171 ) | ( n_n41  &  wire160 ) ;
 assign wire4113 = ( n_n40  &  wire215 ) | ( n_n40  &  n_n155 ) | ( n_n40  &  wire125 ) ;
 assign wire4130 = ( n_n42  &  wire171 ) | ( n_n42  &  wire160 ) ;
 assign wire4143 = ( n_n40  &  n_n176 ) | ( n_n40  &  wire250 ) | ( n_n40  &  wire100 ) ;
 assign wire4151 = ( n_n17  &  n_n48  &  wire714  &  wire240 ) ;
 assign wire17632 = ( wire725  &  n_n156 ) | ( n_n156  &  wire721 ) | ( wire725  &  n_n191 ) ;
 assign wire4158 = ( wire144  &  n_n46 ) | ( n_n46  &  wire222 ) | ( n_n46  &  wire17632 ) ;
 assign wire4159 = ( n_n124  &  n_n220  &  n_n156  &  n_n111 ) ;
 assign wire4172 = ( wire172  &  n_n108 ) | ( n_n138  &  n_n108 ) | ( n_n108  &  wire78 ) ;
 assign wire4185 = ( n_n108  &  wire125 ) | ( wire725  &  n_n216  &  n_n108 ) ;
 assign wire4217 = ( n_n4  &  wire170 ) | ( n_n5  &  wire170 ) | ( n_n6  &  wire170 ) ;
 assign wire17591 = ( (~ i_7_)  &  (~ i_5_)  &  i_6_ ) | ( i_7_  &  (~ i_5_)  &  (~ i_6_) ) ;
 assign wire4220 = ( i_3_  &  i_4_  &  n_n159  &  wire17591 ) ;
 assign wire4221 = ( n_n4  &  wire717  &  n_n149 ) | ( wire717  &  n_n149  &  wire1527 ) ;
 assign wire4228 = ( n_n10  &  wire170 ) | ( n_n9  &  wire170 ) | ( n_n12  &  wire170 ) ;
 assign wire4229 = ( n_n10  &  n_n144 ) | ( n_n14  &  n_n144 ) | ( n_n144  &  n_n12 ) ;
 assign wire4230 = ( n_n218  &  n_n220  &  n_n200  &  wire123 ) ;
 assign wire17569 = ( n_n156  &  wire719 ) | ( wire719  &  n_n149 ) | ( n_n156  &  wire728 ) ;
 assign wire4233 = ( wire152  &  n_n197 ) | ( n_n197  &  wire17569 ) ;
 assign wire17570 = ( wire725  &  n_n156 ) | ( wire725  &  n_n149 ) | ( n_n156  &  wire721 ) ;
 assign wire4234 = ( wire245  &  n_n212 ) | ( wire144  &  n_n212 ) | ( n_n212  &  wire17570 ) ;
 assign wire4252 = ( n_n220  &  n_n111  &  n_n149  &  n_n126 ) ;
 assign wire4253 = ( n_n124  &  n_n220  &  n_n156  &  n_n111 ) ;
 assign wire4263 = ( n_n124  &  n_n48  &  n_n220  &  wire249 ) ;
 assign wire4285 = ( n_n40  &  wire173 ) | ( n_n40  &  wire204 ) ;
 assign wire17535 = ( wire725  &  n_n156 ) | ( wire719  &  n_n149 ) ;
 assign wire4286 = ( wire157  &  n_n41 ) | ( wire152  &  n_n41 ) | ( n_n41  &  wire17535 ) ;
 assign wire4291 = ( n_n40  &  wire215 ) | ( n_n156  &  wire720  &  n_n40 ) ;
 assign wire4323 = ( n_n123  &  wire173 ) | ( n_n123  &  wire204 ) ;
 assign wire17468 = ( wire725  &  n_n156 ) | ( wire719  &  n_n149 ) ;
 assign wire4324 = ( wire152  &  n_n125 ) | ( n_n125  &  wire17468 ) ;
 assign wire4343 = ( wire152  &  n_n108 ) | ( wire719  &  n_n149  &  n_n108 ) ;
 assign wire17480 = ( wire725  &  n_n156 ) | ( wire725  &  n_n149 ) | ( n_n149  &  wire721 ) ;
 assign wire4344 = ( wire157  &  n_n101 ) | ( n_n101  &  wire17480 ) ;
 assign wire4382 = ( n_n125  &  wire215 ) | ( n_n156  &  wire720  &  n_n125 ) ;
 assign wire17447 = ( n_n156  &  wire719 ) | ( wire719  &  n_n149 ) | ( n_n156  &  wire728 ) ;
 assign wire4395 = ( n_n34  &  wire152 ) | ( n_n34  &  wire17447 ) ;
 assign wire17448 = ( wire725  &  n_n156 ) | ( wire725  &  n_n149 ) | ( n_n156  &  wire721 ) ;
 assign wire4396 = ( n_n36  &  wire245 ) | ( n_n36  &  wire144 ) | ( n_n36  &  wire17448 ) ;
 assign wire17428 = ( wire725  &  n_n156 ) | ( n_n156  &  wire721 ) | ( wire725  &  n_n216 ) ;
 assign wire4419 = ( n_n30  &  wire152 ) | ( n_n30  &  wire125 ) | ( n_n30  &  wire17428 ) ;
 assign wire4427 = ( n_n31  &  wire245 ) | ( wire725  &  n_n31  &  n_n149 ) ;
 assign wire4429 = ( n_n31  &  wire55 ) | ( n_n31  &  wire127 ) | ( n_n31  &  wire133 ) ;
 assign wire17391 = ( i_15_  &  n_n211  &  n_n191 ) | ( (~ i_15_)  &  n_n211  &  n_n191 ) | ( (~ i_15_)  &  n_n191  &  n_n201 ) ;
 assign wire4453 = ( wire93  &  n_n123 ) | ( n_n123  &  wire177 ) | ( n_n123  &  wire17391 ) ;
 assign wire4454 = ( wire93  &  n_n125 ) | ( n_n125  &  wire362 ) | ( n_n125  &  wire17391 ) ;
 assign wire4458 = ( n_n123  &  wire94 ) | ( n_n184  &  wire729  &  n_n123 ) ;
 assign wire4459 = ( n_n125  &  wire94 ) | ( n_n125  &  wire177 ) ;
 assign wire17385 = ( i_9_  &  (~ i_10_)  &  i_11_  &  wire725 ) | ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire725 ) | ( (~ i_9_)  &  (~ i_10_)  &  (~ i_11_)  &  wire725 ) ;
 assign wire4470 = ( n_n125  &  wire164 ) | ( n_n125  &  wire358 ) ;
 assign wire4474 = ( n_n212  &  wire306 ) | ( n_n212  &  wire193 ) | ( n_n212  &  wire196 ) ;
 assign wire4475 = ( n_n197  &  wire168 ) | ( n_n197  &  wire193 ) | ( n_n197  &  wire196 ) ;
 assign wire4491 = ( n_n101  &  n_n210 ) | ( n_n101  &  wire374 ) | ( n_n101  &  wire17361 ) ;
 assign wire4496 = ( n_n108  &  wire307 ) | ( wire722  &  n_n191  &  n_n108 ) ;
 assign wire17357 = ( (~ i_9_)  &  (~ i_10_)  &  i_11_  &  wire722 ) | ( i_9_  &  i_10_  &  (~ i_11_)  &  wire722 ) ;
 assign wire4500 = ( n_n108  &  wire69 ) | ( n_n108  &  wire229 ) | ( n_n108  &  wire17357 ) ;
 assign wire4504 = ( n_n108  &  wire90 ) | ( n_n108  &  wire377 ) ;
 assign wire17349 = ( (~ i_9_)  &  (~ i_10_)  &  i_11_  &  wire722 ) | ( (~ i_9_)  &  (~ i_10_)  &  (~ i_11_)  &  wire722 ) ;
 assign wire17350 = ( n_n184  &  wire729 ) | ( wire729  &  n_n191 ) | ( n_n184  &  wire726 ) | ( n_n191  &  wire726 ) ;
 assign wire17352 = ( i_9_  &  (~ i_10_)  &  i_11_  &  wire722 ) | ( (~ i_9_)  &  (~ i_10_)  &  (~ i_11_)  &  wire722 ) ;
 assign wire17353 = ( wire729  &  n_n177 ) | ( wire729  &  n_n191 ) | ( n_n177  &  wire726 ) | ( n_n191  &  wire726 ) ;
 assign wire17343 = ( wire729  &  n_n170 ) | ( wire729  &  n_n191 ) | ( n_n170  &  wire726 ) | ( n_n191  &  wire726 ) ;
 assign wire4510 = ( n_n40  &  n_n168 ) | ( n_n40  &  wire229 ) | ( n_n40  &  wire17343 ) ;
 assign wire4520 = ( n_n41  &  wire307 ) | ( wire722  &  n_n41  &  n_n191 ) ;
 assign wire17336 = ( wire729  &  n_n177 ) | ( n_n177  &  wire722 ) | ( n_n177  &  wire726 ) ;
 assign wire4523 = ( n_n40  &  wire265 ) | ( n_n40  &  wire17336 ) ;
 assign wire4526 = ( n_n41  &  n_n196 ) | ( n_n41  &  wire374 ) | ( n_n41  &  wire263 ) ;
 assign wire17324 = ( i_9_  &  (~ i_10_)  &  i_11_  &  wire729 ) | ( (~ i_9_)  &  (~ i_10_)  &  i_11_  &  wire729 ) ;
 assign wire4539 = ( n_n36  &  wire117 ) | ( n_n36  &  wire366 ) | ( n_n36  &  wire17324 ) ;
 assign wire17317 = ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire729 ) | ( (~ i_9_)  &  (~ i_10_)  &  (~ i_11_)  &  wire729 ) ;
 assign wire4544 = ( n_n34  &  wire93 ) | ( n_n34  &  wire301 ) | ( n_n34  &  wire17317 ) ;
 assign wire17319 = ( i_15_  &  n_n184  &  n_n211 ) | ( (~ i_15_)  &  n_n184  &  n_n211 ) | ( i_15_  &  n_n211  &  n_n177 ) | ( (~ i_15_)  &  n_n211  &  n_n177 ) ;
 assign wire4545 = ( n_n36  &  wire120 ) | ( n_n36  &  wire94 ) | ( n_n36  &  wire17319 ) ;
 assign wire4548 = ( n_n34  &  wire94 ) | ( n_n34  &  wire177 ) ;
 assign wire4549 = ( n_n36  &  wire93 ) | ( wire729  &  n_n36  &  n_n191 ) ;
 assign wire4550 = ( n_n34  &  wire369 ) | ( wire729  &  n_n177  &  n_n34 ) ;
 assign wire4551 = ( n_n36  &  wire116 ) | ( n_n36  &  wire371 ) ;
 assign wire17310 = ( i_9_  &  i_10_  &  (~ i_11_)  &  wire729 ) | ( (~ i_9_)  &  i_10_  &  (~ i_11_)  &  wire729 ) ;
 assign wire4568 = ( n_n36  &  wire164 ) | ( n_n36  &  wire358 ) ;
 assign wire4569 = ( n_n34  &  n_n199  &  _29782 ) | ( n_n34  &  n_n199  &  _29784 ) ;
 assign wire17292 = ( wire722  &  n_n149 ) | ( wire725  &  n_n216 ) ;
 assign wire4572 = ( n_n41  &  wire60 ) | ( n_n41  &  wire351 ) | ( n_n41  &  wire17292 ) ;
 assign wire17294 = ( n_n156  &  wire722 ) | ( wire725  &  n_n216 ) ;
 assign wire17295 = ( wire729  &  n_n156 ) | ( wire729  &  n_n149 ) | ( n_n156  &  wire726 ) | ( n_n149  &  wire726 ) ;
 assign wire4573 = ( n_n40  &  wire377 ) | ( n_n40  &  wire17294 ) | ( n_n40  &  wire17295 ) ;
 assign wire4576 = ( n_n40  &  wire351 ) | ( wire722  &  n_n149  &  n_n40 ) ;
 assign wire17287 = ( n_n177  &  wire722 ) | ( n_n177  &  wire724 ) ;
 assign wire4581 = ( n_n38  &  wire1120 ) | ( n_n38  &  wire17287 ) ;
 assign wire4591 = ( n_n48  &  n_n220  &  n_n126  &  wire1116 ) ;
 assign wire4602 = ( wire120  &  n_n123 ) | ( wire729  &  n_n177  &  n_n123 ) ;
 assign wire4628 = ( n_n30  &  wire149 ) | ( n_n30  &  wire200 ) | ( n_n30  &  wire201 ) ;
 assign wire4638 = ( n_n31  &  wire176 ) | ( n_n31  &  n_n59 ) | ( n_n31  &  wire299 ) ;
 assign wire4639 = ( _5289 ) | ( n_n30  &  wire158 ) | ( n_n30  &  wire308 ) ;
 assign wire4644 = ( n_n31  &  wire130 ) | ( n_n31  &  wire304 ) | ( n_n31  &  wire306 ) ;
 assign wire4649 = ( n_n32  &  wire62 ) | ( n_n32  &  wire202 ) ;
 assign wire17224 = ( (~ i_9_)  &  (~ i_10_)  &  i_11_  &  wire722 ) | ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire722 ) ;
 assign wire4651 = ( n_n33  &  wire229 ) | ( n_n33  &  wire307 ) | ( n_n33  &  wire17224 ) ;
 assign wire4655 = ( n_n33  &  n_n147 ) | ( n_n33  &  wire351 ) | ( n_n33  &  wire69 ) ;
 assign wire17215 = ( (~ i_9_)  &  i_10_  &  (~ i_11_)  &  wire725 ) | ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire725 ) ;
 assign wire4662 = ( wire149  &  n_n46 ) | ( n_n46  &  wire200 ) | ( n_n46  &  wire201 ) ;
 assign wire4663 = ( wire131  &  n_n47 ) | ( n_n47  &  wire308 ) | ( n_n47  &  wire201 ) ;
 assign wire4669 = ( wire896  &  wire301 ) | ( n_n184  &  wire729  &  wire896 ) ;
 assign wire4671 = ( n_n43  &  wire94 ) | ( n_n43  &  wire177 ) ;
 assign wire4676 = ( n_n42  &  wire94 ) | ( n_n42  &  wire177 ) ;
 assign wire4684 = ( n_n47  &  wire168 ) | ( n_n47  &  wire193 ) | ( n_n47  &  wire196 ) ;
 assign wire4685 = ( n_n46  &  wire193 ) | ( n_n46  &  wire196 ) ;
 assign wire4735 = ( n_n101  &  wire100 ) | ( n_n177  &  wire720  &  n_n101 ) ;
 assign wire4743 = ( n_n123  &  wire224 ) | ( n_n123  &  wire250 ) | ( n_n123  &  wire57 ) ;
 assign wire4750 = ( n_n123  &  wire141 ) | ( wire719  &  n_n216  &  n_n123 ) ;
 assign wire4752 = ( n_n125  &  wire225 ) | ( n_n170  &  wire720  &  n_n125 ) ;
 assign wire4753 = ( _5601 ) | ( n_n123  &  wire225 ) | ( n_n123  &  wire100 ) ;
 assign wire4765 = ( wire85  &  n_n123 ) | ( wire720  &  n_n216  &  n_n123 ) ;
 assign wire4768 = ( n_n123  &  wire218 ) | ( wire725  &  n_n199  &  n_n123 ) ;
 assign wire4780 = ( n_n218  &  n_n220  &  n_n126  &  wire219 ) ;
 assign wire4786 = ( n_n17  &  n_n218  &  wire714  &  wire247 ) ;
 assign wire4805 = ( n_n46  &  wire86 ) | ( n_n46  &  wire208 ) | ( n_n46  &  wire148 ) ;
 assign wire4818 = ( n_n48  &  wire714  &  n_n18  &  wire1030 ) ;
 assign wire17089 = ( n_n176 ) | ( wire69 ) | ( wire224 ) | ( wire250 ) ;
 assign wire4819 = ( n_n46  &  wire225 ) | ( n_n46  &  wire100 ) | ( n_n46  &  wire17089 ) ;
 assign wire4820 = ( n_n47  &  wire85 ) | ( wire720  &  n_n47  &  n_n216 ) ;
 assign wire4821 = ( n_n108  &  wire150 ) | ( wire719  &  n_n170  &  n_n108 ) ;
 assign wire17074 = ( wire725  &  n_n177 ) | ( wire725  &  n_n170 ) | ( n_n170  &  wire721 ) ;
 assign wire4822 = ( n_n101  &  wire182 ) | ( n_n101  &  wire17074 ) ;
 assign wire4827 = ( n_n220  &  n_n177  &  n_n111  &  n_n200 ) ;
 assign wire4828 = ( n_n220  &  n_n170  &  n_n111  &  wire17072 ) ;
 assign wire4831 = ( n_n101  &  wire224 ) | ( n_n101  &  wire209 ) ;
 assign wire4832 = ( n_n57  &  n_n108 ) | ( n_n108  &  wire182 ) | ( n_n108  &  wire141 ) ;
 assign wire4838 = ( n_n162  &  n_n124  &  n_n220  &  wire1862 ) ;
 assign wire4839 = ( n_n108  &  wire153 ) | ( n_n108  &  wire135 ) ;
 assign wire4857 = ( n_n47  &  wire182 ) | ( wire725  &  n_n177  &  n_n47 ) ;
 assign wire4858 = ( wire719  &  n_n170  &  _29269 ) | ( n_n170  &  wire728  &  _29269 ) ;
 assign wire4859 = ( n_n47  &  wire153 ) | ( n_n47  &  wire135 ) ;
 assign wire17052 = ( wire725  &  n_n199 ) | ( wire719  &  n_n216 ) ;
 assign wire4860 = ( n_n46  &  wire141 ) | ( n_n46  &  wire17052 ) ;
 assign wire4863 = ( n_n38  &  wire53 ) | ( n_n38  &  wire237 ) ;
 assign wire4888 = ( n_n218  &  wire714  &  n_n157  &  wire151 ) ;
 assign wire4890 = ( n_n41  &  wire225 ) | ( n_n170  &  wire720  &  n_n41 ) ;
 assign wire4891 = ( n_n40  &  wire69 ) | ( n_n40  &  wire250 ) | ( n_n40  &  wire100 ) ;
 assign wire4900 = ( n_n17  &  n_n48  &  wire714  &  wire150 ) ;
 assign wire4904 = ( n_n40  &  wire141 ) | ( wire719  &  n_n40  &  n_n216 ) ;
 assign wire4905 = ( wire725  &  n_n199  &  _29181 ) | ( wire721  &  n_n199  &  _29181 ) ;
 assign wire4908 = ( n_n40  &  wire218 ) | ( wire725  &  n_n40  &  n_n199 ) ;
 assign wire4919 = ( n_n40  &  wire219 ) | ( wire720  &  n_n40  &  n_n199 ) ;
 assign wire4924 = ( n_n108  &  wire100 ) | ( n_n177  &  wire720  &  n_n108 ) ;
 assign wire4933 = ( n_n108  &  wire224 ) | ( n_n108  &  wire57 ) ;
 assign wire4937 = ( n_n101  &  wire219 ) | ( n_n101  &  wire108 ) ;
 assign wire4941 = ( n_n125  &  wire150 ) | ( wire719  &  n_n170  &  n_n125 ) ;
 assign wire16988 = ( wire725  &  n_n177 ) | ( wire725  &  n_n170 ) | ( n_n170  &  wire721 ) ;
 assign wire4942 = ( n_n123  &  wire182 ) | ( n_n123  &  wire209 ) | ( n_n123  &  wire16988 ) ;
 assign wire4950 = ( n_n220  &  n_n111  &  n_n199  &  wire16987 ) ;
 assign wire16972 = ( wire149 ) | ( wire147 ) | ( wire80 ) | ( wire78 ) ;
 assign wire4953 = ( n_n30  &  wire126 ) | ( n_n30  &  wire150 ) | ( n_n30  &  wire16972 ) ;
 assign wire16964 = ( wire719  &  n_n170 ) | ( wire725  &  n_n216 ) ;
 assign wire4961 = ( n_n30  &  wire146 ) | ( n_n30  &  wire125 ) | ( n_n30  &  wire16964 ) ;
 assign wire16946 = ( n_n177  &  wire719 ) | ( wire719  &  n_n170 ) | ( n_n177  &  wire728 ) ;
 assign wire4982 = ( n_n218  &  wire714  &  n_n157  &  wire942 ) ;
 assign wire4986 = ( n_n218  &  wire714  &  n_n157  &  wire247 ) ;
 assign wire16940 = ( wire69 ) | ( wire186 ) | ( wire208 ) | ( wire16936 ) ;
 assign wire4993 = ( n_n33  &  wire225 ) | ( n_n33  &  wire148 ) | ( n_n33  &  wire16940 ) ;
 assign wire4998 = ( n_n124  &  n_n48  &  n_n220  &  wire140 ) ;
 assign wire16908 = ( n_n159  &  n_n35  &  n_n48 ) | ( n_n159  &  n_n35  &  n_n111 ) ;
 assign wire16909 = ( n_n159  &  n_n218  &  n_n35 ) | ( n_n159  &  n_n218  &  n_n124 ) ;
 assign wire5067 = ( n_n184  &  wire725  &  n_n111 ) ;
 assign wire5068 = ( n_n184  &  n_n48  &  wire717 ) ;
 assign wire16861 = ( (~ i_1_)  &  i_2_  &  (~ i_0_) ) ;
 assign wire16857 = ( n_n162  &  n_n163  &  n_n200 ) ;
 assign wire16863 = ( i_3_  &  n_n219 ) | ( n_n219  &  n_n111  &  n_n157 ) ;
 assign wire16865 = ( n_n7263 ) | ( n_n7264 ) | ( n_n135  &  wire16857 ) ;
 assign wire16867 = ( n_n3389 ) | ( n_n7252 ) | ( n_n7262 ) ;
 assign wire16871 = ( i_2_  &  (~ i_0_) ) | ( i_3_  &  (~ i_1_)  &  (~ i_2_)  &  i_0_ ) ;
 assign wire16884 = ( (~ i_7_)  &  i_6_  &  n_n218  &  n_n19 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n218  &  n_n19 ) ;
 assign wire16885 = ( i_3_  &  (~ i_1_)  &  i_2_  &  i_0_ ) | ( i_3_  &  (~ i_1_)  &  (~ i_2_)  &  i_0_ ) ;
 assign wire16888 = ( i_3_  &  (~ i_1_)  &  i_2_  &  i_0_ ) | ( i_3_  &  (~ i_1_)  &  (~ i_2_)  &  i_0_ ) ;
 assign wire16889 = ( n_n17  &  n_n219  &  n_n218 ) | ( n_n17  &  n_n219  &  n_n111 ) ;
 assign wire16890 = ( n_n162  &  n_n219  &  n_n18 ) | ( n_n219  &  n_n111  &  n_n18 ) ;
 assign wire16892 = ( n_n7263 ) | ( wire711 ) | ( n_n7264 ) ;
 assign wire16896 = ( wire388 ) | ( n_n2948 ) | ( wire16889 ) | ( wire16890 ) ;
 assign wire16910 = ( n_n5144 ) | ( wire729  &  n_n9  &  n_n156 ) ;
 assign wire16924 = ( n_n5144 ) | ( n_n39  &  n_n177  &  wire719 ) ;
 assign wire16929 = ( wire390 ) | ( wire393 ) | ( wire712 ) | ( wire16924 ) ;
 assign wire16930 = ( n_n969 ) | ( n_n519 ) | ( n_n4597 ) | ( wire4998 ) ;
 assign wire16936 = ( i_15_  &  n_n170  &  n_n215 ) | ( (~ i_15_)  &  n_n170  &  n_n215 ) ;
 assign wire16941 = ( n_n132  &  n_n33 ) | ( n_n34  &  wire78 ) ;
 assign wire16943 = ( wire443 ) | ( wire16941 ) | ( n_n31  &  wire143 ) ;
 assign wire16950 = ( _29458 ) | ( n_n34  &  wire150 ) | ( n_n34  &  wire16946 ) ;
 assign wire16957 = ( n_n36  &  wire147 ) | ( n_n36  &  wire125 ) ;
 assign wire16960 = ( wire607 ) | ( wire16957 ) | ( n_n36  &  wire149 ) ;
 assign wire16962 = ( n_n4169 ) | ( n_n4419 ) | ( wire4982 ) | ( wire16950 ) ;
 assign wire16966 = ( n_n30  &  wire131 ) | ( n_n31  &  wire125 ) ;
 assign wire16968 = ( wire4965 ) | ( wire4966 ) | ( wire655 ) | ( wire4961 ) ;
 assign wire16976 = ( n_n3510 ) | ( wire16968 ) | ( _29471 ) | ( _29472 ) ;
 assign wire16990 = ( n_n57  &  n_n125 ) | ( n_n108  &  n_n214 ) ;
 assign wire16991 = ( n_n5739 ) | ( n_n5743 ) | ( wire4948 ) | ( wire4950 ) ;
 assign wire16993 = ( wire4941 ) | ( wire16990 ) | ( wire16991 ) ;
 assign wire16994 = ( n_n4904 ) | ( wire4942 ) ;
 assign wire16995 = ( n_n101  &  wire86 ) | ( n_n108  &  wire250 ) ;
 assign wire16996 = ( wire4924 ) | ( n_n101  &  wire208 ) ;
 assign wire16997 = ( n_n5033 ) | ( wire4937 ) | ( wire16995 ) ;
 assign wire17001 = ( wire544 ) | ( wire16993 ) | ( wire16994 ) | ( wire16996 ) ;
 assign wire17003 = ( n_n41  &  n_n102 ) | ( n_n41  &  wire180 ) | ( n_n41  &  n_n202 ) ;
 assign wire17016 = ( n_n41  &  wire135 ) | ( n_n41  &  wire141 ) ;
 assign wire17028 = ( n_n34  &  wire168 ) | ( n_n34  &  wire74 ) ;
 assign wire17038 = ( n_n39  &  n_n132 ) | ( n_n38  &  n_n84 ) ;
 assign wire17039 = ( n_n38  &  n_n134 ) | ( n_n39  &  n_n134 ) | ( n_n38  &  n_n132 ) ;
 assign wire17041 = ( n_n4597 ) | ( wire17038 ) | ( wire17039 ) ;
 assign wire17042 = ( n_n40  &  n_n57 ) | ( n_n39  &  wire104 ) ;
 assign wire17044 = ( n_n38  &  wire279 ) | ( n_n39  &  wire279 ) ;
 assign wire17045 = ( n_n974 ) | ( wire17042 ) | ( n_n40  &  wire182 ) ;
 assign wire17047 = ( wire4869 ) | ( wire4863 ) | ( _29207 ) ;
 assign wire17053 = ( n_n47  &  n_n142 ) | ( n_n46  &  wire57 ) ;
 assign wire17055 = ( n_n5103 ) | ( wire652 ) | ( wire17053 ) ;
 assign wire17056 = ( wire4857 ) | ( wire4858 ) | ( wire4859 ) | ( wire4860 ) ;
 assign wire17058 = ( n_n6271 ) | ( n_n6270 ) | ( n_n57  &  n_n46 ) ;
 assign wire17060 = ( n_n6266 ) | ( n_n6268 ) | ( wire666 ) | ( wire17058 ) ;
 assign wire17061 = ( wire549 ) | ( wire4919 ) | ( wire17003 ) ;
 assign wire17063 = ( wire621 ) | ( wire17055 ) | ( wire17056 ) ;
 assign wire17067 = ( n_n108  &  n_n142 ) | ( n_n101  &  wire57 ) ;
 assign wire17071 = ( wire4832 ) | ( wire4838 ) | ( wire4839 ) | ( wire17067 ) ;
 assign wire17076 = ( wire445 ) | ( wire446 ) | ( wire4827 ) | ( wire4828 ) ;
 assign wire17079 = ( wire4820 ) | ( wire4821 ) | ( wire4822 ) | ( wire17076 ) ;
 assign wire17093 = ( n_n1606 ) | ( n_n46  &  wire142 ) | ( n_n46  &  wire180 ) ;
 assign wire17094 = ( wire4805 ) | ( n_n47  &  wire1170 ) ;
 assign wire17096 = ( wire4818 ) | ( wire4819 ) | ( wire17093 ) | ( wire17094 ) ;
 assign wire17106 = ( n_n125  &  n_n214 ) | ( n_n197  &  n_n63 ) ;
 assign wire17108 = ( wire422 ) | ( wire17106 ) | ( n_n197  &  wire125 ) ;
 assign wire17109 = ( _5628 ) | ( n_n212  &  wire796 ) ;
 assign wire17114 = ( _29315 ) | ( n_n125  &  wire108 ) | ( n_n125  &  wire258 ) ;
 assign wire17115 = ( n_n4674 ) | ( wire4780 ) | ( n_n123  &  wire1853 ) ;
 assign wire17116 = ( wire131  &  n_n197 ) | ( wire149  &  n_n212 ) ;
 assign wire17117 = ( n_n212  &  wire125 ) | ( n_n197  &  wire46 ) ;
 assign wire17119 = ( n_n4686 ) | ( wire704 ) | ( wire4786 ) | ( wire17117 ) ;
 assign wire17121 = ( wire17108 ) | ( wire17109 ) | ( wire17114 ) | ( wire17115 ) ;
 assign wire17122 = ( n_n125  &  wire135 ) | ( n_n125  &  wire141 ) ;
 assign wire17123 = ( wire142  &  n_n123 ) | ( n_n125  &  wire70 ) ;
 assign wire17125 = ( n_n123  &  n_n169 ) | ( n_n125  &  n_n176 ) ;
 assign wire17127 = ( n_n123  &  wire180 ) | ( n_n125  &  wire100 ) ;
 assign wire17128 = ( wire17125 ) | ( wire17127 ) | ( wire86  &  n_n123 ) ;
 assign wire17129 = ( wire394 ) | ( wire4765 ) | ( wire17123 ) ;
 assign wire17134 = ( n_n1708 ) | ( wire698 ) | ( wire4752 ) ;
 assign wire17136 = ( n_n125  &  wire182 ) | ( wire719  &  n_n216  &  n_n125 ) ;
 assign wire17137 = ( wire4768 ) | ( wire17122 ) | ( wire17136 ) ;
 assign wire17140 = ( wire4753 ) | ( wire17128 ) | ( wire17129 ) | ( wire17134 ) ;
 assign wire17141 = ( wire149  &  n_n197 ) | ( wire132  &  n_n212 ) ;
 assign wire17145 = ( wire17141 ) | ( wire132  &  n_n197 ) | ( n_n197  &  wire181 ) ;
 assign wire17146 = ( wire557 ) | ( wire648 ) | ( wire504 ) | ( wire578 ) ;
 assign wire17152 = ( n_n101  &  wire225 ) | ( n_n108  &  wire225 ) | ( n_n101  &  wire148 ) ;
 assign wire17153 = ( n_n5011 ) | ( wire591 ) | ( n_n101  &  wire250 ) ;
 assign wire17154 = ( wire4735 ) | ( wire17152 ) | ( n_n108  &  wire69 ) ;
 assign wire17156 = ( wire17071 ) | ( wire17079 ) | ( _29375 ) ;
 assign wire17158 = ( wire17001 ) | ( wire17096 ) | ( _29424 ) ;
 assign wire17166 = ( n_n5144 ) | ( n_n30  &  wire181 ) ;
 assign wire17170 = ( n_n4161 ) | ( wire695 ) | ( n_n30  &  wire132 ) ;
 assign wire17172 = ( wire599 ) | ( wire4993 ) | ( wire16943 ) ;
 assign wire17174 = ( wire16962 ) | ( wire16976 ) | ( _29474 ) ;
 assign wire17181 = ( n_n135  &  n_n101 ) | ( n_n135  &  n_n108 ) | ( n_n101  &  wire1179 ) ;
 assign wire17184 = ( n_n101  &  wire90 ) | ( n_n101  &  n_n61 ) | ( n_n108  &  n_n61 ) ;
 assign wire17185 = ( wire17181 ) | ( wire17184 ) | ( n_n108  &  wire1178 ) ;
 assign wire17187 = ( n_n51  &  n_n101 ) | ( n_n53  &  n_n101 ) | ( n_n51  &  n_n108 ) ;
 assign wire17191 = ( wire4684 ) | ( wire17187 ) | ( n_n47  &  wire181 ) ;
 assign wire17193 = ( n_n2253 ) | ( wire17185 ) | ( _5207 ) | ( _5208 ) ;
 assign wire17196 = ( n_n47  &  n_n61 ) | ( n_n46  &  n_n61 ) | ( n_n47  &  n_n63 ) ;
 assign wire17201 = ( n_n43  &  wire93 ) | ( wire729  &  n_n191  &  n_n43 ) ;
 assign wire17202 = ( wire725  &  n_n156  &  n_n47 ) | ( wire725  &  n_n156  &  n_n46 ) ;
 assign wire17203 = ( n_n57  &  n_n46 ) | ( n_n47  &  wire894 ) | ( n_n46  &  wire894 ) ;
 assign wire17206 = ( wire4669 ) | ( wire4676 ) | ( wire17201 ) | ( wire17202 ) ;
 assign wire17209 = ( n_n47  &  wire149 ) | ( n_n47  &  wire176 ) ;
 assign wire17212 = ( wire561 ) | ( wire4662 ) | ( wire4663 ) | ( wire17209 ) ;
 assign wire17220 = ( n_n33  &  wire60 ) | ( n_n32  &  n_n182 ) ;
 assign wire17226 = ( wire725  &  n_n156  &  n_n36 ) | ( wire725  &  n_n149  &  n_n36 ) ;
 assign wire17231 = ( n_n30  &  wire181 ) | ( n_n31  &  wire129 ) ;
 assign wire17239 = ( n_n31  &  wire158 ) | ( wire725  &  n_n31  &  n_n216 ) ;
 assign wire17241 = ( wire4638 ) | ( wire17239 ) | ( wire213  &  n_n61 ) ;
 assign wire17243 = ( n_n31  &  wire1189 ) | ( n_n31  &  wire1188 ) | ( n_n30  &  wire1188 ) ;
 assign wire17245 = ( n_n30  &  wire131 ) | ( n_n31  &  wire149 ) ;
 assign wire17246 = ( wire17243 ) | ( wire17245 ) | ( n_n30  &  wire1190 ) ;
 assign wire17247 = ( wire4628 ) | ( n_n31  &  wire902 ) ;
 assign wire17251 = ( n_n135  &  n_n125 ) | ( n_n135  &  n_n123 ) | ( n_n125  &  wire1177 ) ;
 assign wire17265 = ( n_n5739 ) | ( wire440 ) | ( n_n108  &  n_n210 ) ;
 assign wire17266 = ( wire447 ) | ( n_n5743 ) | ( n_n135  &  n_n113 ) ;
 assign wire17271 = ( i_15_  &  n_n211  &  n_n177 ) | ( (~ i_15_)  &  n_n211  &  n_n177 ) | ( i_15_  &  n_n211  &  n_n170 ) | ( (~ i_15_)  &  n_n211  &  n_n170 ) ;
 assign wire17275 = ( n_n77  &  n_n123 ) | ( wire117  &  n_n123 ) | ( n_n123  &  wire17271 ) ;
 assign wire17276 = ( wire4602 ) | ( n_n125  &  wire975 ) | ( n_n125  &  wire1234 ) ;
 assign wire17280 = ( n_n53  &  n_n40 ) | ( n_n38  &  n_n168 ) ;
 assign wire17281 = ( n_n51  &  wire190 ) | ( wire334  &  n_n78 ) ;
 assign wire17284 = ( n_n53  &  n_n41 ) | ( n_n41  &  wire1117 ) | ( n_n40  &  wire1117 ) ;
 assign wire17285 = ( n_n135  &  n_n41 ) | ( n_n135  &  n_n40 ) | ( n_n41  &  n_n57 ) | ( n_n40  &  n_n57 ) ;
 assign wire17288 = ( n_n39  &  wire1120 ) | ( n_n39  &  n_n156  &  wire726 ) ;
 assign wire17289 = ( wire4581 ) | ( wire17284 ) | ( wire17285 ) ;
 assign wire17290 = ( wire4591 ) | ( wire17280 ) | ( wire17281 ) | ( wire17288 ) ;
 assign wire17291 = ( n_n71  &  n_n41 ) | ( n_n41  &  n_n150 ) | ( n_n41  &  wire377 ) ;
 assign wire17297 = ( wire4572 ) | ( wire725  &  n_n199  &  wire190 ) ;
 assign wire17298 = ( wire4573 ) | ( wire4576 ) | ( wire17291 ) ;
 assign wire17299 = ( n_n36  &  n_n102 ) | ( n_n38  &  n_n150 ) ;
 assign wire17301 = ( n_n34  &  n_n102 ) | ( n_n36  &  wire978 ) ;
 assign wire17309 = ( i_15_  &  n_n211  &  n_n149 ) | ( (~ i_15_)  &  n_n211  &  n_n149 ) | ( (~ i_15_)  &  n_n149  &  n_n201 ) ;
 assign wire17325 = ( wire4550 ) | ( wire4551 ) | ( _29890 ) ;
 assign wire17337 = ( n_n41  &  wire69 ) | ( n_n156  &  wire722  &  n_n41 ) ;
 assign wire17338 = ( n_n40  &  n_n102 ) | ( n_n40  &  n_n202 ) | ( n_n40  &  wire263 ) ;
 assign wire17359 = ( wire4500 ) | ( n_n101  &  wire1060 ) ;
 assign wire17360 = ( n_n101  &  wire86 ) | ( n_n101  &  wire263 ) ;
 assign wire17363 = ( wire4491 ) | ( wire4496 ) | ( wire17360 ) ;
 assign wire17364 = ( wire17363 ) | ( n_n108  &  wire1064 ) ;
 assign wire17365 = ( n_n2257 ) | ( wire4504 ) | ( wire17359 ) | ( _29963 ) ;
 assign wire17377 = ( n_n212  &  wire168 ) | ( n_n197  &  wire181 ) | ( n_n212  &  wire181 ) ;
 assign wire17382 = ( n_n51  &  n_n197 ) | ( n_n53  &  n_n197 ) | ( n_n51  &  n_n212 ) | ( n_n53  &  n_n212 ) ;
 assign wire17383 = ( n_n197  &  wire176 ) | ( n_n212  &  n_n63 ) ;
 assign wire17384 = ( n_n197  &  n_n61 ) | ( n_n212  &  n_n61 ) | ( n_n197  &  wire308 ) ;
 assign wire17388 = ( n_n197  &  n_n55 ) | ( n_n212  &  n_n55 ) | ( n_n197  &  wire887 ) ;
 assign wire17389 = ( _30001 ) | ( n_n212  &  wire299 ) | ( n_n212  &  wire17385 ) ;
 assign wire17390 = ( wire17383 ) | ( wire17384 ) | ( wire17388 ) ;
 assign wire17392 = ( n_n117  &  n_n125 ) | ( n_n102  &  n_n123 ) ;
 assign wire17393 = ( wire4458 ) | ( wire4459 ) | ( wire17392 ) ;
 assign wire17394 = ( wire4453 ) | ( wire4454 ) ;
 assign wire17397 = ( n_n102  &  n_n125 ) | ( n_n125  &  wire243 ) | ( n_n125  &  wire17395 ) ;
 assign wire17398 = ( wire4470 ) | ( wire17382 ) | ( n_n123  &  wire1124 ) ;
 assign wire17400 = ( wire17389 ) | ( wire17390 ) | ( wire17393 ) | ( wire17394 ) ;
 assign wire17405 = ( n_n2234 ) | ( wire17397 ) | ( wire17398 ) | ( wire17400 ) ;
 assign wire17417 = ( n_n33  &  wire60 ) | ( wire719  &  n_n149  &  n_n33 ) ;
 assign wire17418 = ( n_n31  &  wire143 ) | ( n_n34  &  wire122 ) ;
 assign wire17433 = ( wire4419 ) | ( wire4427 ) | ( n_n30  &  wire144 ) ;
 assign wire17434 = ( n_n4154 ) | ( wire654 ) | ( _4479 ) | ( _30218 ) ;
 assign wire17435 = ( wire17433 ) | ( _4473 ) | ( _30224 ) | ( _30229 ) ;
 assign wire17436 = ( n_n34  &  wire133 ) | ( n_n34  &  wire181 ) ;
 assign wire17439 = ( wire458 ) | ( wire17436 ) | ( n_n34  &  wire127 ) ;
 assign wire17440 = ( n_n34  &  wire134 ) | ( n_n34  &  wire123 ) ;
 assign wire17441 = ( n_n34  &  wire156 ) | ( n_n34  &  wire176 ) ;
 assign wire17443 = ( n_n36  &  wire55 ) | ( n_n36  &  wire127 ) ;
 assign wire17446 = ( wire17440 ) | ( wire17443 ) | ( n_n36  &  wire158 ) ;
 assign wire17450 = ( n_n34  &  wire125 ) | ( wire725  &  n_n34  &  n_n216 ) ;
 assign wire17452 = ( n_n4564 ) | ( wire709 ) | ( wire4396 ) | ( wire4986 ) ;
 assign wire17453 = ( wire4395 ) | ( wire17450 ) | ( wire17452 ) ;
 assign wire17454 = ( wire17439 ) | ( wire17446 ) | ( _30244 ) ;
 assign wire17456 = ( wire4768 ) | ( wire17122 ) | ( wire157  &  n_n125 ) ;
 assign wire17457 = ( wire4393 ) | ( wire4750 ) | ( _30176 ) ;
 assign wire17458 = ( wire86  &  n_n123 ) | ( wire720  &  n_n149  &  n_n123 ) ;
 assign wire17459 = ( n_n125  &  wire155 ) | ( n_n123  &  wire180 ) ;
 assign wire17462 = ( wire570 ) | ( wire4765 ) | ( wire17123 ) | ( wire17458 ) ;
 assign wire17465 = ( n_n1700 ) | ( n_n125  &  wire803 ) ;
 assign wire17467 = ( wire17456 ) | ( wire17457 ) | ( wire17465 ) ;
 assign wire17469 = ( n_n101  &  wire90 ) | ( n_n108  &  n_n142 ) ;
 assign wire17484 = ( n_n6005 ) | ( wire419 ) | ( n_n1624 ) | ( wire4344 ) ;
 assign wire17493 = ( n_n46  &  wire142 ) | ( n_n46  &  wire799 ) | ( n_n46  &  wire180 ) ;
 assign wire17499 = ( n_n1594 ) | ( n_n47  &  wire808 ) ;
 assign wire17504 = ( n_n5000 ) | ( n_n101  &  wire86 ) | ( n_n101  &  wire84 ) ;
 assign wire17505 = ( n_n4900 ) | ( n_n108  &  wire867 ) ;
 assign wire17507 = ( n_n5739 ) | ( wire4950 ) | ( n_n53  &  n_n123 ) ;
 assign wire17509 = ( n_n5037 ) | ( wire17507 ) | ( wire157  &  n_n123 ) ;
 assign wire17513 = ( n_n4903 ) | ( wire17504 ) | ( wire17505 ) | ( wire17509 ) ;
 assign wire17516 = ( wire55  &  n_n212 ) | ( n_n197  &  wire181 ) ;
 assign wire17518 = ( wire127  &  n_n197 ) | ( n_n212  &  wire123 ) ;
 assign wire17537 = ( wire4285 ) | ( wire4908 ) | ( wire17016 ) ;
 assign wire17541 = ( n_n38  &  n_n156  &  wire728 ) | ( n_n38  &  n_n156  &  wire726 ) ;
 assign wire17542 = ( n_n39  &  n_n54 ) | ( n_n38  &  n_n52 ) | ( n_n39  &  n_n52 ) ;
 assign wire17543 = ( n_n1514 ) | ( wire17541 ) | ( wire17542 ) ;
 assign wire17545 = ( n_n38  &  wire248 ) | ( n_n39  &  wire248 ) ;
 assign wire17548 = ( n_n1520 ) | ( wire571 ) | ( n_n39  &  wire110 ) ;
 assign wire17549 = ( n_n1517 ) | ( wire17545 ) | ( n_n39  &  wire249 ) ;
 assign wire17550 = ( wire457 ) | ( wire4263 ) | ( wire4888 ) | ( wire17028 ) ;
 assign wire17555 = ( n_n46  &  wire90 ) | ( n_n47  &  n_n142 ) ;
 assign wire17557 = ( wire4260 ) | ( wire17554 ) | ( wire652 ) ;
 assign wire17558 = ( n_n4312 ) | ( wire4859 ) | ( wire4860 ) | ( wire17555 ) ;
 assign wire17559 = ( wire4252 ) | ( wire4253 ) | ( n_n53  &  n_n46 ) ;
 assign wire17560 = ( n_n6267 ) | ( n_n6269 ) | ( wire157  &  n_n46 ) ;
 assign wire17562 = ( wire17559 ) | ( wire17560 ) | ( n_n47  &  wire152 ) ;
 assign wire17565 = ( wire621 ) | ( wire17557 ) | ( wire17558 ) ;
 assign wire17568 = ( wire122  &  n_n197 ) | ( n_n125  &  n_n214 ) ;
 assign wire17574 = ( wire422 ) | ( wire4234 ) | ( wire17568 ) ;
 assign wire17575 = ( n_n197  &  wire176 ) | ( n_n212  &  wire125 ) ;
 assign wire17578 = ( n_n4231 ) | ( wire565 ) | ( _4527 ) | ( _30195 ) ;
 assign wire17579 = ( wire17115 ) | ( wire17574 ) | ( _30203 ) ;
 assign wire17581 = ( n_n4116 ) | ( wire17578 ) | ( wire17579 ) ;
 assign wire17585 = ( wire17434 ) | ( wire17435 ) | ( wire17453 ) | ( wire17454 ) ;
 assign wire17592 = ( wire4220 ) | ( wire170  &  wire1527 ) ;
 assign wire17593 = ( n_n5  &  n_n144 ) | ( n_n9  &  n_n144 ) | ( n_n6  &  n_n144 ) ;
 assign wire17594 = ( n_n162  &  n_n219  &  n_n157 ) | ( n_n219  &  n_n48  &  n_n157 ) ;
 assign wire17596 = ( n_n16  &  n_n219  &  n_n218 ) | ( n_n16  &  n_n219  &  n_n48 ) ;
 assign wire17599 = ( wire569 ) | ( wire17594 ) | ( n_n14  &  wire170 ) ;
 assign wire17605 = ( n_n5144 ) | ( n_n19  &  n_n111  &  n_n157 ) ;
 assign wire17606 = ( i_7_  &  i_6_  &  n_n19  &  n_n111 ) | ( (~ i_7_)  &  i_6_  &  n_n19  &  n_n111 ) | ( i_7_  &  (~ i_6_)  &  n_n19  &  n_n111 ) ;
 assign wire17608 = ( wire569 ) | ( wire725  &  n_n13  &  n_n149 ) ;
 assign wire17610 = ( wire529 ) | ( wire568 ) | ( n_n4  &  wire77 ) ;
 assign wire17622 = ( wire445 ) | ( n_n53  &  n_n108 ) | ( wire157  &  n_n108 ) ;
 assign wire17626 = ( n_n4981 ) | ( wire4172 ) ;
 assign wire17627 = ( wire17622 ) | ( n_n101  &  wire1321 ) | ( n_n101  &  wire1488 ) ;
 assign wire17629 = ( n_n3823 ) | ( _30484 ) ;
 assign wire17631 = ( n_n134  &  n_n46 ) | ( n_n47  &  wire78 ) ;
 assign wire17635 = ( n_n6266 ) | ( wire725  &  n_n156  &  n_n47 ) ;
 assign wire17638 = ( wire4159 ) | ( n_n47  &  wire172 ) | ( n_n47  &  wire80 ) ;
 assign wire17639 = ( n_n6271 ) | ( n_n6267 ) | ( wire17635 ) | ( wire17638 ) ;
 assign wire17640 = ( wire651 ) | ( wire4158 ) | ( wire17631 ) ;
 assign wire17646 = ( n_n1553 ) | ( wire500 ) | ( wire361 ) | ( wire4151 ) ;
 assign wire17647 = ( wire497 ) | ( n_n40  &  wire1450 ) ;
 assign wire17650 = ( n_n3542 ) | ( n_n41  &  wire215 ) | ( n_n41  &  n_n155 ) ;
 assign wire17651 = ( wire397 ) | ( wire653 ) | ( wire4143 ) ;
 assign wire17654 = ( n_n41  &  n_n214 ) | ( n_n40  &  n_n214 ) | ( n_n40  &  wire180 ) ;
 assign wire17656 = ( wire359 ) | ( wire537 ) | ( n_n43  &  n_n59 ) ;
 assign wire17659 = ( wire17654 ) | ( wire17656 ) | ( _30358 ) | ( _30359 ) ;
 assign wire17660 = ( wire17646 ) | ( wire17647 ) | ( wire17650 ) | ( wire17651 ) ;
 assign wire17662 = ( n_n41  &  n_n57 ) | ( n_n41  &  wire182 ) | ( n_n41  &  n_n130 ) ;
 assign wire17663 = ( n_n38  &  wire104 ) | ( n_n38  &  wire279 ) ;
 assign wire17667 = ( n_n38  &  n_n134 ) | ( n_n39  &  n_n134 ) | ( n_n38  &  wire110 ) ;
 assign wire17668 = ( n_n38  &  n_n54 ) | ( n_n39  &  n_n54 ) | ( n_n38  &  n_n150 ) | ( n_n39  &  n_n150 ) ;
 assign wire17672 = ( wire605 ) | ( n_n972 ) | ( wire17663 ) | ( wire17667 ) ;
 assign wire17674 = ( n_n71  &  n_n41 ) | ( n_n41  &  n_n150 ) | ( n_n41  &  wire141 ) ;
 assign wire17677 = ( n_n3979 ) | ( wire442 ) | ( wire4113 ) ;
 assign wire17679 = ( n_n40  &  _30386 ) | ( wire725  &  n_n40  &  _29298 ) ;
 assign wire17681 = ( wire17679 ) | ( _4253 ) | ( wire104  &  _30385 ) ;
 assign wire17684 = ( wire4104 ) | ( wire17681 ) | ( _30390 ) | ( _30391 ) ;
 assign wire17685 = ( wire17672 ) | ( wire17677 ) | ( _30404 ) ;
 assign wire17686 = ( n_n47  &  n_n63 ) | ( n_n46  &  wire212 ) ;
 assign wire17688 = ( n_n46  &  wire134 ) | ( n_n47  &  wire125 ) ;
 assign wire17690 = ( n_n5107 ) | ( wire688 ) | ( n_n46  &  wire176 ) ;
 assign wire17691 = ( wire560 ) | ( wire17686 ) | ( wire17688 ) ;
 assign wire17692 = ( n_n43  &  wire52 ) | ( n_n43  &  wire129 ) ;
 assign wire17693 = ( n_n42  &  wire63 ) | ( n_n43  &  wire63 ) | ( n_n42  &  wire48 ) | ( n_n43  &  wire48 ) ;
 assign wire17695 = ( wire4102 ) | ( wire4103 ) | ( wire17692 ) | ( wire17693 ) ;
 assign wire17696 = ( wire17639 ) | ( wire17640 ) | ( wire17690 ) | ( wire17691 ) ;
 assign wire17698 = ( wire17659 ) | ( wire17660 ) | ( wire17684 ) | ( wire17685 ) ;
 assign wire17700 = ( wire419 ) | ( n_n200  &  wire1375 ) ;
 assign wire17701 = ( wire47  &  n_n46 ) | ( n_n46  &  wire181 ) ;
 assign wire17704 = ( wire481 ) | ( wire17700 ) | ( wire17701 ) ;
 assign wire17705 = ( wire131  &  n_n46 ) | ( n_n47  &  wire129 ) ;
 assign wire17706 = ( wire137  &  n_n46 ) | ( wire146  &  n_n46 ) | ( n_n46  &  wire46 ) ;
 assign wire17708 = ( wire4088 ) | ( wire17705 ) | ( n_n47  &  wire46 ) ;
 assign wire17709 = ( n_n3889 ) | ( n_n3561 ) ;
 assign wire17710 = ( wire674 ) | ( wire671 ) | ( wire17706 ) ;
 assign wire17712 = ( wire577 ) | ( wire4080 ) | ( wire17704 ) | ( wire17710 ) ;
 assign wire17721 = ( wire729  &  n_n191 ) | ( wire720  &  n_n191 ) | ( wire715  &  n_n191 ) ;
 assign wire17725 = ( wire157  &  n_n123 ) | ( wire725  &  n_n156  &  n_n123 ) ;
 assign wire17732 = ( n_n125  &  wire141 ) | ( n_n125  &  wire160 ) ;
 assign wire17735 = ( n_n2859 ) | ( n_n4657 ) | ( wire4048 ) | ( wire17732 ) ;
 assign wire17740 = ( wire479 ) | ( wire90  &  n_n125 ) | ( n_n125  &  wire205 ) ;
 assign wire17744 = ( n_n125  &  n_n176 ) | ( n_n125  &  wire51 ) | ( n_n123  &  wire51 ) ;
 assign wire17746 = ( wire394 ) | ( n_n123  &  wire1420 ) ;
 assign wire17748 = ( n_n3912 ) | ( wire4043 ) | ( wire17735 ) | ( wire17740 ) ;
 assign wire17750 = ( n_n134  &  n_n197 ) | ( n_n53  &  n_n212 ) ;
 assign wire17753 = ( wire422 ) | ( wire4026 ) | ( wire17568 ) | ( wire17750 ) ;
 assign wire17757 = ( wire565 ) | ( wire4021 ) | ( wire4230 ) | ( wire17575 ) ;
 assign wire17760 = ( wire86  &  n_n123 ) | ( n_n123  &  wire180 ) ;
 assign wire17761 = ( wire85  &  n_n123 ) | ( wire142  &  n_n123 ) | ( n_n123  &  n_n214 ) ;
 assign wire17764 = ( n_n3592 ) | ( wire4013 ) | ( wire17760 ) | ( wire17761 ) ;
 assign wire17765 = ( wire17753 ) | ( wire17757 ) | ( _30453 ) ;
 assign wire17772 = ( n_n212  &  wire48 ) | ( n_n197  &  wire181 ) ;
 assign wire17773 = ( wire47  &  n_n197 ) | ( n_n212  &  wire181 ) ;
 assign wire17776 = ( n_n4518 ) | ( wire3998 ) | ( wire17772 ) | ( wire17773 ) ;
 assign wire17778 = ( n_n3834 ) | ( n_n3833 ) | ( wire17776 ) ;
 assign wire17779 = ( wire17748 ) | ( wire17765 ) | ( _30455 ) ;
 assign wire17783 = ( n_n31  &  wire125 ) | ( wire725  &  n_n31  &  n_n216 ) ;
 assign wire17786 = ( wire3991 ) | ( wire3996 ) | ( _30491 ) ;
 assign wire17796 = ( n_n30  &  wire137 ) | ( n_n31  &  wire46 ) | ( n_n30  &  wire46 ) ;
 assign wire17800 = ( n_n36  &  _30549 ) | ( wire725  &  n_n36  &  _29298 ) ;
 assign wire17801 = ( n_n34  &  wire134 ) | ( n_n34  &  wire123 ) ;
 assign wire17806 = ( wire541 ) | ( n_n4566 ) | ( wire3964 ) | ( wire17800 ) ;
 assign wire17810 = ( n_n53  &  n_n36 ) | ( n_n134  &  n_n34 ) ;
 assign wire17813 = ( wire636 ) | ( wire3958 ) | ( wire17810 ) ;
 assign wire17816 = ( n_n31  &  wire143 ) | ( n_n33  &  n_n138 ) ;
 assign wire17817 = ( n_n30  &  wire47 ) | ( n_n31  &  wire181 ) ;
 assign wire17818 = ( wire17816 ) | ( n_n31  &  wire154 ) | ( n_n31  &  wire47 ) ;
 assign wire17819 = ( wire17817 ) | ( n_n33  &  wire1519 ) ;
 assign wire17821 = ( wire17806 ) | ( wire17813 ) | ( _30557 ) ;
 assign wire17822 = ( n_n34  &  wire52 ) | ( n_n36  &  wire46 ) ;
 assign wire17824 = ( n_n38  &  n_n134 ) | ( n_n38  &  n_n54 ) | ( n_n39  &  n_n54 ) ;
 assign wire17825 = ( wire143  &  n_n34 ) | ( n_n34  &  wire181 ) ;
 assign wire17826 = ( wire143  &  n_n36 ) | ( wire154  &  n_n34 ) ;
 assign wire17827 = ( wire47  &  n_n34 ) | ( n_n36  &  wire181 ) ;
 assign wire17830 = ( wire432 ) | ( wire17824 ) | ( wire17827 ) ;
 assign wire17837 = ( wire458 ) | ( wire640 ) | ( wire642 ) | ( wire606 ) ;
 assign wire17840 = ( n_n5144 ) | ( wire725  &  n_n156  &  wire213 ) ;
 assign wire17844 = ( n_n3795 ) | ( wire17708 ) | ( wire17709 ) | ( wire17712 ) ;
 assign wire17845 = ( n_n3787 ) | ( wire17818 ) | ( wire17819 ) | ( wire17821 ) ;
 assign wire17850 = ( n_n162  &  n_n17  &  n_n219 ) | ( n_n17  &  n_n219  &  n_n218 ) ;
 assign wire17852 = ( wire463 ) | ( wire17850 ) ;
 assign wire17853 = ( wire568 ) | ( n_n7264 ) | ( n_n14  &  wire145 ) ;
 assign wire17854 = ( wire3899 ) | ( wire145  &  wire1044 ) ;
 assign wire17858 = ( n_n7252 ) | ( n_n7242 ) | ( wire3887 ) ;
 assign wire17864 = ( n_n34  &  wire127 ) | ( n_n36  &  wire123 ) ;
 assign wire17865 = ( wire137  &  n_n34 ) | ( n_n36  &  wire176 ) ;
 assign wire17868 = ( wire458 ) | ( wire17865 ) | ( n_n34  &  wire55 ) ;
 assign wire17870 = ( n_n3525 ) | ( wire17822 ) | ( n_n34  &  wire129 ) ;
 assign wire17872 = ( n_n36  &  wire147 ) | ( n_n34  &  wire147 ) ;
 assign wire17873 = ( n_n36  &  wire149 ) | ( n_n34  &  wire126 ) ;
 assign wire17887 = ( n_n134  &  n_n34 ) | ( n_n36  &  wire186 ) ;
 assign wire17889 = ( n_n34  &  wire176 ) | ( wire725  &  n_n34  &  n_n216 ) ;
 assign wire17891 = ( n_n36  &  wire125 ) | ( n_n34  &  wire125 ) ;
 assign wire17893 = ( n_n4564 ) | ( wire709 ) | ( wire17889 ) ;
 assign wire17894 = ( wire3850 ) | ( wire3851 ) | ( wire17891 ) ;
 assign wire17906 = ( wire636 ) | ( wire3835 ) | ( wire17887 ) ;
 assign wire17908 = ( n_n2626 ) | ( wire17893 ) | ( wire17894 ) ;
 assign wire17911 = ( n_n5144 ) | ( wire725  &  n_n156  &  n_n36 ) ;
 assign wire17916 = ( wire725  &  n_n156 ) | ( wire719  &  n_n149 ) ;
 assign wire17931 = ( n_n31  &  wire129 ) | ( n_n31  &  wire46 ) ;
 assign wire17955 = ( n_n39  &  n_n132 ) | ( n_n39  &  n_n54 ) | ( n_n39  &  n_n52 ) ;
 assign wire17963 = ( n_n36  &  wire52 ) | ( n_n36  &  wire129 ) ;
 assign wire17964 = ( n_n36  &  wire139 ) | ( n_n36  &  wire46 ) ;
 assign wire17965 = ( n_n36  &  wire130 ) | ( n_n36  &  wire124 ) | ( n_n36  &  wire128 ) ;
 assign wire17976 = ( n_n6267 ) | ( n_n6266 ) | ( n_n6270 ) | ( wire3774 ) ;
 assign wire17985 = ( n_n41  &  wire85 ) | ( n_n41  &  n_n214 ) | ( n_n41  &  n_n198 ) ;
 assign wire17987 = ( wire17985 ) | ( n_n41  &  wire142 ) | ( n_n41  &  wire180 ) ;
 assign wire17988 = ( wire524 ) | ( wire359 ) | ( n_n4476 ) | ( wire3759 ) ;
 assign wire17989 = ( i_9_  &  (~ i_10_)  &  i_11_  &  wire720 ) | ( (~ i_9_)  &  (~ i_10_)  &  (~ i_11_)  &  wire720 ) ;
 assign wire17995 = ( wire497 ) | ( n_n41  &  wire51 ) | ( n_n41  &  wire70 ) ;
 assign wire17996 = ( n_n41  &  n_n83 ) | ( n_n41  &  wire69 ) | ( n_n41  &  n_n171 ) ;
 assign wire17999 = ( wire694 ) | ( n_n3542 ) | ( wire17996 ) ;
 assign wire18000 = ( wire426 ) | ( wire3747 ) | ( wire17999 ) ;
 assign wire18001 = ( wire3755 ) | ( wire17987 ) | ( wire17988 ) | ( wire17995 ) ;
 assign wire18003 = ( n_n39  &  wire207 ) | ( n_n39  &  wire248 ) | ( n_n39  &  n_n78 ) ;
 assign wire18010 = ( n_n41  &  n_n57 ) | ( n_n39  &  wire104 ) ;
 assign wire18012 = ( wire18010 ) | ( wire245  &  n_n41 ) | ( n_n41  &  wire182 ) ;
 assign wire18013 = ( n_n41  &  wire1807 ) | ( n_n41  &  wire1811 ) ;
 assign wire18017 = ( n_n71  &  n_n41 ) | ( n_n41  &  n_n150 ) | ( n_n41  &  wire141 ) ;
 assign wire18018 = ( _30710 ) | ( n_n41  &  wire155 ) | ( n_n41  &  wire205 ) ;
 assign wire18019 = ( wire18017 ) | ( n_n41  &  wire1812 ) ;
 assign wire18021 = ( n_n39  &  n_n177  &  wire719 ) | ( n_n39  &  wire719  &  n_n170 ) ;
 assign wire18023 = ( wire434 ) | ( wire18021 ) | ( n_n39  &  wire249 ) ;
 assign wire18026 = ( wire3723 ) | ( wire18023 ) | ( _30702 ) | ( _30703 ) ;
 assign wire18027 = ( wire18012 ) | ( wire18013 ) | ( wire18018 ) | ( wire18019 ) ;
 assign wire18035 = ( n_n47  &  wire129 ) | ( n_n47  &  wire130 ) ;
 assign wire18036 = ( n_n47  &  wire124 ) | ( n_n47  &  wire46 ) ;
 assign wire18071 = ( wire445 ) | ( wire157  &  n_n108 ) ;
 assign wire18074 = ( wire131 ) | ( wire126 ) ;
 assign wire18075 = ( wire132 ) | ( wire149 ) | ( wire147 ) | ( wire134 ) ;
 assign wire18076 = ( n_n108  &  wire1489 ) | ( n_n108  &  wire18074 ) | ( n_n108  &  wire18075 ) ;
 assign wire18085 = ( n_n125  &  wire85 ) | ( n_n125  &  wire142 ) | ( n_n125  &  n_n214 ) ;
 assign wire18089 = ( wire55  &  n_n212 ) | ( wire158  &  n_n212 ) ;
 assign wire18096 = ( n_n3592 ) | ( wire538 ) | ( wire539 ) | ( wire3665 ) ;
 assign wire18097 = ( wire3671 ) | ( wire3676 ) | ( _30799 ) ;
 assign wire18098 = ( wire725  &  n_n199 ) | ( wire719  &  n_n216 ) ;
 assign wire18106 = ( n_n125  &  wire182 ) | ( n_n125  &  wire141 ) ;
 assign wire18107 = ( (~ i_9_)  &  (~ i_10_)  &  i_11_  &  wire720 ) | ( (~ i_9_)  &  (~ i_10_)  &  (~ i_11_)  &  wire720 ) ;
 assign wire18120 = ( wire394 ) | ( wire3662 ) | ( _30816 ) | ( _30817 ) ;
 assign wire18128 = ( n_n212  &  wire168 ) | ( n_n212  &  wire151 ) ;
 assign wire18129 = ( n_n212  &  wire48 ) | ( n_n212  &  wire181 ) ;
 assign wire18132 = ( n_n4518 ) | ( wire3643 ) | ( wire18128 ) | ( wire18129 ) ;
 assign wire18134 = ( n_n3501 ) | ( n_n3500 ) | ( wire18132 ) ;
 assign wire18136 = ( n_n47  &  wire55 ) | ( n_n47  &  wire125 ) ;
 assign wire18145 = ( _30839 ) | ( n_n31  &  wire1601 ) ;
 assign wire18158 = ( n_n5144 ) | ( n_n219  &  n_n48  &  n_n157 ) ;
 assign wire18159 = ( i_7_  &  (~ i_6_)  &  n_n219  &  n_n111 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n219  &  n_n111 ) ;
 assign wire18160 = ( n_n17  &  n_n219  &  n_n218 ) | ( n_n17  &  n_n219  &  n_n48 ) ;
 assign wire18161 = ( n_n162  &  n_n219  &  n_n157 ) | ( n_n219  &  n_n218  &  n_n157 ) ;
 assign wire18163 = ( wire18160 ) | ( wire18161 ) ;
 assign wire18164 = ( wire18158 ) | ( wire18159 ) | ( n_n14  &  wire253 ) ;
 assign wire18178 = ( n_n47  &  wire129 ) | ( n_n47  &  wire124 ) ;
 assign wire18182 = ( wire131  &  n_n46 ) | ( n_n47  &  wire176 ) ;
 assign wire18185 = ( wire546 ) | ( wire18182 ) | ( n_n47  &  wire123 ) ;
 assign wire18187 = ( n_n3889 ) | ( wire4088 ) | ( n_n47  &  wire46 ) ;
 assign wire18190 = ( n_n46  &  wire176 ) | ( n_n47  &  n_n63 ) ;
 assign wire18191 = ( n_n47  &  n_n140 ) | ( n_n47  &  wire247 ) | ( n_n47  &  wire125 ) ;
 assign wire18193 = ( wire3580 ) | ( wire3581 ) | ( wire18191 ) ;
 assign wire18196 = ( n_n184  &  wire725 ) | ( n_n177  &  wire719 ) ;
 assign wire18201 = ( wire3570 ) | ( _3429 ) | ( _3430 ) ;
 assign wire18202 = ( n_n47  &  wire55 ) | ( n_n46  &  wire134 ) ;
 assign wire18205 = ( wire688 ) | ( n_n3555 ) | ( wire3563 ) | ( wire18202 ) ;
 assign wire18209 = ( n_n47  &  wire149 ) | ( n_n46  &  wire46 ) ;
 assign wire18210 = ( wire132  &  n_n47 ) | ( n_n47  &  wire126 ) | ( n_n47  &  wire147 ) ;
 assign wire18220 = ( n_n5144 ) | ( n_n6271 ) | ( wire4252 ) | ( wire4253 ) ;
 assign wire18221 = ( n_n6267 ) | ( n_n6266 ) | ( n_n6270 ) | ( n_n6269 ) ;
 assign wire18222 = ( n_n6268 ) | ( n_n53  &  n_n46 ) | ( wire157  &  n_n46 ) ;
 assign wire18232 = ( n_n6384 ) | ( n_n3419 ) | ( n_n41  &  wire1036 ) ;
 assign wire18234 = ( n_n53  &  n_n46 ) | ( n_n41  &  n_n202 ) ;
 assign wire18237 = ( n_n4308 ) | ( n_n3421 ) | ( wire391 ) | ( wire18234 ) ;
 assign wire18238 = ( wire4260 ) | ( wire17554 ) | ( wire3533 ) | ( wire3607 ) ;
 assign wire18243 = ( wire3526 ) | ( wire3531 ) | ( n_n40  &  n_n95 ) ;
 assign wire18245 = ( wire18237 ) | ( wire18238 ) | ( wire18243 ) ;
 assign wire18252 = ( n_n3417 ) | ( n_n41  &  wire1174 ) ;
 assign wire18264 = ( n_n41  &  n_n83 ) | ( n_n41  &  n_n171 ) | ( n_n41  &  wire469 ) ;
 assign wire18266 = ( n_n3415 ) | ( wire18264 ) | ( n_n40  &  wire1331 ) ;
 assign wire18268 = ( wire3515 ) | ( wire3516 ) | ( wire3520 ) | ( wire18252 ) ;
 assign wire18269 = ( n_n40  &  _30964 ) | ( wire719  &  n_n40  &  _30347 ) ;
 assign wire18270 = ( n_n40  &  wire172 ) | ( n_n41  &  wire182 ) ;
 assign wire18278 = ( n_n156  &  wire717 ) | ( n_n156  &  wire724 ) ;
 assign wire18287 = ( wire673 ) | ( wire3479 ) | ( _30984 ) ;
 assign wire18290 = ( wire18237 ) | ( wire18238 ) | ( wire18243 ) | ( _31044 ) ;
 assign wire18294 = ( wire3550 ) | ( _3273 ) | ( n_n41  &  _31050 ) ;
 assign wire18295 = ( n_n5052 ) | ( n_n5055 ) | ( n_n5058 ) | ( wire4900 ) ;
 assign wire18300 = ( n_n33  &  _31081 ) | ( wire719  &  n_n33  &  _29117 ) ;
 assign wire18307 = ( n_n5144 ) | ( wire719  &  n_n33  &  n_n191 ) ;
 assign wire18318 = ( (~ i_7_)  &  i_6_  &  n_n19  &  n_n111 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n19  &  n_n111 ) ;
 assign wire18321 = ( wire431 ) | ( wire529 ) | ( wire18318 ) ;
 assign wire18324 = ( n_n5144 ) | ( n_n219  &  n_n111  &  n_n157 ) ;
 assign wire18325 = ( wire18324 ) | ( n_n9  &  wire717  &  n_n149 ) ;
 assign wire18328 = ( n_n3389 ) | ( wire388 ) | ( n_n9  &  wire770 ) ;
 assign wire18334 = ( n_n184  &  wire725 ) | ( n_n184  &  wire719 ) | ( n_n184  &  wire728 ) ;
 assign wire18348 = ( wire526 ) | ( wire3397 ) | ( n_n42  &  n_n138 ) ;
 assign wire18353 = ( n_n1575 ) | ( wire3392 ) | ( n_n42  &  wire1782 ) ;
 assign wire18358 = ( n_n41  &  wire182 ) | ( n_n40  &  wire182 ) ;
 assign wire18370 = ( n_n7263 ) | ( n_n5319 ) | ( n_n7264 ) ;
 assign wire18371 = ( n_n7242 ) | ( wire463 ) | ( n_n7262 ) ;
 assign wire18372 = ( wire428 ) | ( n_n3276 ) | ( _31151 ) ;
 assign wire18388 = ( wire729  &  n_n156 ) | ( wire719  &  n_n199 ) ;
 assign wire18393 = ( n_n5107 ) | ( wire3342 ) | ( n_n47  &  wire172 ) ;
 assign wire18397 = ( n_n5103 ) | ( wire666 ) | ( wire3337 ) ;
 assign wire18398 = ( wire3338 ) | ( wire4857 ) | ( n_n46  &  wire209 ) ;
 assign wire18401 = ( n_n5109 ) | ( n_n47  &  wire1326 ) ;
 assign wire18403 = ( wire18397 ) | ( wire18398 ) | ( wire18401 ) ;
 assign wire18409 = ( wire498 ) | ( n_n46  &  wire951 ) ;
 assign wire18411 = ( n_n5319 ) | ( n_n46  &  wire168 ) ;
 assign wire18414 = ( wire481 ) | ( wire18411 ) | ( n_n46  &  wire151 ) ;
 assign wire18418 = ( n_n5319 ) | ( n_n47  &  wire151 ) ;
 assign wire18420 = ( wire3312 ) | ( wire3313 ) | ( wire18418 ) ;
 assign wire18422 = ( wire18409 ) | ( wire18414 ) | ( _31221 ) ;
 assign wire18429 = ( n_n5111 ) | ( _3109 ) | ( _3110 ) ;
 assign wire18433 = ( wire3353 ) | ( _31186 ) ;
 assign wire18434 = ( n_n5113 ) | ( _31193 ) | ( n_n46  &  wire868 ) ;
 assign wire18445 = ( n_n41  &  n_n83 ) | ( n_n41  &  n_n171 ) | ( n_n41  &  wire1544 ) ;
 assign wire18452 = ( wire18445 ) | ( _2970 ) | ( _31272 ) | ( _31276 ) ;
 assign wire18471 = ( n_n41  &  n_n214 ) | ( n_n41  &  n_n210 ) | ( n_n41  &  n_n107 ) ;
 assign wire18474 = ( n_n5319 ) | ( wire725  &  n_n177  &  n_n46 ) ;
 assign wire18475 = ( wire3271 ) | ( wire18471 ) | ( wire18474 ) ;
 assign wire18476 = ( _2981 ) | ( n_n47  &  wire1425 ) ;
 assign wire18482 = ( wire361 ) | ( n_n41  &  wire1493 ) ;
 assign wire18487 = ( wire3264 ) | ( wire18475 ) | ( wire18476 ) | ( wire18482 ) ;
 assign wire18488 = ( wire18452 ) | ( _2976 ) | ( _31264 ) | ( _31278 ) ;
 assign wire18492 = ( n_n7263 ) | ( n_n7265 ) | ( n_n7264 ) ;
 assign wire18493 = ( wire711 ) | ( n_n10  &  wire729  &  n_n191 ) ;
 assign wire18495 = ( wire18492 ) | ( wire18493 ) | ( _2938 ) ;
 assign wire18496 = ( wire529 ) | ( n_n9  &  wire77 ) | ( wire77  &  n_n6 ) ;
 assign wire18504 = ( n_n3276 ) | ( n_n2948 ) | ( _31302 ) ;
 assign wire18507 = ( n_n231 ) | ( wire18504 ) | ( _31318 ) | ( _31319 ) ;
 assign wire18509 = ( n_n5144 ) | ( n_n159  &  n_n218  &  n_n18 ) ;
 assign wire18510 = ( wire18509 ) | ( wire717  &  n_n149  &  n_n3 ) ;
 assign wire18533 = ( wire3219 ) | ( wire3222 ) | ( wire3223 ) ;
 assign wire18537 = ( n_n184  &  wire719 ) | ( wire719  &  n_n199 ) | ( wire728  &  n_n199 ) ;
 assign wire18541 = ( n_n2859 ) | ( n_n125  &  wire1395 ) ;
 assign wire18546 = ( wire133  &  n_n123 ) | ( n_n123  &  wire959 ) ;
 assign wire18548 = ( wire18533 ) | ( wire18541 ) | ( _31365 ) ;
 assign wire18562 = ( _31376 ) | ( _31377 ) ;
 assign wire18564 = ( n_n5144 ) | ( n_n53  &  n_n123 ) | ( wire157  &  n_n123 ) ;
 assign wire18575 = ( n_n212  &  wire48 ) | ( n_n197  &  wire181 ) ;
 assign wire18576 = ( n_n212  &  wire63 ) | ( n_n212  &  wire52 ) | ( n_n212  &  wire129 ) ;
 assign wire18586 = ( n_n197  &  wire52 ) | ( n_n212  &  wire130 ) ;
 assign wire18587 = ( wire127  &  n_n197 ) | ( n_n197  &  wire129 ) ;
 assign wire18588 = ( wire137  &  n_n212 ) | ( n_n212  &  wire46 ) ;
 assign wire18596 = ( n_n134  &  n_n197 ) | ( n_n212  &  wire186 ) ;
 assign wire18598 = ( n_n197  &  wire125 ) | ( wire725  &  n_n197  &  n_n216 ) ;
 assign wire18600 = ( n_n197  &  wire176 ) | ( n_n212  &  wire125 ) ;
 assign wire18602 = ( n_n4686 ) | ( wire704 ) | ( wire18598 ) ;
 assign wire18603 = ( wire3154 ) | ( wire3155 ) | ( wire18600 ) ;
 assign wire18605 = ( wire158  &  n_n197 ) | ( wire133  &  n_n197 ) ;
 assign wire18607 = ( _31423 ) | ( n_n197  &  wire134 ) | ( n_n197  &  wire156 ) ;
 assign wire18608 = ( wire532 ) | ( wire18605 ) | ( n_n197  &  wire123 ) ;
 assign wire18614 = ( wire689 ) | ( wire3142 ) | ( wire18596 ) ;
 assign wire18616 = ( wire18602 ) | ( wire18603 ) | ( wire18607 ) | ( wire18608 ) ;
 assign wire18619 = ( n_n5144 ) | ( wire725  &  n_n156  &  n_n212 ) ;
 assign wire18631 = ( wire672 ) | ( wire3123 ) | ( n_n43  &  n_n59 ) ;
 assign wire18632 = ( wire3124 ) | ( wire4102 ) | ( n_n43  &  wire222 ) ;
 assign wire18637 = ( n_n101  &  wire224 ) | ( n_n101  &  wire250 ) | ( n_n101  &  wire57 ) ;
 assign wire18638 = ( wire4735 ) | ( wire18637 ) | ( n_n108  &  wire69 ) ;
 assign wire18641 = ( wire4839 ) | ( wire17469 ) | ( _31450 ) ;
 assign wire18642 = ( wire3113 ) | ( n_n101  &  wire218 ) | ( n_n101  &  wire141 ) ;
 assign wire18646 = ( n_n184  &  wire719 ) | ( wire725  &  n_n191 ) ;
 assign wire18650 = ( n_n4981 ) | ( _2737 ) | ( _2738 ) ;
 assign wire18652 = ( n_n5000 ) | ( wire511 ) | ( n_n101  &  wire84 ) ;
 assign wire18655 = ( wire3102 ) | ( wire18652 ) | ( _31445 ) | ( _31446 ) ;
 assign wire18656 = ( wire3111 ) | ( wire18641 ) | ( wire18642 ) | ( wire18650 ) ;
 assign wire18663 = ( n_n5021 ) | ( n_n101  &  wire1723 ) ;
 assign wire18665 = ( n_n5739 ) | ( wire440 ) | ( wire760 ) ;
 assign wire18668 = ( n_n4904 ) | ( n_n5037 ) | ( wire657 ) | ( wire18665 ) ;
 assign wire18669 = ( n_n5033 ) | ( n_n4900 ) | ( wire4937 ) ;
 assign wire18670 = ( wire4935 ) | ( wire18668 ) | ( n_n108  &  wire1844 ) ;
 assign wire18671 = ( wire18663 ) | ( wire18669 ) | ( _2726 ) | ( _31468 ) ;
 assign wire18677 = ( n_n5019 ) | ( n_n101  &  wire1689 ) ;
 assign wire18679 = ( n_n101  &  wire208 ) | ( n_n101  &  wire225 ) | ( n_n101  &  wire148 ) ;
 assign wire18688 = ( n_n5144 ) | ( wire719  &  n_n191  &  n_n42 ) ;
 assign wire18691 = ( wire3068 ) | ( wire3080 ) | ( wire3081 ) | ( wire18688 ) ;
 assign wire18692 = ( wire662 ) | ( wire3069 ) | ( wire3078 ) | ( wire3079 ) ;
 assign wire18694 = ( n_n4755 ) | ( wire18631 ) | ( wire18632 ) ;
 assign wire18701 = ( n_n7240 ) | ( n_n7252 ) | ( wire3060 ) ;
 assign wire18702 = ( n_n7242 ) | ( n_n7254 ) | ( n_n7248 ) | ( wire3059 ) ;
 assign wire18703 = ( i_7_  &  i_6_  &  n_n219  &  n_n111 ) | ( (~ i_7_)  &  i_6_  &  n_n219  &  n_n111 ) ;
 assign wire18704 = ( n_n219  &  n_n218  &  n_n18 ) | ( n_n219  &  n_n48  &  n_n18 ) ;
 assign wire18705 = ( n_n16  &  n_n219  &  n_n218 ) | ( n_n16  &  n_n219  &  n_n48 ) ;
 assign wire18709 = ( wire3044 ) | ( wire245  &  n_n41 ) ;
 assign wire18714 = ( n_n9  &  n_n74 ) | ( n_n10  &  wire1389 ) | ( n_n9  &  wire1389 ) ;
 assign wire18715 = ( n_n6  &  wire344 ) | ( n_n12  &  wire1390 ) ;
 assign wire18718 = ( wire3066 ) | ( wire3067 ) | ( wire18714 ) | ( wire18715 ) ;
 assign wire18726 = ( n_n1408 ) | ( n_n30  &  wire789 ) ;
 assign wire18732 = ( n_n1426 ) | ( n_n30  &  wire791 ) ;
 assign wire18735 = ( n_n1416 ) | ( n_n30  &  wire793 ) ;
 assign wire18737 = ( wire18732 ) | ( wire18735 ) | ( _2581 ) | ( _31594 ) ;
 assign wire18749 = ( n_n1442 ) | ( wire18300 ) | ( _31615 ) ;
 assign wire18750 = ( wire3006 ) | ( n_n31  &  wire863 ) ;
 assign wire18755 = ( n_n1434 ) | ( wire3001 ) | ( wire3015 ) ;
 assign wire18757 = ( wire3013 ) | ( wire3014 ) | ( wire18749 ) | ( wire18750 ) ;
 assign wire18760 = ( n_n33  &  wire48 ) | ( wire130  &  n_n32 ) ;
 assign wire18761 = ( wire675 ) | ( n_n2733 ) | ( wire1417  &  n_n32 ) ;
 assign wire18763 = ( n_n101  &  wire381 ) | ( n_n32  &  wire124 ) ;
 assign wire18767 = ( wire3078 ) | ( wire3079 ) | ( wire3080 ) | ( wire3081 ) ;
 assign wire18768 = ( wire587 ) | ( wire564 ) | ( wire566 ) | ( wire670 ) ;
 assign wire18770 = ( wire2995 ) | ( wire18760 ) | ( wire18761 ) | ( wire18768 ) ;
 assign wire18776 = ( wire3996 ) | ( n_n31  &  wire172 ) | ( n_n31  &  n_n138 ) ;
 assign wire18777 = ( wire2981 ) | ( n_n30  &  wire1021 ) ;
 assign wire18786 = ( n_n4240 ) | ( wire2970 ) | ( n_n31  &  wire144 ) ;
 assign wire18788 = ( wire2964 ) | ( wire2974 ) | ( wire2975 ) ;
 assign wire18793 = ( wire18757 ) | ( wire18770 ) | ( _31632 ) ;
 assign wire18801 = ( wire446 ) | ( wire4252 ) | ( wire4253 ) ;
 assign wire18804 = ( n_n5144 ) | ( n_n6266 ) | ( n_n6268 ) | ( n_n6005 ) ;
 assign wire18812 = ( n_n5319 ) | ( n_n4  &  wire729  &  n_n156 ) ;
 assign wire18815 = ( wire2952 ) | ( wire2958 ) | ( wire2959 ) | ( wire18812 ) ;
 assign wire18816 = ( n_n5319 ) | ( n_n2  &  wire95 ) ;
 assign wire18826 = ( n_n34  &  n_n133 ) | ( n_n36  &  wire1247 ) | ( n_n34  &  wire1247 ) ;
 assign wire18828 = ( wire2939 ) | ( wire2940 ) | ( wire18826 ) ;
 assign wire18833 = ( n_n159  &  n_n218  &  wire747 ) ;
 assign wire18837 = ( wire551 ) | ( wire725  &  n_n191  &  wire18833 ) ;
 assign wire18838 = ( n_n51  &  wire18298 ) | ( n_n30  &  n_n129 ) ;
 assign wire18839 = ( wire428 ) | ( wire462 ) | ( n_n7264 ) ;
 assign wire18841 = ( wire18837 ) | ( wire18838 ) | ( wire18839 ) ;
 assign wire18845 = ( n_n31  &  wire321 ) | ( n_n31  &  wire1285 ) | ( n_n30  &  wire1285 ) ;
 assign wire18846 = ( wire18841 ) | ( wire18845 ) | ( _32149 ) ;
 assign wire18850 = ( n_n41  &  n_n115 ) | ( n_n40  &  n_n115 ) | ( n_n40  &  wire989 ) ;
 assign wire18854 = ( n_n40  &  n_n129 ) | ( n_n38  &  n_n82 ) ;
 assign wire18855 = ( n_n127  &  wire190 ) | ( n_n166  &  wire334 ) ;
 assign wire18871 = ( n_n34  &  n_n95 ) | ( n_n34  &  wire74 ) | ( n_n34  &  wire364 ) ;
 assign wire18877 = ( n_n34  &  wire1579 ) | ( n_n36  &  wire1578 ) | ( n_n34  &  wire1578 ) ;
 assign wire18878 = ( n_n201  &  _31977 ) | ( n_n201  &  _31978 ) ;
 assign wire18882 = ( n_n36  &  wire133 ) | ( n_n36  &  wire376 ) | ( n_n36  &  wire18878 ) ;
 assign wire18883 = ( wire2875 ) | ( n_n34  &  wire133 ) | ( n_n34  &  wire123 ) ;
 assign wire18884 = ( wire18877 ) | ( wire18882 ) | ( n_n36  &  wire1580 ) ;
 assign wire18885 = ( n_n36  &  wire313 ) | ( n_n184  &  wire729  &  n_n36 ) ;
 assign wire18889 = ( n_n36  &  wire52 ) | ( n_n34  &  wire52 ) ;
 assign wire18890 = ( wire2865 ) | ( wire2866 ) ;
 assign wire18891 = ( n_n3638 ) | ( wire2870 ) | ( wire18885 ) | ( wire18889 ) ;
 assign wire18895 = ( n_n36  &  wire147 ) | ( n_n34  &  n_n77 ) ;
 assign wire18911 = ( n_n212  &  wire319 ) | ( n_n197  &  wire1135 ) | ( n_n212  &  wire1135 ) ;
 assign wire18913 = ( n_n117  &  n_n125 ) | ( n_n102  &  n_n123 ) ;
 assign wire18914 = ( n_n123  &  wire313 ) | ( n_n125  &  wire383 ) ;
 assign wire18916 = ( n_n125  &  wire52 ) | ( n_n125  &  wire1279 ) | ( n_n123  &  wire1279 ) ;
 assign wire18917 = ( wire18913 ) | ( wire18914 ) | ( n_n123  &  wire52 ) ;
 assign wire18918 = ( wire2842 ) | ( wire2843 ) | ( wire18916 ) ;
 assign wire18919 = ( n_n197  &  n_n139 ) | ( n_n212  &  n_n139 ) | ( n_n212  &  n_n141 ) ;
 assign wire18922 = ( wire2831 ) | ( wire18919 ) | ( wire188  &  n_n131 ) ;
 assign wire18923 = ( wire2828 ) | ( _2270 ) ;
 assign wire18924 = ( n_n197  &  n_n129 ) | ( n_n212  &  n_n129 ) | ( n_n197  &  n_n127 ) | ( n_n212  &  n_n127 ) ;
 assign wire18925 = ( n_n102  &  n_n125 ) | ( n_n123  &  wire74 ) ;
 assign wire18926 = ( n_n125  &  wire74 ) | ( n_n125  &  wire1136 ) | ( n_n123  &  wire1136 ) ;
 assign wire18928 = ( wire2825 ) | ( wire18924 ) | ( wire18926 ) ;
 assign wire18930 = ( wire18917 ) | ( wire18918 ) | ( wire18922 ) | ( wire18923 ) ;
 assign wire18931 = ( n_n125  &  wire376 ) | ( wire729  &  n_n156  &  n_n125 ) ;
 assign wire18932 = ( wire133  &  n_n123 ) | ( n_n123  &  wire904 ) ;
 assign wire18934 = ( n_n125  &  n_n115 ) | ( n_n123  &  n_n115 ) | ( n_n125  &  wire1242 ) ;
 assign wire18936 = ( wire2808 ) | ( wire2809 ) | ( wire18931 ) | ( wire18932 ) ;
 assign wire18941 = ( n_n113  &  n_n122 ) | ( wire255  &  n_n131 ) ;
 assign wire18943 = ( wire2791 ) | ( wire2801 ) | ( wire2802 ) | ( wire18941 ) ;
 assign wire18947 = ( wire147  &  n_n125 ) | ( n_n77  &  n_n123 ) ;
 assign wire18949 = ( wire2814 ) | ( wire2815 ) | ( wire18947 ) ;
 assign wire18951 = ( wire18936 ) | ( wire18943 ) | ( _31801 ) ;
 assign wire18955 = ( n_n101  &  n_n115 ) | ( n_n108  &  n_n115 ) | ( n_n101  &  wire1470 ) ;
 assign wire18965 = ( n_n101  &  n_n129 ) | ( n_n101  &  n_n127 ) | ( n_n108  &  n_n127 ) ;
 assign wire18968 = ( n_n42  &  wire257 ) | ( n_n43  &  wire313 ) ;
 assign wire18969 = ( n_n42  &  n_n117 ) | ( n_n43  &  n_n117 ) | ( n_n43  &  wire139 ) ;
 assign wire18970 = ( n_n43  &  n_n89 ) | ( n_n47  &  n_n129 ) ;
 assign wire18971 = ( n_n46  &  wire1754 ) | ( n_n47  &  wire1753 ) | ( n_n46  &  wire1753 ) ;
 assign wire18972 = ( n_n43  &  wire257 ) | ( n_n42  &  wire313 ) ;
 assign wire18973 = ( n_n43  &  wire52 ) | ( n_n42  &  wire139 ) ;
 assign wire18976 = ( wire18968 ) | ( wire18969 ) | ( wire18970 ) | ( wire18971 ) ;
 assign wire18985 = ( wire18976 ) | ( _2056 ) | ( _32068 ) | ( _32081 ) ;
 assign wire18991 = ( wire2748 ) | ( n_n101  &  wire1194 ) | ( n_n101  &  wire1497 ) ;
 assign wire18998 = ( wire2740 ) | ( wire2743 ) | ( wire2744 ) ;
 assign wire19003 = ( wire2733 ) | ( wire2738 ) | ( wire2739 ) ;
 assign wire19005 = ( wire18991 ) | ( wire18998 ) | ( _32108 ) ;
 assign wire19010 = ( wire2726 ) | ( wire2728 ) | ( wire2729 ) ;
 assign wire19011 = ( n_n42  &  n_n89 ) | ( n_n41  &  n_n107 ) ;
 assign wire19015 = ( wire2717 ) | ( wire2720 ) | ( wire2721 ) | ( wire19011 ) ;
 assign wire19025 = ( wire18930 ) | ( _31833 ) | ( _31834 ) | ( _31887 ) ;
 assign wire19027 = ( wire18985 ) | ( wire19005 ) | ( _32110 ) ;
 assign wire19031 = ( wire708 ) | ( wire473 ) | ( wire2914 ) | ( wire2915 ) ;
 assign wire19034 = ( n_n1811 ) | ( wire2943 ) | ( wire2944 ) | ( wire18828 ) ;
 assign wire19048 = ( n_n71  &  n_n36 ) | ( n_n34  &  wire133 ) ;
 assign wire19050 = ( wire542 ) | ( wire2692 ) | ( wire19048 ) ;
 assign wire19054 = ( n_n36  &  wire850 ) | ( n_n34  &  wire849 ) ;
 assign wire19057 = ( wire2700 ) | ( wire19050 ) | ( _32649 ) ;
 assign wire19062 = ( wire397 ) | ( n_n3417 ) | ( n_n1553 ) ;
 assign wire19063 = ( wire2679 ) | ( n_n41  &  wire1152 ) ;
 assign wire19069 = ( n_n3419 ) | ( wire500 ) | ( n_n40  &  wire1153 ) ;
 assign wire19076 = ( wire2676 ) | ( wire19062 ) | ( wire19063 ) | ( wire19069 ) ;
 assign wire19077 = ( n_n42  &  n_n89 ) | ( n_n43  &  wire65 ) ;
 assign wire19078 = ( n_n41  &  n_n214 ) | ( n_n41  &  n_n107 ) | ( n_n41  &  n_n202 ) ;
 assign wire19079 = ( n_n42  &  n_n115 ) | ( n_n42  &  n_n136 ) | ( n_n43  &  n_n136 ) ;
 assign wire19083 = ( n_n4622 ) | ( n_n3421 ) | ( n_n1566 ) | ( wire2657 ) ;
 assign wire19084 = ( wire2666 ) | ( wire19077 ) | ( wire19078 ) | ( wire19079 ) ;
 assign wire19087 = ( n_n43  &  n_n89 ) | ( n_n42  &  wire139 ) ;
 assign wire19089 = ( wire19087 ) | ( n_n42  &  wire54 ) | ( n_n42  &  wire357 ) ;
 assign wire19090 = ( n_n4808 ) | ( n_n1575 ) | ( n_n43  &  wire1297 ) ;
 assign wire19098 = ( wire19083 ) | ( wire19084 ) | ( wire19089 ) | ( wire19090 ) ;
 assign wire19103 = ( n_n6267 ) | ( n_n47  &  wire1499 ) ;
 assign wire19104 = ( n_n177  &  wire721 ) | ( n_n177  &  wire728 ) | ( wire721  &  n_n191 ) ;
 assign wire19106 = ( n_n6269 ) | ( wire4252 ) | ( wire4253 ) ;
 assign wire19109 = ( wire19103 ) | ( wire19106 ) | ( _32562 ) ;
 assign wire19118 = ( n_n1594 ) | ( wire2630 ) | ( wire2634 ) | ( wire2635 ) ;
 assign wire19123 = ( n_n46  &  wire852 ) | ( n_n47  &  wire1436 ) ;
 assign wire19125 = ( wire19109 ) | ( wire19118 ) | ( _32577 ) ;
 assign wire19127 = ( wire19076 ) | ( wire19098 ) | ( _32625 ) ;
 assign wire19130 = ( n_n52  &  n_n33 ) | ( n_n136  &  n_n32 ) ;
 assign wire19134 = ( wire473 ) | ( wire2615 ) | ( wire2618 ) | ( wire19130 ) ;
 assign wire19146 = ( _32657 ) | ( n_n30  &  wire925 ) ;
 assign wire19147 = ( n_n1442 ) | ( n_n1170 ) | ( wire2614 ) | ( wire19134 ) ;
 assign wire19148 = ( n_n125  &  wire1287 ) | ( n_n123  &  wire1286 ) ;
 assign wire19153 = ( wire2599 ) | ( wire19148 ) | ( n_n113  &  wire276 ) ;
 assign wire19158 = ( n_n1700 ) | ( wire2594 ) | ( wire133  &  n_n123 ) ;
 assign wire19164 = ( n_n2881 ) | ( n_n1708 ) | ( n_n123  &  wire916 ) ;
 assign wire19169 = ( n_n117  &  n_n125 ) | ( n_n123  &  wire52 ) ;
 assign wire19178 = ( wire2584 ) | ( wire19164 ) | ( wire19169 ) | ( _32351 ) ;
 assign wire19182 = ( n_n184  &  wire729 ) | ( wire727  &  n_n191 ) ;
 assign wire19186 = ( n_n5019 ) | ( n_n108  &  wire1070 ) ;
 assign wire19189 = ( n_n113  &  n_n115 ) | ( n_n108  &  wire111 ) ;
 assign wire19190 = ( wire760 ) | ( wire2567 ) | ( n_n112  &  wire65 ) ;
 assign wire19193 = ( n_n5033 ) | ( wire2568 ) | ( wire19189 ) ;
 assign wire19200 = ( n_n5021 ) | ( wire2560 ) | ( wire2565 ) ;
 assign wire19202 = ( wire19186 ) | ( wire19193 ) | ( _32380 ) ;
 assign wire19208 = ( wire2557 ) | ( wire2559 ) | ( _32304 ) ;
 assign wire19210 = ( wire19153 ) | ( wire19158 ) | ( _32327 ) ;
 assign wire19212 = ( wire19178 ) | ( wire19202 ) | ( _32382 ) ;
 assign wire19213 = ( n_n212  &  n_n127 ) | ( n_n197  &  wire83 ) ;
 assign wire19216 = ( n_n184  &  wire720 ) | ( wire729  &  n_n216 ) ;
 assign wire19220 = ( n_n212  &  wire63 ) | ( n_n212  &  wire1145 ) ;
 assign wire19227 = ( n_n197  &  wire52 ) | ( n_n212  &  wire1147 ) ;
 assign wire19232 = ( wire2532 ) | ( n_n212  &  wire1150 ) ;
 assign wire19234 = ( wire19220 ) | ( wire19227 ) | ( _32426 ) ;
 assign wire19238 = ( n_n102  &  n_n123 ) | ( n_n125  &  wire51 ) ;
 assign wire19239 = ( wire142  &  n_n123 ) | ( n_n125  &  wire52 ) ;
 assign wire19241 = ( wire2526 ) | ( n_n125  &  wire1255 ) ;
 assign wire19249 = ( wire2523 ) | ( wire2525 ) | ( _32408 ) ;
 assign wire19256 = ( wire127  &  n_n197 ) | ( n_n212  &  wire1289 ) ;
 assign wire19263 = ( _1516 ) | ( _1517 ) | ( wire133  &  _32447 ) ;
 assign wire19268 = ( wire126  &  n_n212 ) | ( wire147  &  n_n212 ) | ( n_n212  &  wire1293 ) ;
 assign wire19270 = ( wire19256 ) | ( wire19263 ) | ( _32450 ) ;
 assign wire19272 = ( n_n123  &  wire74 ) | ( n_n123  &  wire68 ) | ( n_n123  &  wire81 ) ;
 assign wire19273 = ( n_n4674 ) | ( wire2498 ) | ( n_n102  &  n_n125 ) ;
 assign wire19276 = ( wire19241 ) | ( wire19249 ) | ( _32410 ) ;
 assign wire19278 = ( wire19234 ) | ( wire19270 ) | ( _32452 ) ;
 assign wire19281 = ( n_n170  &  wire727 ) | ( n_n170  &  wire717 ) ;
 assign wire19285 = ( wire685 ) | ( n_n101  &  wire250 ) ;
 assign wire19286 = ( wire2493 ) | ( _1845 ) | ( _1846 ) ;
 assign wire19294 = ( n_n5000 ) | ( wire2490 ) | ( n_n108  &  wire234 ) ;
 assign wire19301 = ( wire2487 ) | ( _32230 ) | ( wire384  &  _32227 ) ;
 assign wire19302 = ( wire2489 ) | ( wire19285 ) | ( wire19286 ) | ( wire19294 ) ;
 assign wire19304 = ( n_n6005 ) | ( wire419 ) | ( n_n101  &  n_n129 ) ;
 assign wire19306 = ( wire729  &  n_n216 ) | ( wire717  &  n_n216 ) | ( wire726  &  n_n216 ) ;
 assign wire19307 = ( n_n108  &  n_n129 ) | ( n_n101  &  wire378 ) ;
 assign wire19308 = ( n_n46  &  wire1343 ) | ( wire1345  &  wire1342 ) ;
 assign wire19309 = ( wire19307 ) | ( n_n47  &  wire162 ) | ( n_n47  &  wire19306 ) ;
 assign wire19310 = ( n_n1624 ) | ( wire2475 ) | ( wire19304 ) | ( wire19308 ) ;
 assign wire19316 = ( wire2464 ) | ( n_n101  &  wire90 ) ;
 assign wire19317 = ( wire2463 ) | ( wire2468 ) | ( n_n101  &  wire1405 ) ;
 assign wire19324 = ( wire2462 ) | ( n_n46  &  wire1214 ) | ( n_n46  &  wire1581 ) ;
 assign wire19325 = ( n_n4641 ) | ( wire693 ) | ( wire19324 ) ;
 assign wire19326 = ( wire19309 ) | ( wire19310 ) | ( wire19316 ) | ( wire19317 ) ;
 assign wire19332 = ( n_n5113 ) | ( n_n1606 ) | ( wire2451 ) ;
 assign wire19338 = ( wire498 ) | ( wire2448 ) ;
 assign wire19343 = ( n_n5111 ) | ( wire137  &  n_n46 ) | ( wire146  &  n_n46 ) ;
 assign wire19344 = ( wire2442 ) | ( n_n47  &  wire1216 ) ;
 assign wire19346 = ( wire2449 ) | ( wire2452 ) | ( wire19332 ) | ( wire19338 ) ;
 assign wire19347 = ( wire19301 ) | ( wire19302 ) | ( wire19325 ) | ( wire19326 ) ;
 assign wire19351 = ( n_n36  &  n_n102 ) | ( n_n34  &  wire81 ) ;
 assign wire19354 = ( wire17541 ) | ( _32677 ) | ( wire68  &  _32675 ) ;
 assign wire19355 = ( wire2435 ) | ( wire19351 ) | ( n_n38  &  wire248 ) ;
 assign wire19359 = ( n_n39  &  wire248 ) | ( n_n39  &  wire249 ) ;
 assign wire19362 = ( n_n1517 ) | ( wire457 ) | ( wire19359 ) ;
 assign wire19363 = ( n_n1520 ) | ( wire572 ) | ( wire2427 ) | ( wire2428 ) ;
 assign wire19364 = ( n_n36  &  wire98 ) | ( n_n34  &  n_n102 ) ;
 assign wire19366 = ( n_n34  &  wire74 ) | ( n_n36  &  n_n198 ) ;
 assign wire19368 = ( wire2418 ) | ( wire2424 ) | ( wire19364 ) ;
 assign wire19369 = ( wire2417 ) | ( wire19366 ) | ( wire19368 ) ;
 assign wire19370 = ( wire19354 ) | ( wire19355 ) | ( wire19362 ) | ( wire19363 ) ;
 assign wire19376 = ( n_n1426 ) | ( n_n30  &  wire913 ) ;
 assign wire19380 = ( n_n1416 ) | ( n_n31  &  wire126 ) | ( n_n31  &  wire147 ) ;
 assign wire19381 = ( wire2410 ) | ( n_n30  &  wire1069 ) ;
 assign wire19389 = ( wire2415 ) | ( wire19376 ) | ( wire19380 ) | ( wire19381 ) ;
 assign wire19393 = ( n_n36  &  _32478 ) | ( wire720  &  n_n36  &  _29155 ) ;
 assign wire19395 = ( wire19393 ) | ( n_n34  &  wire63 ) | ( n_n34  &  wire52 ) ;
 assign wire19396 = ( wire2398 ) | ( n_n34  &  wire1077 ) ;
 assign wire19400 = ( n_n36  &  wire52 ) | ( n_n34  &  n_n183 ) ;
 assign wire19401 = ( wire19400 ) | ( n_n36  &  wire63 ) ;
 assign wire19402 = ( wire2393 ) | ( n_n36  &  wire1079 ) ;
 assign wire19403 = ( n_n34  &  _32474 ) | ( wire729  &  n_n34  &  _29755 ) ;
 assign wire19405 = ( n_n36  &  wire126 ) | ( n_n36  &  wire53 ) | ( n_n36  &  wire69 ) ;
 assign wire19406 = ( wire2384 ) | ( wire19403 ) | ( n_n36  &  wire147 ) ;
 assign wire19409 = ( wire19395 ) | ( wire19396 ) | ( wire19401 ) | ( wire19402 ) ;
 assign wire19423 = ( n_n6492 ) | ( n_n3413 ) | ( n_n1542 ) | ( wire2374 ) ;
 assign wire19429 = ( wire2370 ) | ( wire2372 ) | ( _32510 ) ;
 assign wire19431 = ( wire2382 ) | ( wire19423 ) | ( _32526 ) | ( _32529 ) ;
 assign wire19437 = ( n_n1408 ) | ( n_n30  &  wire1504 ) ;
 assign wire19454 = ( wire19146 ) | ( wire19147 ) | ( wire19369 ) | ( wire19370 ) ;
 assign wire19455 = ( wire19389 ) | ( wire19409 ) | ( _32488 ) ;
 assign wire19456 = ( wire19431 ) | ( wire19437 ) | ( _32540 ) | ( _32541 ) ;
 assign wire19466 = ( wire2345 ) | ( wire2349 ) | ( n_n31  &  wire1012 ) ;
 assign wire19471 = ( wire2340 ) | ( wire2343 ) | ( wire2344 ) ;
 assign wire19479 = ( wire19466 ) | ( wire19471 ) | ( _33138 ) ;
 assign wire19485 = ( n_n36  &  wire1708 ) | ( n_n36  &  wire1707 ) | ( n_n34  &  wire1707 ) ;
 assign wire19491 = ( wire2323 ) | ( wire19485 ) | ( n_n34  &  wire1709 ) ;
 assign wire19494 = ( n_n156  &  wire719  &  n_n34 ) | ( n_n177  &  wire719  &  n_n34 ) ;
 assign wire19496 = ( n_n33  &  wire48 ) | ( n_n32  &  wire124 ) ;
 assign wire19497 = ( wire226  &  n_n128 ) | ( n_n32  &  wire165 ) ;
 assign wire19498 = ( wire19494 ) | ( wire19496 ) | ( n_n36  &  wire1738 ) ;
 assign wire19499 = ( wire19497 ) | ( n_n33  &  wire1739 ) ;
 assign wire19513 = ( n_n212  &  wire48 ) | ( n_n212  &  wire151 ) ;
 assign wire19520 = ( n_n36  &  wire219 ) | ( wire720  &  n_n36  &  n_n199 ) ;
 assign wire19521 = ( n_n36  &  wire100 ) | ( n_n177  &  wire720  &  n_n36 ) ;
 assign wire19527 = ( wire2287 ) | ( wire19521 ) | ( n_n36  &  wire1605 ) ;
 assign wire19536 = ( n_n38  &  n_n134 ) | ( n_n39  &  n_n132 ) ;
 assign wire19538 = ( wire2269 ) | ( wire19536 ) | ( n_n34  &  n_n198 ) ;
 assign wire19539 = ( wire2290 ) | ( wire2293 ) | ( wire2294 ) | ( wire19520 ) ;
 assign wire19541 = ( wire2277 ) | ( wire2278 ) | ( wire19527 ) | ( _33013 ) ;
 assign wire19542 = ( n_n41  &  n_n130 ) | ( n_n39  &  wire104 ) ;
 assign wire19543 = ( n_n40  &  wire1160 ) | ( n_n41  &  wire1159 ) | ( n_n40  &  wire1159 ) ;
 assign wire19544 = ( n_n40  &  n_n138 ) | ( n_n41  &  n_n142 ) ;
 assign wire19545 = ( n_n41  &  n_n140 ) | ( n_n40  &  n_n140 ) | ( n_n40  &  wire407 ) ;
 assign wire19548 = ( n_n4602 ) | ( wire19542 ) | ( wire19543 ) | ( wire19544 ) ;
 assign wire19549 = ( wire4863 ) | ( wire19545 ) | ( _32808 ) ;
 assign wire19552 = ( n_n38  &  wire110 ) | ( n_n38  &  n_n177  &  wire719 ) ;
 assign wire19567 = ( n_n42  &  n_n138 ) | ( n_n41  &  n_n210 ) ;
 assign wire19576 = ( i_9_  &  (~ i_10_)  &  i_11_  &  wire719 ) | ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire719 ) | ( (~ i_9_)  &  (~ i_10_)  &  (~ i_11_)  &  wire719 ) ;
 assign wire19580 = ( n_n47  &  n_n140 ) | ( n_n46  &  n_n140 ) | ( n_n47  &  n_n142 ) ;
 assign wire19581 = ( n_n47  &  wire55 ) | ( n_n46  &  wire134 ) ;
 assign wire19589 = ( n_n6266 ) | ( n_n6268 ) | ( n_n43  &  wire107 ) ;
 assign wire19603 = ( n_n108  &  wire401 ) | ( wire719  &  n_n216  &  n_n108 ) ;
 assign wire19610 = ( wire445 ) | ( wire719  &  n_n170  &  wire228 ) ;
 assign wire19612 = ( wire2190 ) | ( wire2195 ) | ( wire2197 ) | ( wire19603 ) ;
 assign wire19613 = ( wire446 ) | ( wire4827 ) | ( wire4828 ) ;
 assign wire19623 = ( wire2176 ) | ( wire2179 ) | ( wire2180 ) ;
 assign wire19629 = ( wire2174 ) | ( n_n101  &  wire1706 ) | ( n_n101  &  wire1740 ) ;
 assign wire19636 = ( wire2169 ) | ( n_n108  &  wire1742 ) | ( n_n108  &  wire1756 ) ;
 assign wire19638 = ( wire19623 ) | ( wire19629 ) | ( _33048 ) ;
 assign wire19644 = ( n_n125  &  n_n142 ) | ( n_n125  &  n_n116 ) | ( n_n123  &  n_n116 ) ;
 assign wire19645 = ( wire2157 ) | ( wire19644 ) ;
 assign wire19646 = ( wire2163 ) | ( n_n123  &  wire856 ) | ( n_n123  &  wire859 ) ;
 assign wire19647 = ( n_n113  &  n_n116 ) | ( n_n112  &  wire1084 ) ;
 assign wire19648 = ( i_15_  &  n_n184  &  n_n207 ) | ( (~ i_15_)  &  n_n184  &  n_n207 ) | ( i_15_  &  n_n184  &  n_n215 ) ;
 assign wire19650 = ( n_n132  &  n_n125 ) | ( n_n132  &  n_n123 ) | ( n_n123  &  wire1087 ) ;
 assign wire19652 = ( wire19650 ) | ( n_n113  &  wire107 ) | ( n_n113  &  wire19648 ) ;
 assign wire19653 = ( wire2146 ) | ( wire2149 ) | ( wire2153 ) | ( wire19647 ) ;
 assign wire19656 = ( wire2141 ) | ( wire2155 ) | ( wire2156 ) ;
 assign wire19658 = ( wire19645 ) | ( wire19646 ) | ( wire19652 ) | ( wire19653 ) ;
 assign wire19659 = ( n_n197  &  n_n130 ) | ( n_n212  &  n_n130 ) | ( n_n197  &  n_n128 ) | ( n_n212  &  n_n128 ) ;
 assign wire19666 = ( wire2136 ) | ( n_n125  &  wire1259 ) | ( n_n125  &  wire1260 ) ;
 assign wire19667 = ( n_n197  &  n_n140 ) | ( n_n212  &  n_n140 ) | ( n_n212  &  n_n142 ) ;
 assign wire19668 = ( n_n134  &  n_n197 ) | ( wire55  &  n_n212 ) ;
 assign wire19670 = ( wire2124 ) | ( wire2130 ) | ( wire19667 ) ;
 assign wire19671 = ( wire2125 ) | ( wire19668 ) | ( n_n132  &  wire188 ) ;
 assign wire19674 = ( wire2119 ) | ( wire2139 ) | ( wire19659 ) ;
 assign wire19676 = ( wire2134 ) | ( wire19666 ) | ( wire19670 ) | ( wire19671 ) ;
 assign wire19677 = ( n_n752 ) | ( wire19538 ) | ( wire19539 ) | ( wire19541 ) ;
 assign wire19680 = ( wire19638 ) | ( wire19658 ) | ( _33099 ) ;
 assign wire19687 = ( n_n31  &  wire777 ) | ( n_n30  &  wire776 ) ;
 assign wire19691 = ( n_n31  &  wire1416 ) | ( n_n31  &  wire1414 ) | ( n_n30  &  wire1414 ) ;
 assign wire19693 = ( n_n7242 ) | ( n_n156  &  n_n30  &  wire728 ) ;
 assign wire19694 = ( n_n7263 ) | ( n_n3276 ) | ( n_n2948 ) ;
 assign wire19695 = ( n_n52  &  n_n31 ) | ( wire751  &  wire1367 ) ;
 assign wire19698 = ( wire2108 ) | ( wire19691 ) | ( wire19693 ) | ( wire19694 ) ;
 assign wire19702 = ( _635 ) | ( _636 ) | ( n_n41  &  _30974 ) ;
 assign wire19704 = ( n_n41  &  n_n62 ) | ( n_n40  &  n_n62 ) | ( n_n40  &  wire1476 ) ;
 assign wire19706 = ( n_n177  &  wire720 ) | ( n_n170  &  wire720 ) | ( n_n177  &  wire727 ) | ( n_n170  &  wire727 ) ;
 assign wire19707 = ( n_n40  &  n_n58 ) | ( n_n41  &  wire1478 ) | ( n_n40  &  wire1478 ) ;
 assign wire19708 = ( n_n54  &  wire1480 ) | ( n_n38  &  wire1479 ) ;
 assign wire19710 = ( wire19704 ) | ( wire19708 ) | ( n_n41  &  wire1477 ) ;
 assign wire19717 = ( n_n34  &  n_n183 ) | ( n_n36  &  n_n176 ) ;
 assign wire19718 = ( n_n34  &  wire63 ) | ( n_n36  &  wire348 ) ;
 assign wire19722 = ( wire2070 ) | ( wire2078 ) | ( wire2079 ) | ( wire19717 ) ;
 assign wire19725 = ( n_n34  &  wire126 ) | ( n_n34  &  wire933 ) ;
 assign wire19726 = ( wire720  &  n_n149 ) | ( n_n177  &  wire718 ) ;
 assign wire19730 = ( n_n36  &  wire126 ) | ( n_n34  &  n_n176 ) ;
 assign wire19731 = ( wire137  &  n_n34 ) | ( n_n34  &  n_n171 ) | ( n_n34  &  wire19726 ) ;
 assign wire19733 = ( wire2062 ) | ( wire2068 ) | ( wire19725 ) ;
 assign wire19734 = ( n_n36  &  n_n198 ) | ( n_n34  &  wire385 ) ;
 assign wire19735 = ( n_n36  &  wire68 ) | ( n_n34  &  wire68 ) ;
 assign wire19738 = ( n_n369 ) | ( n_n371 ) | ( wire19734 ) | ( wire19735 ) ;
 assign wire19739 = ( wire19722 ) | ( wire19733 ) | ( _33261 ) ;
 assign wire19746 = ( wire720  &  n_n41  &  n_n216 ) | ( n_n41  &  wire726  &  n_n216 ) ;
 assign wire19747 = ( n_n42  &  n_n136 ) | ( n_n43  &  n_n136 ) | ( n_n42  &  n_n60 ) ;
 assign wire19750 = ( n_n41  &  wire296 ) | ( n_n40  &  wire296 ) | ( n_n40  &  wire332 ) ;
 assign wire19752 = ( wire2045 ) | ( wire19746 ) | ( wire19747 ) | ( wire19750 ) ;
 assign wire19756 = ( n_n41  &  wire1617 ) | ( n_n177  &  n_n41  &  wire726 ) ;
 assign wire19757 = ( _33291 ) | ( n_n40  &  wire1684 ) | ( n_n40  &  _33287 ) ;
 assign wire19758 = ( wire2041 ) | ( wire19752 ) | ( wire19756 ) | ( _33293 ) ;
 assign wire19765 = ( wire1992 ) | ( wire1995 ) | ( wire1996 ) ;
 assign wire19769 = ( wire1987 ) | ( wire1990 ) | ( wire1991 ) ;
 assign wire19775 = ( wire1982 ) | ( wire1997 ) | ( wire1998 ) ;
 assign wire19777 = ( wire19765 ) | ( wire19769 ) | ( _33477 ) ;
 assign wire19779 = ( n_n101  &  n_n136 ) | ( n_n108  &  n_n136 ) | ( n_n108  &  wire1357 ) ;
 assign wire19792 = ( n_n6005 ) | ( wire4354 ) | ( wire4355 ) ;
 assign wire19800 = ( n_n43  &  n_n183 ) | ( n_n42  &  wire346 ) ;
 assign wire19801 = ( n_n42  &  wire128 ) | ( n_n43  &  wire128 ) ;
 assign wire19802 = ( n_n42  &  n_n183 ) | ( n_n46  &  n_n58 ) ;
 assign wire19803 = ( i_8_  &  n_n16  &  wire739 ) | ( (~ i_8_)  &  n_n16  &  wire739 ) | ( i_8_  &  n_n16  &  wire759 ) | ( (~ i_8_)  &  n_n16  &  wire759 ) ;
 assign wire19804 = ( n_n43  &  n_n190 ) | ( wire189  &  wire1666 ) ;
 assign wire19807 = ( wire2004 ) | ( wire19802 ) | ( n_n54  &  wire1668 ) ;
 assign wire19808 = ( wire19800 ) | ( wire19801 ) | ( wire19803 ) | ( wire19804 ) ;
 assign wire19813 = ( n_n302 ) | ( wire1983 ) | ( wire19775 ) | ( wire19777 ) ;
 assign wire19823 = ( n_n212  &  wire166 ) | ( n_n197  &  wire1366 ) | ( n_n212  &  wire1366 ) ;
 assign wire19825 = ( n_n197  &  n_n62 ) | ( n_n212  &  n_n62 ) | ( n_n212  &  n_n64 ) ;
 assign wire19828 = ( wire1979 ) | ( wire19825 ) | ( wire188  &  n_n56 ) ;
 assign wire19829 = ( wire1976 ) | ( _217 ) ;
 assign wire19830 = ( n_n54  &  n_n197 ) | ( n_n52  &  n_n197 ) | ( n_n54  &  n_n212 ) | ( n_n52  &  n_n212 ) ;
 assign wire19834 = ( wire1971 ) | ( n_n123  &  wire1510 ) | ( n_n123  &  wire1512 ) ;
 assign wire19837 = ( wire1962 ) | ( wire1972 ) | ( wire19830 ) ;
 assign wire19839 = ( wire1968 ) | ( wire19828 ) | ( wire19829 ) | ( wire19834 ) ;
 assign wire19841 = ( n_n113  &  n_n183 ) | ( wire255  &  n_n56 ) ;
 assign wire19842 = ( n_n125  &  wire1717 ) | ( n_n123  &  wire1716 ) ;
 assign wire19843 = ( i_15_  &  n_n184  &  n_n205 ) | ( (~ i_15_)  &  n_n184  &  n_n205 ) | ( (~ i_15_)  &  n_n184  &  n_n215 ) ;
 assign wire19845 = ( wire63  &  n_n112 ) | ( n_n112  &  wire1720 ) ;
 assign wire19858 = ( wire1940 ) | ( wire1960 ) | ( wire1961 ) ;
 assign wire19861 = ( wire19839 ) | ( _33496 ) | ( _33497 ) | ( _33535 ) ;
 assign wire19867 = ( wire19707 ) | ( wire19710 ) | ( _33185 ) | ( _33220 ) ;
 assign wire19875 = ( n_n34  &  n_n58 ) | ( n_n36  &  n_n56 ) ;
 assign wire19876 = ( n_n54  &  n_n36 ) | ( n_n52  &  n_n36 ) | ( n_n54  &  n_n34 ) | ( n_n52  &  n_n34 ) ;
 assign wire19878 = ( wire1914 ) | ( wire19875 ) | ( wire19876 ) ;
 assign wire19880 = ( n_n52  &  n_n33 ) | ( n_n31  &  wire335 ) ;
 assign wire19884 = ( wire1907 ) | ( wire1910 ) | ( wire1912 ) | ( wire19880 ) ;
 assign wire19886 = ( n_n36  &  wire1778 ) | ( n_n36  &  wire1777 ) | ( n_n34  &  wire1777 ) ;
 assign wire19887 = ( n_n36  &  wire127 ) | ( n_n34  &  wire1780 ) ;
 assign wire19890 = ( wire556 ) | ( n_n34  &  wire156 ) | ( n_n34  &  wire1570 ) ;
 assign wire19891 = ( wire542 ) | ( wire1906 ) | ( wire19886 ) | ( wire19887 ) ;
 assign wire19893 = ( wire19878 ) | ( wire19884 ) | ( _33626 ) ;
 assign wire19898 = ( wire520 ) | ( n_n30  &  wire1311 ) | ( n_n30  &  wire1482 ) ;
 assign wire19904 = ( wire507 ) | ( wire510 ) | ( wire513 ) ;
 assign wire19907 = ( wire499 ) | ( wire552 ) | ( n_n31  &  wire1090 ) ;
 assign wire19909 = ( wire19898 ) | ( wire19904 ) | ( _33578 ) ;
 assign wire19910 = ( n_n5144 ) | ( n_n159  &  n_n218  &  n_n18 ) ;
 assign wire19911 = ( wire19910 ) | ( wire185  &  n_n3 ) ;
 assign wire19917 = ( n_n5144 ) | ( n_n162  &  n_n219  &  n_n18 ) ;
 assign wire19920 = ( wire389 ) | ( wire19917 ) | ( _33670 ) ;
 assign wire19923 = ( n_n5144 ) | ( n_n219  &  n_n111  &  n_n157 ) ;
 assign wire19925 = ( wire388 ) | ( wire267  &  wire781 ) ;
 assign wire19926 = ( n_n3389 ) | ( wire19923 ) | ( n_n135  &  wire783 ) ;
 assign wire19930 = ( i_7_  &  (~ i_6_)  &  n_n219  &  n_n218 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n219  &  n_n218 ) ;
 assign wire19938 = ( wire551 ) | ( wire725  &  n_n191  &  wire18833 ) ;
 assign wire19939 = ( n_n7242 ) | ( wire462 ) | ( wire751  &  n_n59 ) ;
 assign wire19943 = ( n_n5144 ) | ( n_n159  &  n_n218  &  n_n18 ) ;
 assign wire19944 = ( wire19943 ) | ( wire77  &  n_n3 ) ;
 assign _86 = ( n_n5  &  wire95 ) | ( n_n5  &  _33681 ) ;
 assign _87 = ( n_n5  &  wire87 ) | ( n_n5  &  wire729  &  n_n149 ) ;
 assign _143 = ( n_n33  &  wire166 ) | ( n_n33  &  wire283 ) | ( n_n33  &  wire235 ) ;
 assign _217 = ( n_n212  &  wire235 ) | ( n_n212  &  wire236 ) | ( n_n212  &  _33528 ) ;
 assign _252 = ( n_n212  &  wire269 ) | ( n_n212  &  wire275 ) | ( n_n212  &  wire278 ) ;
 assign _255 = ( n_n197  &  wire282 ) | ( n_n197  &  wire236 ) | ( n_n197  &  wire354 ) ;
 assign _285 = ( n_n101  &  wire161 ) | ( n_n101  &  wire337 ) | ( n_n101  &  _288 ) ;
 assign _288 = ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire726 ) ;
 assign _314 = ( n_n108  &  wire110 ) | ( n_n108  &  wire329 ) | ( n_n108  &  _317 ) ;
 assign _317 = ( (~ i_9_)  &  (~ i_10_)  &  i_11_  &  wire726 ) ;
 assign _360 = ( n_n218  &  n_n220  &  n_n126  &  wire1761 ) ;
 assign _409 = ( n_n184  &  wire728  &  wire255 ) ;
 assign _422 = ( wire207  &  n_n123 ) | ( n_n123  &  wire249 ) | ( n_n123  &  _425 ) ;
 assign _425 = ( i_9_  &  i_10_  &  i_11_  &  wire728 ) ;
 assign _453 = ( n_n47  &  wire282 ) | ( n_n47  &  wire283 ) | ( n_n47  &  wire354 ) ;
 assign _461 = ( wire244  &  n_n46 ) | ( wire140  &  n_n46 ) | ( n_n46  &  wire414 ) ;
 assign _462 = ( n_n46  &  wire235 ) | ( n_n46  &  wire236 ) | ( n_n46  &  _465 ) ;
 assign _465 = ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire728 ) ;
 assign _499 = ( n_n41  &  wire166 ) | ( n_n41  &  wire269 ) | ( n_n41  &  wire332 ) ;
 assign _511 = ( n_n40  &  wire282 ) | ( n_n40  &  wire283 ) | ( n_n40  &  wire325 ) ;
 assign _596 = ( n_n124  &  n_n48  &  n_n220  &  wire140 ) ;
 assign _635 = ( wire140  &  n_n40 ) | ( n_n40  &  wire354 ) ;
 assign _636 = ( wire244  &  n_n40 ) | ( n_n40  &  wire235 ) | ( n_n40  &  wire236 ) ;
 assign _696 = ( n_n31  &  wire53 ) | ( n_n31  &  wire237 ) | ( n_n31  &  _699 ) ;
 assign _699 = ( i_9_  &  (~ i_10_)  &  i_11_  &  wire724 ) ;
 assign _745 = ( n_n218  &  n_n220  &  n_n126  &  wire1758 ) ;
 assign _778 = ( n_n162  &  n_n124  &  n_n220  &  wire1743 ) ;
 assign _823 = ( n_n184  &  wire720  &  n_n34 ) ;
 assign _969 = ( n_n48  &  n_n220  &  n_n161  &  wire46 ) ;
 assign _976 = ( wire132  &  n_n47 ) | ( n_n47  &  wire280 ) | ( n_n47  &  wire121 ) ;
 assign _1018 = ( wire132  &  n_n40 ) | ( n_n40  &  wire46 ) | ( n_n40  &  wire121 ) ;
 assign _1021 = ( n_n41  &  wire48 ) | ( n_n41  &  wire167 ) | ( n_n41  &  wire192 ) ;
 assign _1126 = ( n_n34  &  wire215 ) | ( n_n34  &  wire438 ) | ( n_n34  &  _1129 ) ;
 assign _1129 = ( i_9_  &  i_10_  &  (~ i_11_)  &  wire720 ) ;
 assign _1208 = ( n_n31  &  wire63 ) | ( n_n31  &  wire330 ) | ( n_n31  &  _1211 ) ;
 assign _1211 = ( (~ i_9_)  &  i_10_  &  i_11_  &  wire720 ) ;
 assign _1239 = ( n_n36  &  wire155 ) | ( n_n36  &  wire315 ) | ( n_n36  &  wire300 ) ;
 assign _1242 = ( n_n218  &  n_n35  &  n_n220  &  wire1207 ) ;
 assign _1262 = ( n_n33  &  wire118 ) | ( n_n33  &  wire277 ) | ( n_n33  &  _1265 ) ;
 assign _1263 = ( n_n162  &  n_n220  &  n_n200  &  wire274 ) ;
 assign _1264 = ( n_n162  &  n_n220  &  n_n200  &  wire148 ) ;
 assign _1265 = ( (~ i_9_)  &  (~ i_10_)  &  i_11_  &  wire729 ) ;
 assign _1289 = ( n_n40  &  wire142 ) | ( n_n40  &  wire233 ) | ( n_n40  &  wire56 ) ;
 assign _1307 = ( n_n40  &  wire179 ) | ( n_n40  &  wire148 ) | ( n_n40  &  wire274 ) ;
 assign _1308 = ( n_n40  &  wire223 ) | ( n_n40  &  wire239 ) ;
 assign _1347 = ( n_n46  &  wire198 ) | ( n_n46  &  wire175 ) | ( n_n46  &  wire88 ) ;
 assign _1401 = ( n_n31  &  wire52 ) | ( n_n31  &  wire51 ) | ( n_n31  &  wire271 ) ;
 assign _1404 = ( n_n162  &  wire714  &  wire1006  &  _29429 ) ;
 assign _1411 = ( n_n31  &  wire315 ) | ( n_n31  &  wire300 ) | ( n_n31  &  _1414 ) ;
 assign _1414 = ( (~ i_9_)  &  i_10_  &  (~ i_11_)  &  wire720 ) ;
 assign _1455 = ( n_n41  &  wire155 ) | ( n_n41  &  wire50 ) | ( n_n41  &  wire300 ) ;
 assign _1516 = ( n_n212  &  wire49 ) | ( n_n212  &  wire300 ) | ( n_n212  &  _1519 ) ;
 assign _1517 = ( n_n212  &  wire221 ) | ( n_n212  &  wire315 ) ;
 assign _1519 = ( (~ i_9_)  &  i_10_  &  (~ i_11_)  &  wire720 ) ;
 assign _1533 = ( n_n218  &  n_n220  &  n_n200  &  wire1294 ) ;
 assign _1544 = ( n_n197  &  wire142 ) | ( n_n197  &  wire251 ) | ( n_n197  &  wire19216 ) ;
 assign _1549 = ( n_n197  &  wire98 ) | ( n_n197  &  wire254 ) | ( n_n197  &  wire51 ) ;
 assign _1581 = ( n_n218  &  n_n220  &  n_n200  &  wire1257 ) ;
 assign _1643 = ( n_n101  &  wire257 ) | ( n_n101  &  wire271 ) | ( n_n101  &  wire19182 ) ;
 assign _1648 = ( n_n162  &  n_n220  &  n_n126  &  wire1075 ) ;
 assign _1676 = ( wire63  &  n_n123 ) | ( wire98  &  n_n123 ) | ( n_n123  &  wire254 ) ;
 assign _1679 = ( wire126  &  n_n125 ) | ( wire53  &  n_n125 ) | ( n_n125  &  wire239 ) ;
 assign _1721 = ( n_n218  &  n_n220  &  n_n161  &  wire63 ) ;
 assign _1845 = ( n_n108  &  wire281 ) | ( n_n108  &  wire69 ) | ( n_n108  &  wire59 ) ;
 assign _1846 = ( n_n108  &  wire19281 ) | ( n_n108  &  _1848 ) | ( n_n108  &  _1849 ) ;
 assign _1848 = ( i_14_  &  i_13_  &  (~ i_12_)  &  _32240 ) ;
 assign _1849 = ( i_14_  &  i_13_  &  (~ i_12_)  &  _32241 ) ;
 assign _1862 = ( n_n101  &  wire156 ) | ( n_n101  &  wire59 ) | ( n_n101  &  wire300 ) ;
 assign _1871 = ( n_n162  &  n_n220  &  n_n126  &  wire250 ) ;
 assign _1972 = ( n_n2  &  wire95 ) | ( n_n2  &  _32140 ) ;
 assign _1978 = ( n_n162  &  wire714  &  wire1197  &  _29429 ) ;
 assign _1990 = ( n_n162  &  wire714  &  wire993  &  _29429 ) ;
 assign _1992 = ( n_n30  &  wire321 ) | ( n_n30  &  _32115 ) ;
 assign _1993 = ( n_n30  &  wire302 ) | ( n_n30  &  wire303 ) | ( n_n30  &  wire316 ) ;
 assign _2020 = ( n_n108  &  wire380 ) | ( n_n108  &  wire305 ) | ( n_n108  &  _2023 ) ;
 assign _2023 = ( i_9_  &  (~ i_10_)  &  i_11_  &  wire715 ) ;
 assign _2026 = ( n_n162  &  n_n220  &  n_n126  &  wire1205 ) ;
 assign _2056 = ( n_n47  &  wire326 ) | ( n_n47  &  wire327 ) | ( n_n47  &  wire312 ) ;
 assign _2059 = ( n_n46  &  wire303 ) | ( n_n46  &  wire321 ) | ( n_n46  &  wire410 ) ;
 assign _2060 = ( n_n46  &  wire302 ) | ( n_n46  &  wire316 ) | ( n_n46  &  _2071 ) ;
 assign _2071 = ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire721 ) ;
 assign _2123 = ( n_n40  &  wire380 ) | ( n_n40  &  wire352 ) | ( n_n40  &  _2126 ) ;
 assign _2126 = ( i_9_  &  (~ i_10_)  &  i_11_  &  wire715 ) ;
 assign _2182 = ( n_n218  &  n_n35  &  n_n220  &  wire911 ) ;
 assign _2199 = ( n_n218  &  wire714  &  wire840  &  _29212 ) ;
 assign _2250 = ( wire721  &  n_n199  &  wire190 ) ;
 assign _2264 = ( n_n40  &  wire260 ) | ( n_n40  &  wire373 ) | ( n_n40  &  _2265 ) ;
 assign _2265 = ( i_9_  &  i_10_  &  i_11_  &  wire721 ) ;
 assign _2270 = ( n_n212  &  wire302 ) | ( n_n212  &  wire316 ) | ( n_n212  &  _31883 ) ;
 assign _2332 = ( n_n212  &  wire292 ) | ( n_n212  &  wire311 ) | ( n_n212  &  wire317 ) ;
 assign _2335 = ( n_n197  &  wire316 ) | ( n_n197  &  wire331 ) | ( n_n197  &  wire312 ) ;
 assign _2519 = ( wire725  &  n_n41  &  _29611 ) ;
 assign _2561 = ( n_n162  &  wire714  &  wire865  &  _29429 ) ;
 assign _2581 = ( n_n31  &  wire324 ) | ( n_n31  &  wire94 ) | ( n_n31  &  wire104 ) ;
 assign _2591 = ( n_n31  &  wire59 ) | ( n_n31  &  wire289 ) | ( n_n31  &  _2594 ) ;
 assign _2594 = ( (~ i_9_)  &  (~ i_10_)  &  i_11_  &  wire729 ) ;
 assign _2597 = ( n_n31  &  wire117 ) | ( n_n31  &  wire281 ) | ( n_n31  &  wire294 ) ;
 assign _2661 = ( wire730  &  wire1229  &  _31512 ) ;
 assign _2679 = ( n_n48  &  wire714  &  wire122  &  _29131 ) ;
 assign _2726 = ( n_n108  &  wire51 ) | ( n_n108  &  wire210 ) | ( n_n108  &  _2729 ) ;
 assign _2729 = ( (~ i_9_)  &  (~ i_10_)  &  (~ i_11_)  &  wire720 ) ;
 assign _2737 = ( n_n101  &  wire256 ) | ( n_n101  &  wire222 ) | ( n_n101  &  _2740 ) ;
 assign _2738 = ( n_n101  &  wire150 ) | ( n_n101  &  _31455 ) ;
 assign _2740 = ( (~ i_9_)  &  (~ i_10_)  &  i_11_  &  wire719 ) ;
 assign _2752 = ( n_n108  &  wire78 ) | ( n_n108  &  wire252 ) | ( n_n108  &  wire18646 ) ;
 assign _2775 = ( n_n108  &  wire155 ) | ( n_n108  &  wire215 ) | ( n_n108  &  _2778 ) ;
 assign _2778 = ( i_9_  &  i_10_  &  (~ i_11_)  &  wire720 ) ;
 assign _2781 = ( n_n108  &  wire100 ) | ( n_n108  &  wire272 ) | ( n_n108  &  _2784 ) ;
 assign _2784 = ( i_9_  &  (~ i_10_)  &  i_11_  &  wire720 ) ;
 assign _2787 = ( n_n162  &  n_n220  &  n_n126  &  wire250 ) ;
 assign _2858 = ( n_n218  &  n_n124  &  n_n220  &  wire74 ) ;
 assign _2863 = ( wire168  &  n_n125 ) | ( n_n125  &  wire74 ) | ( n_n125  &  wire68 ) ;
 assign _2866 = ( wire143  &  n_n125 ) | ( wire47  &  n_n125 ) | ( n_n125  &  wire151 ) ;
 assign _2884 = ( wire176  &  n_n123 ) | ( n_n123  &  wire153 ) | ( n_n123  &  wire18537 ) ;
 assign _2890 = ( n_n218  &  n_n220  &  n_n126  &  wire960 ) ;
 assign _2894 = ( n_n218  &  n_n220  &  n_n126  &  wire1730 ) ;
 assign _2901 = ( n_n218  &  n_n124  &  n_n220  &  wire52 ) ;
 assign _2906 = ( wire137  &  n_n123 ) | ( wire131  &  n_n123 ) | ( wire55  &  n_n123 ) ;
 assign _2909 = ( wire137  &  n_n125 ) | ( wire131  &  n_n125 ) | ( n_n125  &  wire130 ) ;
 assign _2912 = ( n_n218  &  n_n220  &  n_n126  &  wire147 ) ;
 assign _2919 = ( wire132  &  n_n123 ) | ( wire149  &  n_n123 ) | ( wire126  &  n_n123 ) ;
 assign _2938 = ( wire877  &  _31297 ) | ( wire877  &  _31298 ) ;
 assign _2970 = ( n_n40  &  wire130 ) | ( n_n40  &  wire139 ) | ( n_n40  &  wire128 ) ;
 assign _2973 = ( wire132  &  n_n40 ) | ( n_n40  &  wire126 ) | ( n_n40  &  wire52 ) ;
 assign _2976 = ( wire137  &  n_n40 ) | ( wire131  &  n_n40 ) | ( n_n40  &  wire149 ) ;
 assign _2981 = ( wire152  &  n_n46 ) | ( wire122  &  n_n46 ) | ( n_n46  &  _31251 ) ;
 assign _2990 = ( wire143  &  n_n40 ) | ( wire47  &  n_n40 ) | ( n_n40  &  _2993 ) ;
 assign _2993 = ( i_9_  &  i_10_  &  i_11_  &  wire724 ) ;
 assign _3004 = ( n_n41  &  wire55 ) | ( n_n41  &  wire156 ) | ( n_n41  &  _3007 ) ;
 assign _3007 = ( i_9_  &  i_10_  &  (~ i_11_)  &  wire724 ) ;
 assign _3035 = ( n_n47  &  wire93 ) | ( n_n47  &  wire273 ) | ( n_n47  &  wire54 ) ;
 assign _3077 = ( n_n46  &  wire198 ) | ( n_n46  &  wire212 ) | ( n_n46  &  wire18388 ) ;
 assign _3082 = ( n_n46  &  wire115 ) | ( n_n46  &  wire221 ) | ( n_n46  &  wire298 ) ;
 assign _3089 = ( n_n47  &  wire324 ) | ( n_n47  &  wire94 ) | ( n_n47  &  _3092 ) ;
 assign _3092 = ( (~ i_9_)  &  (~ i_10_)  &  (~ i_11_)  &  wire729 ) ;
 assign _3095 = ( n_n47  &  wire117 ) | ( n_n47  &  wire294 ) | ( n_n47  &  _3098 ) ;
 assign _3098 = ( i_9_  &  (~ i_10_)  &  i_11_  &  wire729 ) ;
 assign _3109 = ( n_n46  &  wire118 ) | ( n_n46  &  wire324 ) | ( n_n46  &  _3112 ) ;
 assign _3110 = ( n_n46  &  wire120 ) | ( n_n46  &  wire179 ) ;
 assign _3112 = ( i_9_  &  (~ i_10_)  &  i_11_  &  wire729 ) ;
 assign _3127 = ( n_n2  &  _31166 ) | ( n_n2  &  _31167 ) ;
 assign _3149 = ( wire130  &  n_n113 ) | ( wire139  &  n_n113 ) | ( n_n113  &  wire18334 ) ;
 assign _3158 = ( wire720  &  n_n191  &  n_n42 ) ;
 assign _3273 = ( n_n48  &  n_n220  &  n_n200  &  wire182 ) ;
 assign _3304 = ( n_n40  &  wire268 ) | ( n_n40  &  wire54 ) | ( n_n40  &  wire399 ) ;
 assign _3312 = ( n_n40  &  wire111 ) | ( n_n40  &  wire206 ) | ( n_n40  &  wire368 ) ;
 assign _3332 = ( n_n40  &  wire93 ) | ( n_n40  &  wire273 ) | ( n_n40  &  _3335 ) ;
 assign _3335 = ( (~ i_9_)  &  (~ i_10_)  &  (~ i_11_)  &  wire729 ) ;
 assign _3344 = ( wire729  &  n_n40  &  _29904 ) ;
 assign _3392 = ( n_n41  &  wire118 ) | ( n_n41  &  wire298 ) | ( n_n41  &  wire18278 ) ;
 assign _3429 = ( n_n47  &  wire186 ) | ( n_n47  &  wire209 ) | ( n_n47  &  wire174 ) ;
 assign _3430 = ( n_n47  &  wire217 ) | ( n_n47  &  wire18196 ) ;
 assign _3440 = ( n_n177  &  wire719  &  n_n46 ) ;
 assign _3486 = ( n_n48  &  wire714  &  wire130  &  _29234 ) ;
 assign _3568 = ( n_n36  &  wire153 ) | ( n_n36  &  wire135 ) | ( n_n36  &  _30848 ) ;
 assign _3637 = ( wire157  &  n_n212 ) | ( n_n212  &  wire204 ) | ( n_n212  &  _30792 ) ;
 assign _3638 = ( n_n212  &  wire80 ) | ( n_n212  &  wire78 ) | ( n_n212  &  _30794 ) ;
 assign _3639 = ( n_n212  &  wire150 ) | ( n_n212  &  wire217 ) ;
 assign _3809 = ( n_n47  &  _30656 ) | ( n_n47  &  _30657 ) ;
 assign _3810 = ( n_n47  &  wire78 ) | ( n_n47  &  wire217 ) | ( n_n47  &  _3812 ) ;
 assign _3811 = ( n_n47  &  wire150 ) | ( n_n47  &  _30659 ) ;
 assign _3812 = ( (~ i_9_)  &  (~ i_10_)  &  i_11_  &  wire719 ) ;
 assign _3827 = ( n_n47  &  wire153 ) | ( n_n47  &  wire135 ) | ( n_n47  &  _30650 ) ;
 assign _3899 = ( n_n218  &  wire714  &  wire130  &  _29212 ) ;
 assign _3948 = ( i_7_  &  i_6_  &  n_n159  &  _30571 ) ;
 assign _4048 = ( wire93  &  n_n112 ) | ( n_n112  &  wire171 ) | ( n_n112  &  wire17721 ) ;
 assign _4072 = ( n_n162  &  n_n35  &  n_n220  &  wire157 ) ;
 assign _4088 = ( n_n101  &  wire156 ) | ( n_n101  &  wire176 ) | ( n_n101  &  wire212 ) ;
 assign _4188 = ( n_n218  &  n_n220  &  n_n126  &  wire100 ) ;
 assign _4253 = ( n_n48  &  n_n220  &  n_n200  &  wire172 ) ;
 assign _4363 = ( n_n4  &  _30322 ) | ( n_n4  &  _30323 ) ;
 assign _4473 = ( n_n30  &  wire127 ) | ( n_n30  &  wire158 ) | ( n_n30  &  wire134 ) ;
 assign _4479 = ( n_n162  &  wire714  &  wire125  &  _29429 ) ;
 assign _4492 = ( wire152  &  n_n33 ) | ( n_n33  &  wire220 ) | ( n_n33  &  _4495 ) ;
 assign _4495 = ( (~ i_9_)  &  i_10_  &  (~ i_11_)  &  wire720 ) ;
 assign _4527 = ( n_n218  &  wire714  &  wire158  &  _29276 ) ;
 assign _4585 = ( wire234  &  n_n123 ) | ( wire84  &  n_n123 ) | ( n_n123  &  wire220 ) ;
 assign _4657 = ( n_n48  &  n_n220  &  n_n200  &  wire1173 ) ;
 assign _4707 = ( n_n46  &  wire155 ) | ( n_n46  &  wire60 ) | ( n_n46  &  wire220 ) ;
 assign _4718 = ( n_n48  &  wire714  &  wire85  &  _29234 ) ;
 assign _4739 = ( n_n162  &  n_n220  &  n_n126  &  wire220 ) ;
 assign _4740 = ( n_n162  &  n_n220  &  n_n126  &  wire84 ) ;
 assign _4890 = ( n_n41  &  wire229 ) | ( n_n41  &  wire265 ) | ( n_n41  &  _29934 ) ;
 assign _4924 = ( n_n40  &  wire70 ) | ( n_n40  &  wire374 ) | ( n_n40  &  _29913 ) ;
 assign _4944 = ( n_n34  &  wire120 ) | ( n_n34  &  wire117 ) | ( n_n34  &  _29895 ) ;
 assign _4984 = ( n_n34  &  wire116 ) | ( n_n34  &  wire371 ) | ( n_n34  &  _4987 ) ;
 assign _4987 = ( (~ i_9_)  &  i_10_  &  i_11_  &  wire725 ) ;
 assign _4992 = ( wire725  &  wire226  &  _29849 ) | ( wire725  &  wire226  &  _29851 ) ;
 assign _5193 = ( n_n47  &  wire158 ) | ( n_n47  &  wire299 ) | ( n_n47  &  _29659 ) ;
 assign _5201 = ( wire158  &  n_n46 ) | ( n_n46  &  wire299 ) | ( n_n46  &  _5204 ) ;
 assign _5204 = ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire725 ) ;
 assign _5207 = ( n_n101  &  wire60 ) | ( n_n101  &  wire377 ) | ( n_n101  &  _29643 ) ;
 assign _5208 = ( n_n108  &  wire60 ) | ( n_n108  &  wire351 ) | ( n_n108  &  _29645 ) ;
 assign _5289 = ( n_n30  &  wire176 ) | ( n_n30  &  wire299 ) | ( n_n30  &  wire418 ) ;
 assign _5329 = ( n_n218  &  n_n35  &  n_n220  &  wire1056 ) ;
 assign _5528 = ( n_n46  &  wire85 ) | ( n_n46  &  _29379 ) ;
 assign _5529 = ( n_n46  &  wire219 ) | ( n_n46  &  wire108 ) | ( n_n46  &  wire258 ) ;
 assign _5561 = ( wire720  &  n_n46  &  n_n199 ) ;
 assign _5601 = ( n_n123  &  wire69 ) | ( n_n123  &  wire208 ) | ( n_n123  &  wire148 ) ;
 assign _5628 = ( n_n197  &  wire150 ) | ( n_n197  &  wire78 ) | ( n_n197  &  _29313 ) ;
 assign _5825 = ( wire719  &  n_n41  &  _29189 ) ;
 assign _5873 = ( n_n48  &  n_n220  &  n_n200  &  wire1789 ) ;
 assign _5959 = ( wire1041  &  _29052 ) | ( wire1041  &  _29053 ) ;
 assign _5996 = ( i_5_  &  (~ i_3_)  &  (~ i_4_)  &  wire736 ) ;
 assign _28911 = ( (~ i_9_)  &  (~ i_10_)  &  (~ i_11_) ) ;
 assign _28939 = ( wire5057 ) | ( wire16872 ) | ( wire463 ) | ( wire16863 ) ;
 assign _29017 = ( wire569 ) | ( wire16888 ) ;
 assign _29024 = ( wire16898 ) | ( wire16892 ) | ( wire16896 ) | ( _29017 ) ;
 assign _29028 = ( (~ i_9_)  &  i_10_  &  (~ i_11_) ) ;
 assign _29046 = ( i_9_  &  i_10_  &  (~ i_11_)  &  wire729 ) ;
 assign _29052 = ( n_n162  &  n_n159  &  n_n161 ) | ( n_n159  &  n_n48  &  n_n161 ) ;
 assign _29053 = ( n_n162  &  n_n159  &  n_n124 ) | ( n_n159  &  n_n124  &  n_n48 ) ;
 assign _29117 = ( (~ i_9_)  &  (~ i_10_)  &  i_11_ ) ;
 assign _29131 = ( (~ i_6_)  &  i_7_ ) ;
 assign _29155 = ( i_9_  &  (~ i_10_)  &  i_11_ ) ;
 assign _29156 = ( n_n41  &  wire100 ) | ( wire720  &  n_n41  &  _29155 ) ;
 assign _29181 = ( i_7_  &  (~ i_6_)  &  n_n48  &  wire714 ) ;
 assign _29189 = ( i_9_  &  i_10_  &  i_11_ ) ;
 assign _29191 = ( wire653 ) | ( n_n41  &  wire208 ) | ( n_n41  &  wire148 ) ;
 assign _29192 = ( wire518 ) | ( wire4890 ) | ( wire4891 ) | ( _5825 ) ;
 assign _29193 = ( wire17019 ) | ( wire17018 ) ;
 assign _29197 = ( (~ i_7_)  &  (~ i_6_)  &  n_n218  &  wire714 ) ;
 assign _29204 = ( i_9_  &  (~ i_10_)  &  i_11_  &  wire724 ) ;
 assign _29206 = ( n_n124  &  n_n48  &  n_n220 ) ;
 assign _29207 = ( n_n39  &  _29204 ) | ( wire104  &  _29206 ) ;
 assign _29210 = ( wire17028 ) | ( wire17044 ) | ( wire151  &  _29197 ) ;
 assign _29212 = ( (~ i_6_)  &  (~ i_7_) ) ;
 assign _29222 = ( i_9_  &  (~ i_10_)  &  i_11_ ) ;
 assign _29234 = ( i_6_  &  i_7_ ) ;
 assign _29252 = ( i_9_  &  i_10_  &  i_11_ ) ;
 assign _29269 = ( n_n48  &  n_n220  &  n_n161 ) ;
 assign _29274 = ( wire17050 ) | ( wire17047 ) | ( _29210 ) ;
 assign _29276 = ( (~ i_6_)  &  i_7_ ) ;
 assign _29298 = ( i_9_  &  i_10_  &  i_11_ ) ;
 assign _29305 = ( wire17116 ) | ( wire137  &  n_n197 ) | ( wire146  &  n_n197 ) ;
 assign _29309 = ( (~ i_9_)  &  (~ i_10_)  &  i_11_ ) ;
 assign _29313 = ( n_n177  &  wire719 ) | ( n_n177  &  wire728 ) | ( wire719  &  _29117 ) ;
 assign _29315 = ( n_n125  &  wire86 ) | ( n_n125  &  wire180 ) ;
 assign _29327 = ( n_n218  &  n_n220  &  n_n126 ) ;
 assign _29332 = ( wire4743 ) | ( wire4750 ) | ( wire153  &  _29327 ) ;
 assign _29343 = ( wire17119 ) | ( wire17137 ) | ( _29305 ) | ( _29332 ) ;
 assign _29353 = ( n_n101  &  wire218 ) | ( n_n101  &  wire141 ) ;
 assign _29356 = ( n_n162  &  n_n124  &  n_n220 ) ;
 assign _29375 = ( wire4829 ) | ( wire4831 ) | ( _5561 ) | ( _29353 ) ;
 assign _29379 = ( wire729  &  n_n199 ) | ( n_n199  &  wire726 ) ;
 assign _29381 = ( _5529 ) | ( n_n46  &  wire85 ) | ( n_n46  &  _29379 ) ;
 assign _29383 = ( (~ i_9_)  &  (~ i_10_)  &  i_11_  &  wire720 ) ;
 assign _29386 = ( n_n4900 ) | ( wire4933 ) | ( n_n101  &  _29383 ) ;
 assign _29424 = ( wire17082 ) | ( wire16997 ) | ( _29381 ) | ( _29386 ) ;
 assign _29427 = ( wire17153 ) | ( wire17154 ) | ( wire17156 ) ;
 assign _29429 = ( (~ i_6_)  &  (~ i_7_) ) ;
 assign _29431 = ( n_n31  &  wire137 ) | ( n_n31  &  wire46 ) ;
 assign _29448 = ( wire584 ) | ( wire137  &  n_n34 ) | ( n_n34  &  wire46 ) ;
 assign _29458 = ( n_n34  &  wire125 ) | ( wire725  &  n_n34  &  _29298 ) ;
 assign _29464 = ( wire690 ) | ( n_n31  &  wire149 ) ;
 assign _29471 = ( n_n31  &  wire252 ) | ( wire725  &  n_n31  &  _29309 ) ;
 assign _29472 = ( wire16966 ) | ( n_n31  &  wire80 ) | ( n_n31  &  wire78 ) ;
 assign _29474 = ( wire4953 ) | ( wire16960 ) | ( _29448 ) | ( _29464 ) ;
 assign _29477 = ( wire17166 ) | ( wire17170 ) | ( wire17172 ) | ( _29431 ) ;
 assign _29478 = ( n_n4399 ) | ( n_n4404 ) | ( wire17064 ) | ( _29274 ) ;
 assign _29479 = ( wire17158 ) | ( wire17174 ) | ( _29427 ) | ( _29477 ) ;
 assign _29480 = ( i_7_  &  (~ i_6_)  &  i_3_  &  i_4_ ) ;
 assign _29539 = ( (~ i_9_)  &  i_10_  &  (~ i_11_) ) ;
 assign _29544 = ( wire4649 ) | ( wire17226 ) | ( wire17231 ) | ( _5329 ) ;
 assign _29545 = ( wire4644 ) | ( wire4651 ) | ( wire4655 ) | ( wire17220 ) ;
 assign _29607 = ( n_n2239 ) | ( wire4643 ) | ( _29544 ) | ( _29545 ) ;
 assign _29608 = ( n_n46  &  wire168 ) | ( n_n46  &  wire181 ) ;
 assign _29611 = ( (~ i_9_)  &  i_10_  &  (~ i_11_) ) ;
 assign _29613 = ( i_9_  &  i_10_  &  (~ i_11_) ) ;
 assign _29641 = ( i_9_  &  i_10_  &  (~ i_11_) ) ;
 assign _29643 = ( wire725  &  _29298 ) | ( wire722  &  _29641 ) ;
 assign _29645 = ( wire725  &  _29298 ) | ( wire722  &  _29539 ) ;
 assign _29649 = ( n_n5144 ) | ( wire4685 ) | ( wire17191 ) | ( _29608 ) ;
 assign _29651 = ( n_n46  &  wire308 ) | ( n_n46  &  wire418 ) ;
 assign _29653 = ( n_n48  &  n_n220  &  n_n161 ) ;
 assign _29659 = ( i_9_  &  (~ i_10_)  &  i_11_  &  wire725 ) | ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire725 ) | ( (~ i_9_)  &  (~ i_10_)  &  (~ i_11_)  &  wire725 ) ;
 assign _29694 = ( wire17198 ) | ( _5201 ) | ( _29651 ) ;
 assign _29711 = ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire722 ) ;
 assign _29722 = ( wire4619 ) | ( n_n112  &  wire307 ) | ( n_n112  &  _29711 ) ;
 assign _29731 = ( i_9_  &  i_10_  &  (~ i_11_) ) ;
 assign _29755 = ( (~ i_9_)  &  (~ i_10_)  &  i_11_ ) ;
 assign _29771 = ( wire17256 ) | ( n_n2340 ) | ( wire17268 ) | ( _29722 ) ;
 assign _29772 = ( wire17257 ) | ( wire17275 ) | ( wire17276 ) ;
 assign _29782 = ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  (~ i_15_) ) ;
 assign _29784 = ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  i_15_ ) ;
 assign _29832 = ( wire4561 ) | ( wire4562 ) | ( wire17303 ) ;
 assign _29849 = ( (~ i_9_)  &  (~ i_10_)  &  (~ i_11_) ) ;
 assign _29851 = ( (~ i_9_)  &  (~ i_10_)  &  i_11_ ) ;
 assign _29864 = ( wire4558 ) | ( wire17307 ) | ( wire17314 ) | ( _4992 ) ;
 assign _29870 = ( (~ i_9_)  &  (~ i_10_)  &  (~ i_11_)  &  wire729 ) ;
 assign _29885 = ( i_9_  &  i_10_  &  (~ i_11_)  &  wire729 ) ;
 assign _29886 = ( (~ i_9_)  &  (~ i_10_)  &  i_11_  &  wire729 ) ;
 assign _29890 = ( n_n36  &  _29885 ) | ( n_n34  &  _29886 ) ;
 assign _29895 = ( i_15_  &  n_n211  &  n_n177 ) | ( (~ i_15_)  &  n_n211  &  n_n177 ) | ( i_15_  &  n_n211  &  n_n170 ) | ( (~ i_15_)  &  n_n211  &  n_n170 ) ;
 assign _29896 = ( _4944 ) | ( wire4539 ) ;
 assign _29897 = ( wire17322 ) | ( wire4544 ) | ( n_n36  &  _29870 ) ;
 assign _29898 = ( wire4554 ) | ( wire17325 ) | ( _29864 ) | ( _29896 ) ;
 assign _29899 = ( wire17305 ) | ( _29771 ) | ( _29772 ) | ( _29832 ) ;
 assign _29900 = ( wire17213 ) | ( _29694 ) | ( _29897 ) | ( _29898 ) ;
 assign _29904 = ( i_9_  &  (~ i_10_)  &  (~ i_11_) ) ;
 assign _29913 = ( i_9_  &  i_10_  &  i_11_  &  wire722 ) | ( (~ i_9_)  &  i_10_  &  i_11_  &  wire722 ) ;
 assign _29934 = ( i_9_  &  (~ i_10_)  &  i_11_  &  wire722 ) | ( (~ i_9_)  &  (~ i_10_)  &  i_11_  &  wire722 ) ;
 assign _29936 = ( wire397 ) | ( wire4510 ) | ( wire4523 ) | ( wire17337 ) ;
 assign _29938 = ( wire17341 ) | ( wire17342 ) | ( _4890 ) | ( _29936 ) ;
 assign _29962 = ( (~ i_9_)  &  i_10_  &  (~ i_11_)  &  wire722 ) ;
 assign _29963 = ( n_n101  &  wire351 ) | ( n_n101  &  wire57 ) | ( n_n101  &  _29962 ) ;
 assign _30001 = ( wire158  &  n_n197 ) | ( wire158  &  n_n212 ) ;
 assign _30030 = ( n_n2249 ) | ( wire17364 ) | ( wire17365 ) | ( _29938 ) ;
 assign _30031 = ( wire17249 ) | ( wire17193 ) | ( _29607 ) | ( _29649 ) ;
 assign _30032 = ( _29899 ) | ( _29900 ) | ( _30031 ) ;
 assign _30036 = ( n_n162  &  n_n220  &  n_n126 ) ;
 assign _30037 = ( wire1862  &  _29356 ) | ( wire141  &  _30036 ) ;
 assign _30039 = ( wire17470 ) | ( n_n101  &  wire205 ) | ( n_n101  &  wire204 ) ;
 assign _30040 = ( wire17471 ) | ( wire4839 ) | ( wire17469 ) | ( _30037 ) ;
 assign _30042 = ( i_9_  &  i_10_  &  (~ i_11_) ) ;
 assign _30050 = ( n_n162  &  n_n220  &  n_n126 ) ;
 assign _30071 = ( wire4829 ) | ( wire720  &  n_n46  &  n_n199 ) ;
 assign _30073 = ( wire17479 ) | ( wire511 ) | ( _4739 ) | ( _4740 ) ;
 assign _30076 = ( n_n46  &  wire205 ) | ( n_n46  &  wire215 ) ;
 assign _30081 = ( i_7_  &  i_6_  &  n_n48  &  wire714 ) ;
 assign _30087 = ( _4707 ) | ( _30076 ) | ( wire800  &  _30081 ) ;
 assign _30101 = ( n_n4904 ) | ( wire544 ) | ( wire4323 ) | ( wire4324 ) ;
 assign _30102 = ( wire17082 ) | ( wire17501 ) | ( _5528 ) | ( _5529 ) ;
 assign _30108 = ( n_n41  &  wire155 ) | ( n_n41  &  wire205 ) ;
 assign _30113 = ( n_n41  &  wire60 ) | ( n_n41  &  wire220 ) ;
 assign _30119 = ( wire4286 ) | ( wire4904 ) | ( wire153  &  _29181 ) ;
 assign _30120 = ( wire17534 ) | ( wire4291 ) | ( _30113 ) ;
 assign _30153 = ( i_9_  &  i_10_  &  (~ i_11_)  &  wire725 ) ;
 assign _30155 = ( (~ i_9_)  &  i_10_  &  (~ i_11_) ) ;
 assign _30162 = ( wire549 ) | ( wire4919 ) | ( wire17003 ) | ( wire17562 ) ;
 assign _30163 = ( n_n4460 ) | ( wire17033 ) | ( wire17553 ) | ( wire17550 ) ;
 assign _30166 = ( wire215  &  n_n123 ) | ( wire720  &  n_n123  &  _30042 ) ;
 assign _30172 = ( wire4382 ) | ( wire17459 ) | ( _4585 ) | ( _30166 ) ;
 assign _30175 = ( i_9_  &  i_10_  &  i_11_  &  wire719 ) ;
 assign _30176 = ( wire153  &  _29327 ) | ( n_n125  &  _30175 ) ;
 assign _30194 = ( n_n218  &  n_n220  &  n_n200 ) ;
 assign _30195 = ( wire17575 ) | ( wire123  &  _30194 ) ;
 assign _30198 = ( n_n197  &  wire125 ) | ( wire725  &  n_n197  &  _29298 ) ;
 assign _30203 = ( wire538 ) | ( wire4233 ) | ( _29315 ) | ( _30198 ) ;
 assign _30206 = ( wire17462 ) | ( wire17467 ) | ( _30172 ) ;
 assign _30217 = ( (~ i_7_)  &  (~ i_6_)  &  n_n162  &  wire714 ) ;
 assign _30218 = ( n_n4240 ) | ( wire144  &  _30217 ) ;
 assign _30221 = ( (~ i_7_)  &  (~ i_6_)  &  n_n162  &  wire714 ) ;
 assign _30224 = ( n_n30  &  wire133 ) | ( n_n30  &  wire156 ) ;
 assign _30229 = ( wire4429 ) | ( wire158  &  _30221 ) ;
 assign _30240 = ( n_n34  &  wire55 ) | ( n_n34  &  wire158 ) ;
 assign _30242 = ( n_n36  &  wire133 ) | ( n_n36  &  wire125 ) ;
 assign _30244 = ( wire541 ) | ( wire17441 ) | ( _30240 ) | ( _30242 ) ;
 assign _30248 = ( n_n4106 ) | ( n_n5144 ) ;
 assign _30250 = ( wire17581 ) | ( wire17585 ) | ( _30206 ) | ( _30248 ) ;
 assign _30273 = ( n_n7267 ) | ( wire684 ) | ( wire17596 ) ;
 assign _30296 = ( n_n5144 ) | ( n_n2956 ) | ( _30273 ) ;
 assign _30322 = ( (~ i_9_)  &  i_10_  &  (~ i_11_)  &  wire729 ) | ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire729 ) ;
 assign _30323 = ( n_n156  &  wire730 ) | ( n_n156  &  wire717 ) | ( wire730  &  n_n191 ) | ( wire717  &  n_n191 ) ;
 assign _30347 = ( i_9_  &  (~ i_10_)  &  (~ i_11_) ) ;
 assign _30353 = ( i_7_  &  (~ i_6_)  &  n_n48  &  wire714 ) ;
 assign _30358 = ( n_n41  &  wire142 ) | ( n_n41  &  wire180 ) ;
 assign _30359 = ( wire4130 ) | ( wire85  &  _30353 ) ;
 assign _30362 = ( i_7_  &  (~ i_6_)  &  n_n48  &  wire714 ) ;
 assign _30371 = ( i_9_  &  (~ i_10_)  &  (~ i_11_) ) ;
 assign _30385 = ( n_n48  &  n_n220  &  n_n126 ) ;
 assign _30386 = ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire719 ) ;
 assign _30390 = ( wire157  &  n_n40 ) | ( wire725  &  n_n40  &  _29613 ) ;
 assign _30391 = ( wire17662 ) | ( n_n40  &  wire80 ) | ( n_n40  &  wire78 ) ;
 assign _30395 = ( n_n38  &  wire248 ) | ( n_n39  &  wire248 ) ;
 assign _30401 = ( n_n40  &  wire155 ) | ( n_n40  &  wire205 ) ;
 assign _30404 = ( wire17668 ) | ( wire17674 ) | ( _30395 ) | ( _30401 ) ;
 assign _30450 = ( n_n212  &  wire176 ) | ( wire725  &  n_n212  &  _29298 ) ;
 assign _30453 = ( wire689 ) | ( wire4020 ) | ( wire4027 ) | ( _30450 ) ;
 assign _30455 = ( wire17744 ) | ( wire17746 ) | ( wire17764 ) | ( _4188 ) ;
 assign _30457 = ( wire17695 ) | ( wire17696 ) | ( wire17778 ) ;
 assign _30468 = ( wire17831 ) | ( wire17832 ) | ( wire17836 ) ;
 assign _30471 = ( wire725  &  n_n156 ) | ( n_n156  &  wire721 ) ;
 assign _30482 = ( n_n101  &  wire134 ) | ( n_n101  &  wire123 ) ;
 assign _30484 = ( n_n3570 ) | ( wire4185 ) | ( _4088 ) | ( _30482 ) ;
 assign _30488 = ( (~ i_7_)  &  (~ i_6_)  &  n_n162  &  wire714 ) ;
 assign _30490 = ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire719 ) ;
 assign _30491 = ( wire172  &  _30488 ) | ( n_n31  &  _30490 ) ;
 assign _30495 = ( wire3990 ) | ( wire17783 ) | ( wire17840 ) | ( _4072 ) ;
 assign _30497 = ( wire17626 ) | ( wire17627 ) | ( wire17786 ) | ( _30495 ) ;
 assign _30546 = ( n_n34  &  wire156 ) | ( n_n34  &  wire176 ) ;
 assign _30549 = ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire719 ) ;
 assign _30553 = ( n_n33  &  wire187 ) | ( wire720  &  n_n33  &  _30371 ) ;
 assign _30557 = ( wire3957 ) | ( wire17801 ) | ( _30546 ) | ( _30553 ) ;
 assign _30561 = ( wire17839 ) | ( wire17629 ) | ( _30468 ) | ( _30497 ) ;
 assign _30565 = ( (~ i_6_)  &  i_7_ ) ;
 assign _30568 = ( (~ i_1_)  &  i_2_  &  i_0_ ) ;
 assign _30569 = ( i_6_  &  i_7_ ) ;
 assign _30571 = ( i_5_  &  i_3_  &  i_4_ ) ;
 assign _30578 = ( wire462 ) | ( n_n19  &  wire817  &  _30565 ) ;
 assign _30595 = ( i_5_  &  i_3_  &  i_4_ ) ;
 assign _30599 = ( n_n5144 ) | ( wire3886 ) | ( wire17858 ) | ( _30578 ) ;
 assign _30604 = ( wire146  &  n_n34 ) | ( wire131  &  n_n34 ) ;
 assign _30607 = ( wire640 ) | ( wire17864 ) | ( _3899 ) | ( _30604 ) ;
 assign _30622 = ( n_n218  &  n_n35  &  n_n220 ) ;
 assign _30623 = ( wire151  &  _29197 ) | ( wire181  &  _30622 ) ;
 assign _30650 = ( wire725  &  _29298 ) | ( wire719  &  _30347 ) ;
 assign _30652 = ( n_n47  &  wire176 ) | ( n_n47  &  wire123 ) ;
 assign _30656 = ( i_9_  &  i_10_  &  (~ i_11_)  &  wire725 ) | ( (~ i_9_)  &  (~ i_10_)  &  (~ i_11_)  &  wire725 ) ;
 assign _30657 = ( n_n177  &  wire719 ) | ( wire719  &  n_n149 ) | ( n_n177  &  wire728 ) | ( n_n149  &  wire728 ) ;
 assign _30659 = ( wire725  &  n_n149 ) | ( n_n149  &  wire721 ) ;
 assign _30665 = ( wire17976 ) | ( wire157  &  n_n47 ) | ( n_n47  &  wire172 ) ;
 assign _30668 = ( n_n3555 ) | ( wire18136 ) | ( _3827 ) | ( _30652 ) ;
 assign _30673 = ( i_9_  &  (~ i_10_)  &  i_11_ ) ;
 assign _30694 = ( i_9_  &  i_10_  &  (~ i_11_)  &  wire726 ) ;
 assign _30702 = ( n_n39  &  wire279 ) | ( n_n39  &  wire724  &  _29222 ) ;
 assign _30703 = ( wire18003 ) | ( n_n39  &  wire110 ) | ( n_n39  &  _30694 ) ;
 assign _30710 = ( n_n41  &  wire234 ) | ( n_n41  &  wire84 ) ;
 assign _30763 = ( n_n177  &  wire719 ) | ( wire719  &  n_n149 ) | ( n_n177  &  wire728 ) | ( n_n149  &  wire728 ) ;
 assign _30765 = ( wire725  &  n_n177 ) | ( n_n177  &  wire721 ) | ( wire725  &  n_n199 ) | ( wire721  &  n_n199 ) ;
 assign _30792 = ( wire725  &  n_n149 ) | ( n_n149  &  wire721 ) | ( wire725  &  _29613 ) ;
 assign _30794 = ( wire725  &  _28911 ) | ( wire719  &  _29117 ) ;
 assign _30798 = ( n_n212  &  wire176 ) | ( n_n212  &  wire125 ) ;
 assign _30799 = ( wire18085 ) | ( wire18089 ) | ( _30798 ) ;
 assign _30811 = ( n_n125  &  wire211 ) | ( n_n125  &  wire272 ) ;
 assign _30816 = ( n_n125  &  wire51 ) | ( n_n125  &  wire100 ) ;
 assign _30817 = ( wire18106 ) | ( _30811 ) | ( n_n125  &  wire18111 ) ;
 assign _30819 = ( wire479 ) | ( wire698 ) | ( wire3653 ) | ( wire18096 ) ;
 assign _30821 = ( wire18097 ) | ( wire18120 ) | ( wire18134 ) | ( _30819 ) ;
 assign _30824 = ( wire143  &  n_n36 ) | ( n_n36  &  wire181 ) ;
 assign _30833 = ( wire725  &  _28911 ) | ( wire719  &  _29117 ) ;
 assign _30839 = ( n_n5144 ) | ( n_n31  &  wire172 ) | ( n_n31  &  wire125 ) ;
 assign _30848 = ( wire725  &  _29298 ) | ( wire719  &  _30347 ) ;
 assign _30850 = ( n_n36  &  wire176 ) | ( n_n36  &  wire123 ) ;
 assign _30851 = ( n_n36  &  wire55 ) | ( n_n36  &  wire125 ) ;
 assign _30861 = ( n_n177  &  wire719 ) | ( wire719  &  n_n149 ) | ( n_n177  &  wire728 ) | ( n_n149  &  wire728 ) ;
 assign _30865 = ( n_n2642 ) | ( _3568 ) | ( _30850 ) | ( _30851 ) ;
 assign _30866 = ( n_n3470 ) | ( wire3810 ) | ( wire3811 ) | ( _30865 ) ;
 assign _30869 = ( wire18141 ) | ( wire18142 ) | ( wire18148 ) ;
 assign _30896 = ( i_5_  &  (~ i_3_)  &  (~ i_4_) ) ;
 assign _30923 = ( wire55  &  n_n46 ) | ( wire127  &  n_n46 ) ;
 assign _30926 = ( wire674 ) | ( wire671 ) | ( _3486 ) | ( _30923 ) ;
 assign _30948 = ( wire651 ) | ( wire3575 ) | ( wire18190 ) | ( _3440 ) ;
 assign _30950 = ( wire18193 ) | ( wire18201 ) | ( wire18205 ) | ( _30948 ) ;
 assign _30958 = ( wire18220 ) | ( wire18221 ) | ( wire18222 ) ;
 assign _30959 = ( wire18212 ) | ( n_n3085 ) | ( _30958 ) ;
 assign _30964 = ( (~ i_9_)  &  (~ i_10_)  &  (~ i_11_)  &  wire725 ) ;
 assign _30973 = ( n_n41  &  wire198 ) | ( n_n41  &  wire221 ) ;
 assign _30974 = ( i_9_  &  i_10_  &  (~ i_11_)  &  wire726 ) ;
 assign _30980 = ( i_7_  &  (~ i_6_)  &  n_n48  &  wire714 ) ;
 assign _30983 = ( i_7_  &  (~ i_6_)  &  n_n48  &  wire714 ) ;
 assign _30984 = ( wire115  &  _30980 ) | ( wire212  &  _30983 ) ;
 assign _30987 = ( n_n5075 ) | ( n_n5070 ) | ( wire3471 ) ;
 assign _30988 = ( wire18283 ) | ( _3392 ) | ( _30973 ) ;
 assign _31018 = ( n_n40  &  wire341 ) | ( n_n40  &  wire243 ) ;
 assign _31021 = ( n_n40  &  wire184 ) | ( n_n40  &  wire162 ) ;
 assign _31022 = ( i_9_  &  i_10_  &  i_11_  &  wire726 ) ;
 assign _31026 = ( _3304 ) | ( _3312 ) | ( _31018 ) | ( _31021 ) ;
 assign _31044 = ( n_n5144 ) | ( wire18232 ) | ( _31026 ) ;
 assign _31045 = ( wire3524 ) | ( wire18266 ) | ( wire18268 ) | ( _3344 ) ;
 assign _31049 = ( i_7_  &  (~ i_6_)  &  n_n48  &  wire714 ) ;
 assign _31050 = ( (~ i_9_)  &  i_10_  &  (~ i_11_)  &  wire725 ) ;
 assign _31059 = ( wire18214 ) | ( wire18297 ) | ( n_n3033 ) | ( _30950 ) ;
 assign _31078 = ( i_7_  &  (~ i_6_)  &  n_n162  &  wire714 ) ;
 assign _31080 = ( (~ i_9_)  &  (~ i_10_)  &  (~ i_11_)  &  wire721 ) ;
 assign _31081 = ( (~ i_9_)  &  i_10_  &  (~ i_11_)  &  wire728 ) ;
 assign _31082 = ( wire1417  &  _31078 ) | ( n_n32  &  _31080 ) ;
 assign _31115 = ( (~ i_9_)  &  i_10_  &  (~ i_11_)  &  wire725 ) ;
 assign _31116 = ( wire185  &  n_n14 ) | ( wire270  &  n_n14 ) ;
 assign _31117 = ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire720 ) ;
 assign _31127 = ( wire3403 ) | ( wire18342 ) | ( n_n43  &  _31117 ) ;
 assign _31128 = ( (~ i_9_)  &  (~ i_10_)  &  (~ i_11_)  &  wire725 ) ;
 assign _31132 = ( n_n1566 ) | ( n_n42  &  wire217 ) | ( n_n42  &  _31128 ) ;
 assign _31135 = ( n_n218  &  n_n220  &  n_n161 ) ;
 assign _31139 = ( n_n113  &  wire124 ) | ( n_n113  &  wire128 ) ;
 assign _31143 = ( wire3409 ) | ( wire63  &  _31135 ) ;
 assign _31145 = ( n_n5144 ) | ( wire18345 ) | ( _31127 ) ;
 assign _31151 = ( i_7_  &  i_6_  &  n_n218  &  n_n19 ) | ( (~ i_7_)  &  i_6_  &  n_n218  &  n_n19 ) | ( i_7_  &  (~ i_6_)  &  n_n218  &  n_n19 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n218  &  n_n19 ) ;
 assign _31153 = ( i_5_  &  i_3_  &  i_4_ ) ;
 assign _31166 = ( i_9_  &  i_10_  &  (~ i_11_)  &  wire717 ) | ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire717 ) ;
 assign _31167 = ( wire729  &  n_n156 ) | ( n_n156  &  wire730 ) | ( wire729  &  n_n191 ) | ( wire730  &  n_n191 ) ;
 assign _31173 = ( n_n159  &  n_n48  &  n_n161 ) ;
 assign _31175 = ( wire3374 ) | ( wire3375 ) | ( wire185  &  _31173 ) ;
 assign _31176 = ( wire18375 ) | ( wire18372 ) | ( wire270  &  n_n14 ) ;
 assign _31182 = ( i_7_  &  i_6_  &  n_n48  &  wire714 ) ;
 assign _31186 = ( n_n47  &  wire53 ) | ( n_n46  &  wire53 ) | ( n_n46  &  wire294 ) ;
 assign _31188 = ( n_n47  &  wire120 ) | ( n_n47  &  wire281 ) ;
 assign _31190 = ( n_n47  &  wire179 ) | ( n_n47  &  wire184 ) ;
 assign _31193 = ( _3089 ) | ( _3095 ) | ( _31188 ) | ( _31190 ) ;
 assign _31195 = ( wire18429 ) | ( wire18433 ) | ( wire1576  &  _31182 ) ;
 assign _31197 = ( n_n46  &  wire59 ) | ( n_n46  &  wire289 ) ;
 assign _31199 = ( n_n46  &  wire247 ) | ( n_n46  &  wire116 ) ;
 assign _31203 = ( _3077 ) | ( _3082 ) | ( _31197 ) | ( _31199 ) ;
 assign _31214 = ( wire3325 ) | ( n_n47  &  wire98 ) ;
 assign _31216 = ( n_n47  &  wire241 ) | ( n_n47  &  wire268 ) ;
 assign _31219 = ( n_n46  &  wire74 ) | ( n_n46  &  wire68 ) ;
 assign _31221 = ( wire577 ) | ( _3035 ) | ( _31216 ) | ( _31219 ) ;
 assign _31223 = ( wire18393 ) | ( wire18420 ) | ( _31203 ) | ( _31214 ) ;
 assign _31229 = ( n_n5319 ) | ( wire212  &  _30983 ) ;
 assign _31237 = ( wire363 ) | ( n_n40  &  wire1383 ) ;
 assign _31238 = ( n_n5070 ) | ( wire18461 ) | ( wire3279 ) | ( wire3280 ) ;
 assign _31243 = ( wire359 ) | ( n_n40  &  wire1386 ) ;
 assign _31251 = ( n_n156  &  wire719 ) | ( n_n156  &  wire728 ) | ( wire719  &  _30155 ) ;
 assign _31262 = ( i_7_  &  (~ i_6_)  &  n_n48  &  wire714 ) ;
 assign _31264 = ( wire146  &  n_n40 ) | ( n_n40  &  wire46 ) ;
 assign _31266 = ( n_n40  &  wire147 ) | ( n_n40  &  wire129 ) ;
 assign _31270 = ( i_7_  &  (~ i_6_)  &  n_n48  &  wire714 ) ;
 assign _31272 = ( n_n40  &  wire63 ) | ( n_n40  &  wire48 ) ;
 assign _31276 = ( _2973 ) | ( _31266 ) | ( wire1520  &  _31270 ) ;
 assign _31278 = ( n_n5144 ) | ( wire1381  &  _31262 ) ;
 assign _31279 = ( _2976 ) | ( _31264 ) | ( _31278 ) ;
 assign _31280 = ( wire3258 ) | ( wire18487 ) | ( _31243 ) ;
 assign _31283 = ( n_n3166 ) | ( wire18437 ) | ( wire18434 ) | ( _31195 ) ;
 assign _31285 = ( (~ i_9_)  &  i_10_  &  (~ i_11_)  &  wire729 ) | ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire729 ) ;
 assign _31286 = ( n_n5  &  wire87 ) | ( n_n6  &  wire87 ) | ( n_n5  &  _31285 ) | ( n_n6  &  _31285 ) ;
 assign _31297 = ( (~ i_9_)  &  i_10_  &  (~ i_11_)  &  wire729 ) | ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire729 ) ;
 assign _31298 = ( wire730  &  n_n149 ) | ( wire717  &  n_n149 ) | ( wire730  &  n_n191 ) | ( wire717  &  n_n191 ) ;
 assign _31302 = ( i_7_  &  i_6_  &  n_n218  &  n_n19 ) | ( (~ i_7_)  &  i_6_  &  n_n218  &  n_n19 ) | ( i_7_  &  (~ i_6_)  &  n_n218  &  n_n19 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n218  &  n_n19 ) ;
 assign _31305 = ( (~ i_1_)  &  (~ i_2_)  &  i_0_ ) ;
 assign _31318 = ( i_7_  &  i_6_  &  n_n111  &  _31305 ) | ( (~ i_7_)  &  i_6_  &  n_n111  &  _31305 ) | ( i_7_  &  (~ i_6_)  &  n_n111  &  _31305 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n111  &  _31305 ) ;
 assign _31319 = ( i_7_  &  i_6_  &  n_n219  &  _30896 ) | ( (~ i_7_)  &  i_6_  &  n_n219  &  _30896 ) | ( i_7_  &  (~ i_6_)  &  n_n219  &  _30896 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n219  &  _30896 ) ;
 assign _31321 = ( wire3257 ) | ( wire3256 ) ;
 assign _31328 = ( wire18499 ) | ( wire18512 ) | ( wire3244 ) | ( _31286 ) ;
 assign _31330 = ( wire147  &  n_n123 ) | ( n_n123  &  wire46 ) ;
 assign _31334 = ( wire146  &  n_n125 ) | ( n_n125  &  wire46 ) ;
 assign _31338 = ( n_n218  &  n_n220  &  n_n126 ) ;
 assign _31340 = ( wire146  &  n_n123 ) | ( wire127  &  n_n123 ) ;
 assign _31342 = ( _2909 ) | ( _31334 ) | ( wire1465  &  _31338 ) ;
 assign _31343 = ( wire3229 ) | ( _2901 ) | ( _2906 ) | ( _31340 ) ;
 assign _31356 = ( n_n123  &  wire125 ) | ( n_n123  &  wire242 ) ;
 assign _31360 = ( n_n218  &  n_n220  &  n_n126 ) ;
 assign _31365 = ( _2884 ) | ( _31356 ) | ( wire1336  &  _31360 ) ;
 assign _31368 = ( wire154  &  n_n125 ) | ( n_n125  &  wire181 ) ;
 assign _31372 = ( n_n218  &  n_n124  &  n_n220 ) ;
 assign _31374 = ( wire63  &  n_n125 ) | ( wire48  &  n_n125 ) ;
 assign _31376 = ( _2866 ) | ( _31368 ) | ( wire1695  &  _31372 ) ;
 assign _31377 = ( wire3201 ) | ( _2858 ) | ( _2863 ) | ( _31374 ) ;
 assign _31378 = ( wire18555 ) | ( wire18546 ) | ( _2890 ) | ( _2894 ) ;
 assign _31381 = ( wire18526 ) | ( wire18565 ) | ( _31342 ) | ( _31343 ) ;
 assign _31382 = ( i_5_  &  i_3_  &  i_4_ ) ;
 assign _31392 = ( (~ i_7_)  &  i_6_  &  i_3_  &  i_4_ ) ;
 assign _31423 = ( wire55  &  n_n212 ) | ( wire158  &  n_n212 ) ;
 assign _31433 = ( n_n5011 ) | ( wire591 ) | ( wire18679 ) | ( _2787 ) ;
 assign _31435 = ( n_n108  &  wire211 ) | ( n_n108  &  wire107 ) ;
 assign _31437 = ( n_n108  &  wire205 ) | ( n_n108  &  wire225 ) ;
 assign _31442 = ( _2775 ) | ( _2781 ) | ( _31435 ) | ( _31437 ) ;
 assign _31445 = ( n_n108  &  wire84 ) | ( n_n108  &  wire220 ) ;
 assign _31446 = ( n_n4996 ) | ( wire234  &  _30050 ) ;
 assign _31450 = ( wire1862  &  _29356 ) | ( wire141  &  _30036 ) ;
 assign _31455 = ( n_n184  &  wire719 ) | ( n_n184  &  wire728 ) ;
 assign _31468 = ( n_n108  &  wire240 ) | ( n_n108  &  wire187 ) ;
 assign _31494 = ( wire18692 ) | ( wire18691 ) ;
 assign _31496 = ( wire18682 ) | ( wire18683 ) | ( wire18694 ) | ( _31494 ) ;
 assign _31512 = ( i_9_  &  (~ i_10_)  &  (~ i_11_) ) ;
 assign _31554 = ( wire3469 ) | ( wire18711 ) | ( wire18712 ) | ( _2679 ) ;
 assign _31555 = ( wire18214 ) | ( wire18719 ) | ( _31554 ) ;
 assign _31567 = ( n_n162  &  n_n35  &  n_n220 ) ;
 assign _31569 = ( n_n162  &  n_n35  &  n_n220 ) ;
 assign _31572 = ( wire4427 ) | ( wire144  &  _31569 ) ;
 assign _31586 = ( n_n31  &  wire120 ) | ( wire729  &  n_n31  &  _30673 ) ;
 assign _31588 = ( n_n31  &  wire116 ) | ( n_n31  &  wire198 ) ;
 assign _31592 = ( _2591 ) | ( _2597 ) | ( _31586 ) | ( _31588 ) ;
 assign _31594 = ( n_n31  &  wire179 ) | ( n_n31  &  wire184 ) ;
 assign _31600 = ( n_n5144 ) | ( wire18726 ) | ( _31592 ) ;
 assign _31614 = ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire725 ) ;
 assign _31615 = ( n_n32  &  _31080 ) | ( n_n33  &  _31614 ) ;
 assign _31624 = ( wire18763 ) | ( n_n33  &  wire147 ) | ( n_n33  &  wire158 ) ;
 assign _31632 = ( wire18755 ) | ( wire18767 ) | ( _2561 ) | ( _31624 ) ;
 assign _31662 = ( wire2953 ) | ( wire3550 ) | ( wire18816 ) | ( _2519 ) ;
 assign _31663 = ( _31662 ) | ( wire18815 ) ;
 assign _31664 = ( n_n3179 ) | ( wire18434 ) | ( _31195 ) | ( _31663 ) ;
 assign _31754 = ( wire2785 ) | ( wire147  &  n_n123 ) | ( n_n123  &  wire18944 ) ;
 assign _31770 = ( n_n123  &  wire1242 ) | ( wire729  &  n_n123  &  _29731 ) ;
 assign _31801 = ( wire18938 ) | ( wire18939 ) | ( wire18934 ) | ( _31770 ) ;
 assign _31819 = ( i_7_  &  (~ i_6_)  &  n_n218  &  wire714 ) ;
 assign _31826 = ( n_n197  &  wire326 ) | ( n_n197  &  wire327 ) ;
 assign _31830 = ( n_n218  &  n_n220  &  n_n200 ) ;
 assign _31832 = ( n_n212  &  wire331 ) | ( n_n212  &  wire312 ) ;
 assign _31833 = ( wire1132  &  _31819 ) | ( wire1129  &  _31830 ) ;
 assign _31834 = ( _2332 ) | ( _2335 ) | ( _31826 ) | ( _31832 ) ;
 assign _31883 = ( i_9_  &  (~ i_10_)  &  i_11_  &  wire721 ) | ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire721 ) | ( (~ i_9_)  &  (~ i_10_)  &  (~ i_11_)  &  wire721 ) ;
 assign _31887 = ( wire2817 ) | ( wire18911 ) | ( wire18925 ) | ( wire18928 ) ;
 assign _31890 = ( n_n1803 ) | ( wire18949 ) | ( wire18951 ) | ( _31754 ) ;
 assign _31892 = ( (~ i_9_)  &  i_10_  &  (~ i_11_) ) ;
 assign _31894 = ( n_n40  &  wire347 ) | ( wire715  &  n_n40  &  _31892 ) ;
 assign _31899 = ( wire2900 ) | ( n_n41  &  wire347 ) | ( n_n41  &  wire18859 ) ;
 assign _31900 = ( wire2897 ) | ( _2250 ) | ( _2264 ) | ( _31894 ) ;
 assign _31910 = ( n_n48  &  n_n220  &  n_n126 ) ;
 assign _31923 = ( i_7_  &  (~ i_6_)  &  n_n48  &  wire714 ) ;
 assign _31932 = ( wire1126  &  _31910 ) | ( wire988  &  _31923 ) ;
 assign _31940 = ( wire143  &  n_n34 ) | ( wire729  &  n_n34  &  _29252 ) ;
 assign _31946 = ( wire18857 ) | ( wire2910 ) | ( wire18850 ) | ( _31932 ) ;
 assign _31961 = ( wire146  &  n_n34 ) | ( n_n34  &  wire147 ) ;
 assign _31977 = ( (~ i_9_)  &  i_10_  &  (~ i_11_)  &  (~ i_15_) ) ;
 assign _31978 = ( i_9_  &  i_10_  &  i_11_  &  i_15_ ) ;
 assign _31998 = ( wire2853 ) | ( wire18895 ) | ( _2182 ) | ( _31961 ) ;
 assign _32003 = ( n_n40  &  wire230 ) | ( n_n40  &  wire400 ) ;
 assign _32019 = ( i_7_  &  (~ i_6_)  &  n_n48  &  wire714 ) ;
 assign _32025 = ( n_n40  &  wire261 ) | ( n_n40  &  wire375 ) ;
 assign _32040 = ( wire2724 ) | ( _32025 ) | ( wire1735  &  _32019 ) ;
 assign _32062 = ( _2060 ) | ( _2059 ) ;
 assign _32066 = ( n_n48  &  n_n220  &  n_n161 ) ;
 assign _32068 = ( n_n47  &  wire303 ) | ( n_n47  &  wire321 ) ;
 assign _32081 = ( wire18972 ) | ( wire18973 ) | ( wire1201  &  _32066 ) ;
 assign _32090 = ( n_n108  &  wire310 ) | ( n_n108  &  wire400 ) ;
 assign _32094 = ( n_n162  &  n_n220  &  n_n126 ) ;
 assign _32108 = ( _2020 ) | ( _32090 ) | ( wire1498  &  _32094 ) ;
 assign _32110 = ( wire18981 ) | ( wire19003 ) | ( _2026 ) | ( _32062 ) ;
 assign _32114 = ( (~ i_9_)  &  i_10_  &  i_11_  &  wire721 ) ;
 assign _32115 = ( i_9_  &  i_10_  &  i_11_  &  wire721 ) | ( (~ i_9_)  &  (~ i_10_)  &  (~ i_11_)  &  wire721 ) ;
 assign _32140 = ( i_9_  &  i_10_  &  (~ i_11_)  &  wire729 ) | ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire729 ) ;
 assign _32141 = ( n_n2  &  wire87 ) | ( wire729  &  n_n2  &  _29028 ) ;
 assign _32149 = ( wire18834 ) | ( _1972 ) | ( _1978 ) | ( _32141 ) ;
 assign _32161 = ( wire2704 ) | ( wire2705 ) ;
 assign _32183 = ( wire18832 ) | ( wire19031 ) | ( _1990 ) | ( _32161 ) ;
 assign _32185 = ( n_n5144 ) | ( wire18846 ) | ( wire19034 ) | ( _32183 ) ;
 assign _32227 = ( n_n162  &  n_n220  &  n_n126 ) ;
 assign _32230 = ( n_n5011 ) | ( wire2480 ) | ( wire2481 ) | ( _1871 ) ;
 assign _32240 = ( (~ i_9_)  &  (~ i_10_)  &  i_11_  &  (~ i_15_) ) ;
 assign _32241 = ( (~ i_9_)  &  (~ i_10_)  &  i_11_  &  i_15_ ) ;
 assign _32250 = ( i_7_  &  i_6_  &  n_n48  &  wire714 ) ;
 assign _32288 = ( wire19343 ) | ( wire19344 ) | ( wire19346 ) ;
 assign _32293 = ( n_n218  &  n_n220  &  n_n126 ) ;
 assign _32297 = ( n_n218  &  n_n124  &  n_n220 ) ;
 assign _32302 = ( n_n218  &  n_n124  &  n_n220 ) ;
 assign _32304 = ( wire1562  &  _32297 ) | ( wire1251  &  _32302 ) ;
 assign _32314 = ( n_n218  &  n_n124  &  n_n220 ) ;
 assign _32327 = ( wire2598 ) | ( _1721 ) | ( wire844  &  _32314 ) ;
 assign _32330 = ( wire2548 ) | ( wire19208 ) | ( wire928  &  _32293 ) ;
 assign _32331 = ( (~ i_9_)  &  (~ i_10_)  &  i_11_  &  wire729 ) ;
 assign _32341 = ( n_n1717 ) | ( wire2578 ) | ( n_n123  &  _32331 ) ;
 assign _32343 = ( n_n123  &  wire184 ) | ( n_n123  &  wire246 ) ;
 assign _32344 = ( n_n125  &  wire155 ) | ( wire729  &  n_n125  &  _29731 ) ;
 assign _32351 = ( wire2588 ) | ( _1676 ) | ( _32343 ) | ( _32344 ) ;
 assign _32363 = ( n_n101  &  wire276 ) | ( n_n101  &  wire211 ) ;
 assign _32372 = ( wire143  &  n_n108 ) | ( wire154  &  n_n108 ) ;
 assign _32380 = ( wire19190 ) | ( _1643 ) | ( _32363 ) | ( _32372 ) ;
 assign _32382 = ( wire2579 ) | ( wire19200 ) | ( _1648 ) | ( _32341 ) ;
 assign _32401 = ( i_7_  &  (~ i_6_)  &  n_n218  &  wire714 ) ;
 assign _32406 = ( i_7_  &  (~ i_6_)  &  n_n218  &  wire714 ) ;
 assign _32408 = ( wire1560  &  _32401 ) | ( wire1558  &  _32406 ) ;
 assign _32410 = ( wire2518 ) | ( wire19238 ) | ( wire19239 ) | ( _1581 ) ;
 assign _32412 = ( wire2545 ) | ( wire19213 ) | ( wire19272 ) | ( wire19273 ) ;
 assign _32417 = ( wire2537 ) | ( n_n197  &  wire70 ) ;
 assign _32419 = ( n_n197  &  wire63 ) | ( n_n197  &  wire184 ) ;
 assign _32421 = ( n_n197  &  wire246 ) | ( n_n197  &  wire233 ) ;
 assign _32426 = ( _1544 ) | ( _1549 ) | ( _32419 ) | ( _32421 ) ;
 assign _32437 = ( n_n218  &  n_n220  &  n_n200 ) ;
 assign _32442 = ( n_n218  &  n_n220  &  n_n200 ) ;
 assign _32447 = ( n_n218  &  n_n220  &  n_n200 ) ;
 assign _32450 = ( wire1292  &  _32437 ) | ( wire1290  &  _32442 ) ;
 assign _32452 = ( wire19232 ) | ( wire19268 ) | ( _1533 ) | ( _32417 ) ;
 assign _32454 = ( wire19210 ) | ( wire19276 ) | ( _32330 ) | ( _32412 ) ;
 assign _32472 = ( (~ i_7_)  &  (~ i_6_)  &  n_n218  &  wire714 ) ;
 assign _32474 = ( i_9_  &  (~ i_10_)  &  i_11_  &  wire720 ) ;
 assign _32477 = ( wire2404 ) | ( wire19405 ) | ( wire227  &  _32472 ) ;
 assign _32478 = ( (~ i_9_)  &  (~ i_10_)  &  (~ i_11_)  &  wire729 ) ;
 assign _32488 = ( wire2407 ) | ( wire19406 ) | ( _1404 ) | ( _32477 ) ;
 assign _32495 = ( n_n31  &  wire1537 ) | ( n_n31  &  wire19440 ) | ( n_n31  &  wire19441 ) ;
 assign _32504 = ( i_7_  &  (~ i_6_)  &  n_n48  &  wire714 ) ;
 assign _32509 = ( i_7_  &  (~ i_6_)  &  n_n48  &  wire714 ) ;
 assign _32510 = ( wire1556  &  _32504 ) | ( wire1404  &  _32509 ) ;
 assign _32514 = ( n_n41  &  wire227 ) | ( n_n41  &  wire221 ) ;
 assign _32515 = ( i_9_  &  i_10_  &  (~ i_11_)  &  (~ i_15_) ) ;
 assign _32516 = ( (~ i_9_)  &  (~ i_10_)  &  (~ i_11_)  &  i_15_ ) ;
 assign _32521 = ( n_n48  &  n_n220  &  n_n200 ) ;
 assign _32526 = ( n_n41  &  wire315 ) | ( n_n41  &  wire19411 ) | ( n_n41  &  wire19412 ) ;
 assign _32529 = ( _1455 ) | ( _32514 ) | ( wire1211  &  _32521 ) ;
 assign _32536 = ( n_n31  &  wire232 ) | ( n_n31  &  wire221 ) ;
 assign _32540 = ( wire2352 ) | ( wire2353 ) | ( _1411 ) | ( _32536 ) ;
 assign _32541 = ( n_n1163 ) | ( wire2364 ) | ( wire2365 ) | ( wire19429 ) ;
 assign _32548 = ( n_n46  &  wire49 ) | ( n_n46  &  wire19113 ) ;
 assign _32550 = ( n_n46  &  wire72 ) | ( n_n46  &  wire19104 ) ;
 assign _32554 = ( i_7_  &  i_6_  &  n_n48  &  wire714 ) ;
 assign _32558 = ( n_n48  &  n_n220  &  n_n161 ) ;
 assign _32562 = ( wire1503  &  _32554 ) | ( wire1500  &  _32558 ) ;
 assign _32577 = ( wire2636 ) | ( _1347 ) | ( _32548 ) | ( _32550 ) ;
 assign _32580 = ( n_n5109 ) | ( wire677 ) | ( wire19123 ) ;
 assign _32583 = ( wire518 ) | ( n_n3415 ) | ( wire2669 ) | ( _1307 ) ;
 assign _32603 = ( n_n4620 ) | ( wire2645 ) | ( n_n40  &  _31022 ) ;
 assign _32625 = ( wire2646 ) | ( _1308 ) | ( _32583 ) | ( _32603 ) ;
 assign _32636 = ( n_n36  &  wire232 ) | ( n_n36  &  wire221 ) ;
 assign _32643 = ( n_n218  &  n_n35  &  n_n220 ) ;
 assign _32647 = ( n_n36  &  wire845 ) | ( wire1143  &  _32643 ) ;
 assign _32649 = ( wire2703 ) | ( _1239 ) | ( _32636 ) | ( _32647 ) ;
 assign _32651 = ( n_n5144 ) | ( _1262 ) | ( _1263 ) | ( _1264 ) ;
 assign _32652 = ( wire2691 ) | ( wire19054 ) | ( _1242 ) | ( _32651 ) ;
 assign _32654 = ( n_n31  &  wire206 ) | ( n_n31  &  wire328 ) ;
 assign _32657 = ( n_n1434 ) | ( _1208 ) | ( _32654 ) ;
 assign _32665 = ( (~ i_9_)  &  i_10_  &  (~ i_11_)  &  i_15_ ) ;
 assign _32666 = ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  (~ i_15_) ) ;
 assign _32675 = ( n_n218  &  n_n35  &  n_n220 ) ;
 assign _32677 = ( n_n38  &  n_n54 ) | ( n_n39  &  n_n54 ) | ( n_n38  &  n_n52 ) | ( n_n39  &  n_n52 ) ;
 assign _32682 = ( n_n48  &  n_n220  &  n_n126 ) ;
 assign _32695 = ( wire19057 ) | ( wire19125 ) | ( _32580 ) | ( _32652 ) ;
 assign _32697 = ( wire19347 ) | ( wire19455 ) | ( wire19456 ) | ( _32288 ) ;
 assign _32719 = ( (~ i_7_)  &  (~ i_6_)  &  n_n162  &  wire714 ) ;
 assign _32764 = ( n_n799 ) | ( wire2310 ) | ( wire1809  &  _32719 ) ;
 assign _32769 = ( n_n124  &  n_n48  &  n_n220 ) ;
 assign _32771 = ( n_n124  &  n_n48  &  n_n220 ) ;
 assign _32772 = ( wire279  &  _32769 ) | ( wire207  &  _32771 ) ;
 assign _32802 = ( i_7_  &  (~ i_6_)  &  n_n48  &  wire714 ) ;
 assign _32808 = ( n_n39  &  _29204 ) | ( wire1630  &  _32802 ) ;
 assign _32812 = ( n_n817 ) | ( wire19556 ) | ( wire19557 ) ;
 assign _32815 = ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire719 ) ;
 assign _32818 = ( n_n42  &  n_n190 ) | ( n_n42  &  wire187 ) | ( n_n42  &  wire339 ) ;
 assign _32832 = ( wire2232 ) | ( n_n41  &  wire151 ) | ( n_n41  &  wire322 ) ;
 assign _32837 = ( n_n48  &  n_n220  &  n_n200 ) ;
 assign _32839 = ( n_n41  &  wire124 ) | ( n_n41  &  wire165 ) ;
 assign _32841 = ( n_n40  &  wire48 ) | ( n_n40  &  wire167 ) ;
 assign _32844 = ( _1021 ) | ( _32839 ) | ( wire1628  &  _32837 ) ;
 assign _32845 = ( n_n832 ) | ( wire19569 ) | ( wire19574 ) | ( _32832 ) ;
 assign _32856 = ( wire19588 ) | ( wire19587 ) ;
 assign _32877 = ( n_n47  &  wire134 ) | ( n_n47  &  wire194 ) ;
 assign _32880 = ( n_n834 ) | ( wire19591 ) | ( wire19582 ) | ( _32856 ) ;
 assign _32881 = ( wire19596 ) | ( wire19581 ) | ( n_n46  &  wire1674 ) ;
 assign _32918 = ( wire2182 ) | ( wire19614 ) | ( wire19617 ) ;
 assign _32919 = ( wire19560 ) | ( _32812 ) | ( _32844 ) | ( _32845 ) ;
 assign _32920 = ( wire19619 ) | ( _32880 ) | ( _32881 ) | ( _32918 ) ;
 assign _32999 = ( i_9_  &  (~ i_10_)  &  i_11_  &  wire724 ) ;
 assign _33004 = ( n_n34  &  n_n176 ) | ( n_n34  &  wire19528 ) | ( n_n34  &  _32999 ) ;
 assign _33013 = ( wire2282 ) | ( wire2283 ) | ( _823 ) | ( _33004 ) ;
 assign _33033 = ( n_n162  &  n_n220  &  n_n126 ) ;
 assign _33038 = ( n_n162  &  n_n124  &  n_n220 ) ;
 assign _33048 = ( wire1741  &  _33033 ) | ( wire1017  &  _33038 ) ;
 assign _33099 = ( wire19636 ) | ( wire19656 ) | ( _745 ) | ( _778 ) ;
 assign _33101 = ( wire19674 ) | ( wire19676 ) | ( n_n123  &  wire1775 ) ;
 assign _33104 = ( n_n31  &  wire104 ) | ( n_n31  &  wire279 ) ;
 assign _33117 = ( n_n162  &  n_n35  &  n_n220 ) ;
 assign _33122 = ( (~ i_7_)  &  (~ i_6_)  &  n_n162  &  wire714 ) ;
 assign _33138 = ( wire1305  &  _33117 ) | ( wire1302  &  _33122 ) ;
 assign _33161 = ( n_n5144 ) | ( wire213  &  wire775 ) ;
 assign _33162 = ( wire19687 ) | ( _696 ) | ( _33104 ) | ( _33161 ) ;
 assign _33163 = ( wire2335 ) | ( wire2350 ) | ( wire2351 ) | ( _33162 ) ;
 assign _33164 = ( wire19504 ) | ( wire19479 ) | ( _32764 ) | ( _33163 ) ;
 assign _33165 = ( _32919 ) | ( _32920 ) | ( _33164 ) ;
 assign _33185 = ( wire244  &  n_n39 ) | ( n_n39  &  wire19706 ) ;
 assign _33212 = ( n_n38  &  n_n54 ) | ( n_n39  &  n_n54 ) | ( n_n38  &  n_n52 ) | ( n_n39  &  n_n52 ) ;
 assign _33214 = ( n_n48  &  n_n220  &  n_n126 ) ;
 assign _33216 = ( n_n124  &  n_n48  &  n_n220 ) ;
 assign _33217 = ( wire140  &  _33214 ) | ( wire244  &  _33216 ) ;
 assign _33218 = ( n_n38  &  wire235 ) | ( n_n39  &  wire235 ) | ( n_n38  &  wire236 ) | ( n_n39  &  wire236 ) ;
 assign _33220 = ( _596 ) | ( _33212 ) | ( _33217 ) | ( _33218 ) ;
 assign _33223 = ( wire19702 ) | ( n_n41  &  wire1446 ) ;
 assign _33239 = ( wire137  &  n_n36 ) | ( n_n36  &  wire63 ) ;
 assign _33261 = ( wire19718 ) | ( wire19730 ) | ( wire19731 ) | ( _33239 ) ;
 assign _33275 = ( n_n40  &  wire166 ) | ( n_n40  &  wire278 ) ;
 assign _33286 = ( n_n41  &  wire275 ) | ( n_n41  &  wire278 ) ;
 assign _33287 = ( i_9_  &  i_10_  &  i_11_  &  wire726 ) ;
 assign _33291 = ( _499 ) | ( _511 ) | ( _33275 ) | ( _33286 ) ;
 assign _33293 = ( n_n42  &  wire63 ) | ( n_n42  &  n_n190 ) | ( n_n42  &  wire348 ) ;
 assign _33351 = ( wire19799 ) | ( _461 ) | ( _462 ) ;
 assign _33353 = ( n_n123  &  wire408 ) | ( n_n123  &  wire19850 ) ;
 assign _33354 = ( (~ i_9_)  &  i_10_  &  (~ i_11_)  &  wire726 ) ;
 assign _33361 = ( wire1949 ) | ( n_n125  &  wire249 ) | ( n_n125  &  _33354 ) ;
 assign _33362 = ( wire1945 ) | ( _409 ) | ( _422 ) | ( _33353 ) ;
 assign _33400 = ( wire19846 ) | ( wire19841 ) | ( wire19842 ) | ( wire19845 ) ;
 assign _33401 = ( wire19858 ) | ( _360 ) | ( _33361 ) | ( _33362 ) ;
 assign _33461 = ( n_n162  &  n_n124  &  n_n220 ) ;
 assign _33464 = ( n_n101  &  wire329 ) | ( n_n101  &  wire284 ) ;
 assign _33477 = ( _285 ) | ( _33464 ) | ( wire1613  &  _33461 ) ;
 assign _33487 = ( i_7_  &  (~ i_6_)  &  n_n218  &  wire714 ) ;
 assign _33489 = ( n_n197  &  wire283 ) | ( n_n197  &  wire325 ) ;
 assign _33493 = ( n_n218  &  n_n220  &  n_n200 ) ;
 assign _33495 = ( n_n212  &  wire325 ) | ( n_n212  &  wire354 ) ;
 assign _33496 = ( wire1363  &  _33487 ) | ( wire1354  &  _33493 ) ;
 assign _33497 = ( _252 ) | ( _255 ) | ( _33489 ) | ( _33495 ) ;
 assign _33528 = ( i_9_  &  (~ i_10_)  &  i_11_  &  wire728 ) | ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire728 ) | ( (~ i_9_)  &  (~ i_10_)  &  (~ i_11_)  &  wire728 ) ;
 assign _33535 = ( wire19823 ) | ( wire19837 ) | ( n_n123  &  wire1587 ) ;
 assign _33537 = ( wire19812 ) | ( _33351 ) | ( _33400 ) | ( _33401 ) ;
 assign _33543 = ( (~ i_7_)  &  (~ i_6_)  &  n_n162  &  wire714 ) ;
 assign _33561 = ( n_n162  &  n_n35  &  n_n220 ) ;
 assign _33568 = ( (~ i_7_)  &  (~ i_6_)  &  n_n162  &  wire714 ) ;
 assign _33578 = ( wire1590  &  _33561 ) | ( wire1483  &  _33568 ) ;
 assign _33612 = ( (~ i_7_)  &  (~ i_6_)  &  n_n162  &  wire714 ) ;
 assign _33614 = ( n_n33  &  wire282 ) | ( n_n33  &  wire236 ) ;
 assign _33626 = ( _143 ) | ( _33614 ) | ( wire1568  &  _33612 ) ;
 assign _33656 = ( wire2099 ) | ( wire19695 ) | ( wire19911 ) ;
 assign _33658 = ( wire19698 ) | ( wire19890 ) | ( wire19891 ) | ( _33656 ) ;
 assign _33659 = ( wire19907 ) | ( wire1592  &  _33543 ) ;
 assign _33662 = ( wire19869 ) | ( wire19914 ) | ( wire19867 ) | ( _33223 ) ;
 assign _33670 = ( (~ i_7_)  &  i_6_  &  n_n162  &  n_n219 ) | ( i_7_  &  (~ i_6_)  &  n_n162  &  n_n219 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n162  &  n_n219 ) ;
 assign _33681 = ( i_9_  &  i_10_  &  (~ i_11_)  &  wire729 ) | ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire729 ) ;
 assign _33709 = ( i_9_  &  i_10_  &  (~ i_11_)  &  wire729 ) | ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire729 ) ;
 assign _33710 = ( n_n3  &  wire87 ) | ( wire729  &  n_n3  &  _29028 ) ;


endmodule

