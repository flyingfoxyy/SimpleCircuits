module i10 (
	PV302_0_, PV301_0_, PV295_0_, PV294_0_, PV293_0_, PV292_0_, PV291_0_, PV290_0_, 
	PV289_0_, PV288_7_, PV288_6_, PV288_5_, PV288_4_, PV288_3_, PV288_2_, PV288_1_, PV288_0_, PV280_0_, 
	PV279_0_, PV278_0_, PV277_0_, PV275_0_, PV274_0_, PV272_0_, PV271_0_, PV270_0_, PV269_0_, PV268_5_, 
	PV268_4_, PV268_3_, PV268_2_, PV268_1_, PV268_0_, PV262_0_, PV261_0_, PV260_0_, PV259_0_, PV258_0_, 
	PV257_7_, PV257_6_, PV257_5_, PV257_4_, PV257_3_, PV257_2_, PV257_1_, PV257_0_, PV249_0_, PV248_0_, 
	PV247_0_, PV246_0_, PV245_0_, PV244_0_, PV243_0_, PV242_0_, PV241_0_, PV240_0_, PV239_4_, PV239_3_, 
	PV239_2_, PV239_1_, PV239_0_, PV234_4_, PV234_3_, PV234_2_, PV234_1_, PV234_0_, PV229_5_, PV229_4_, 
	PV229_3_, PV229_2_, PV229_1_, PV229_0_, PV223_5_, PV223_4_, PV223_3_, PV223_2_, PV223_1_, PV223_0_, 
	PV216_0_, PV215_0_, PV214_0_, PV213_5_, PV213_4_, PV213_3_, PV213_2_, PV213_1_, PV213_0_, PV207_0_, 
	PV205_0_, PV204_0_, PV203_0_, PV202_0_, PV199_4_, PV199_3_, PV199_2_, PV199_1_, PV199_0_, PV194_4_, 
	PV194_3_, PV194_2_, PV194_1_, PV194_0_, PV189_5_, PV189_4_, PV189_3_, PV189_2_, PV189_1_, PV189_0_, 
	PV183_5_, PV183_4_, PV183_3_, PV183_2_, PV183_1_, PV183_0_, PV177_0_, PV175_0_, PV174_0_, PV172_0_, 
	PV171_0_, PV169_1_, PV169_0_, PV165_7_, PV165_6_, PV165_5_, PV165_4_, PV165_3_, PV165_2_, PV165_1_, 
	PV165_0_, PV149_7_, PV149_6_, PV149_5_, PV149_4_, PV149_3_, PV149_2_, PV149_1_, PV149_0_, PV134_1_, 
	PV134_0_, PV132_7_, PV132_6_, PV132_5_, PV132_4_, PV132_3_, PV132_2_, PV132_1_, PV132_0_, PV124_5_, 
	PV124_4_, PV124_3_, PV124_2_, PV124_1_, PV124_0_, PV118_7_, PV118_6_, PV118_5_, PV118_4_, PV118_3_, 
	PV118_2_, PV118_1_, PV118_0_, PV110_0_, PV109_0_, PV108_5_, PV108_4_, PV108_3_, PV108_2_, PV108_1_, 
	PV108_0_, PV102_0_, PV101_0_, PV100_5_, PV100_4_, PV100_3_, PV100_2_, PV100_1_, PV100_0_, PV94_1_, 
	PV94_0_, PV91_1_, PV91_0_, PV88_3_, PV88_2_, PV88_1_, PV88_0_, PV84_5_, PV84_4_, PV84_3_, 
	PV84_2_, PV84_1_, PV84_0_, PV78_5_, PV78_4_, PV78_3_, PV78_2_, PV78_1_, PV78_0_, PV71_0_, 
	PV70_0_, PV69_0_, PV68_0_, PV67_0_, PV66_0_, PV65_0_, PV63_0_, PV62_0_, PV60_0_, PV59_0_, 
	PV57_0_, PV56_0_, PV55_0_, PV53_0_, PV52_0_, PV51_0_, PV50_0_, PV48_0_, PV46_0_, PV45_0_, 
	PV44_0_, PV43_0_, PV42_0_, PV41_0_, PV40_0_, PV39_0_, PV38_0_, PV37_0_, PV35_0_, PV34_0_, 
	PV33_0_, PV32_11_, PV32_10_, PV32_9_, PV32_8_, PV32_7_, PV32_6_, PV32_5_, PV32_4_, PV32_3_, 
	PV32_2_, PV32_1_, PV32_0_, PV16_0_, PV15_0_, PV14_0_, PV13_0_, PV12_0_, PV11_0_, PV10_0_, 
	PV9_0_, PV8_0_, PV7_0_, PV6_0_, PV5_0_, PV4_0_, PV3_0_, PV2_0_, PV1_0_, PV1992_1_, 
	PV1992_0_, PV1968_0_, PV1960_1_, PV1960_0_, PV1953_7_, PV1953_6_, PV1953_5_, PV1953_4_, PV1953_3_, PV1953_2_, 
	PV1953_1_, PV1953_0_, PV1921_5_, PV1921_4_, PV1921_3_, PV1921_2_, PV1921_1_, PV1921_0_, PV1901_0_, PV1900_0_, 
	PV1899_0_, PV1898_0_, PV1897_0_, PV1896_0_, PV1864_0_, PV1863_0_, PV1833_0_, PV1832, PV1829_9_, PV1829_8_, 
	PV1829_7_, PV1829_6_, PV1829_5_, PV1829_4_, PV1829_3_, PV1829_2_, PV1829_1_, PV1829_0_, PV1781_1_, PV1781_0_, 
	PV1771_1_, PV1771_0_, PV1760_0_, PV1759_0_, PV1758_0_, PV1757_0_, PV1745_0_, PV1741_0_, PV1736, PV1726_0_, 
	PV1719, PV1717_0_, PV1709_4_, PV1709_3_, PV1709_2_, PV1709_1_, PV1709_0_, PV1693_0_, PV1679_0_, PV1671_0_, 
	PV1669, PV1652_0_, PV1645_0_, PV1629_0_, PV1620_0_, PV1613_1_, PV1613_0_, PV1552_1_, PV1552_0_, PV1539, 
	PV1537, PV1536_0_, PV1512_3_, PV1512_2_, PV1512_1_, PV1495_0_, PV1492_0_, PV1481_0_, PV1480_0_, PV1470, 
	PV1467_0_, PV1459_0_, PV1451_0_, PV1440_0_, PV1439_0_, PV1432, PV1431, PV1429, PV1428, PV1426, 
	PV1423, PV1392_0_, PV1387, PV1386, PV1384, PV1382, PV1380, PV1378, PV1375, PV1374, 
	PV1373, PV1372, PV1371, PV1370, PV1365, PV1297_4_, PV1297_3_, PV1297_2_, PV1297_1_, PV1297_0_, 
	PV1281_0_, PV1274_0_, PV1267, PV1266, PV1265, PV1264, PV1263, PV1262, PV1261, PV1260, 
	PV1259, PV1258, PV1257, PV1256, PV1243_9_, PV1243_8_, PV1243_7_, PV1243_6_, PV1243_5_, PV1243_4_, 
	PV1243_3_, PV1243_2_, PV1243_1_, PV1243_0_, PV1213_11_, PV1213_10_, PV1213_9_, PV1213_8_, PV1213_7_, PV1213_6_, 
	PV1213_5_, PV1213_4_, PV1213_3_, PV1213_2_, PV1213_1_, PV1213_0_, PV986, PV966, PV826_0_, PV821_0_, 
	PV802_0_, PV801, PV798_0_, PV789, PV787, PV784, PV783, PV782, PV781, PV780, 
	PV779, PV778, PV775, PV763, PV707, PV657, PV656, PV655, PV654, PV653, 
	PV652, PV651, PV650, PV640_0_, PV634_0_, PV630, PV621, PV620, PV609_0_, PV603_0_, 
	PV597_0_, PV591_0_, PV587, PV585_0_, PV572_9_, PV572_8_, PV572_7_, PV572_6_, PV572_5_, PV572_4_, 
	PV572_3_, PV572_2_, PV572_1_, PV572_0_, PV548, PV547, PV546, PV545, PV544, PV543, 
	PV542, PV541, PV540, PV539, PV538, PV537, PV527, PV512, PV511_0_, PV508_0_, 
	PV500_0_, PV435_0_, PV432, PV423_0_, PV410_0_, PV398_0_, PV393_0_, PV377, PV375_0_, PV373, 
	PV357, PV356, PV321_2_);

input PV302_0_, PV301_0_, PV295_0_, PV294_0_, PV293_0_, PV292_0_, PV291_0_, PV290_0_, PV289_0_, PV288_7_, PV288_6_, PV288_5_, PV288_4_, PV288_3_, PV288_2_, PV288_1_, PV288_0_, PV280_0_, PV279_0_, PV278_0_, PV277_0_, PV275_0_, PV274_0_, PV272_0_, PV271_0_, PV270_0_, PV269_0_, PV268_5_, PV268_4_, PV268_3_, PV268_2_, PV268_1_, PV268_0_, PV262_0_, PV261_0_, PV260_0_, PV259_0_, PV258_0_, PV257_7_, PV257_6_, PV257_5_, PV257_4_, PV257_3_, PV257_2_, PV257_1_, PV257_0_, PV249_0_, PV248_0_, PV247_0_, PV246_0_, PV245_0_, PV244_0_, PV243_0_, PV242_0_, PV241_0_, PV240_0_, PV239_4_, PV239_3_, PV239_2_, PV239_1_, PV239_0_, PV234_4_, PV234_3_, PV234_2_, PV234_1_, PV234_0_, PV229_5_, PV229_4_, PV229_3_, PV229_2_, PV229_1_, PV229_0_, PV223_5_, PV223_4_, PV223_3_, PV223_2_, PV223_1_, PV223_0_, PV216_0_, PV215_0_, PV214_0_, PV213_5_, PV213_4_, PV213_3_, PV213_2_, PV213_1_, PV213_0_, PV207_0_, PV205_0_, PV204_0_, PV203_0_, PV202_0_, PV199_4_, PV199_3_, PV199_2_, PV199_1_, PV199_0_, PV194_4_, PV194_3_, PV194_2_, PV194_1_, PV194_0_, PV189_5_, PV189_4_, PV189_3_, PV189_2_, PV189_1_, PV189_0_, PV183_5_, PV183_4_, PV183_3_, PV183_2_, PV183_1_, PV183_0_, PV177_0_, PV175_0_, PV174_0_, PV172_0_, PV171_0_, PV169_1_, PV169_0_, PV165_7_, PV165_6_, PV165_5_, PV165_4_, PV165_3_, PV165_2_, PV165_1_, PV165_0_, PV149_7_, PV149_6_, PV149_5_, PV149_4_, PV149_3_, PV149_2_, PV149_1_, PV149_0_, PV134_1_, PV134_0_, PV132_7_, PV132_6_, PV132_5_, PV132_4_, PV132_3_, PV132_2_, PV132_1_, PV132_0_, PV124_5_, PV124_4_, PV124_3_, PV124_2_, PV124_1_, PV124_0_, PV118_7_, PV118_6_, PV118_5_, PV118_4_, PV118_3_, PV118_2_, PV118_1_, PV118_0_, PV110_0_, PV109_0_, PV108_5_, PV108_4_, PV108_3_, PV108_2_, PV108_1_, PV108_0_, PV102_0_, PV101_0_, PV100_5_, PV100_4_, PV100_3_, PV100_2_, PV100_1_, PV100_0_, PV94_1_, PV94_0_, PV91_1_, PV91_0_, PV88_3_, PV88_2_, PV88_1_, PV88_0_, PV84_5_, PV84_4_, PV84_3_, PV84_2_, PV84_1_, PV84_0_, PV78_5_, PV78_4_, PV78_3_, PV78_2_, PV78_1_, PV78_0_, PV71_0_, PV70_0_, PV69_0_, PV68_0_, PV67_0_, PV66_0_, PV65_0_, PV63_0_, PV62_0_, PV60_0_, PV59_0_, PV57_0_, PV56_0_, PV55_0_, PV53_0_, PV52_0_, PV51_0_, PV50_0_, PV48_0_, PV46_0_, PV45_0_, PV44_0_, PV43_0_, PV42_0_, PV41_0_, PV40_0_, PV39_0_, PV38_0_, PV37_0_, PV35_0_, PV34_0_, PV33_0_, PV32_11_, PV32_10_, PV32_9_, PV32_8_, PV32_7_, PV32_6_, PV32_5_, PV32_4_, PV32_3_, PV32_2_, PV32_1_, PV32_0_, PV16_0_, PV15_0_, PV14_0_, PV13_0_, PV12_0_, PV11_0_, PV10_0_, PV9_0_, PV8_0_, PV7_0_, PV6_0_, PV5_0_, PV4_0_, PV3_0_, PV2_0_, PV1_0_;

output PV1992_1_, PV1992_0_, PV1968_0_, PV1960_1_, PV1960_0_, PV1953_7_, PV1953_6_, PV1953_5_, PV1953_4_, PV1953_3_, PV1953_2_, PV1953_1_, PV1953_0_, PV1921_5_, PV1921_4_, PV1921_3_, PV1921_2_, PV1921_1_, PV1921_0_, PV1901_0_, PV1900_0_, PV1899_0_, PV1898_0_, PV1897_0_, PV1896_0_, PV1864_0_, PV1863_0_, PV1833_0_, PV1832, PV1829_9_, PV1829_8_, PV1829_7_, PV1829_6_, PV1829_5_, PV1829_4_, PV1829_3_, PV1829_2_, PV1829_1_, PV1829_0_, PV1781_1_, PV1781_0_, PV1771_1_, PV1771_0_, PV1760_0_, PV1759_0_, PV1758_0_, PV1757_0_, PV1745_0_, PV1741_0_, PV1736, PV1726_0_, PV1719, PV1717_0_, PV1709_4_, PV1709_3_, PV1709_2_, PV1709_1_, PV1709_0_, PV1693_0_, PV1679_0_, PV1671_0_, PV1669, PV1652_0_, PV1645_0_, PV1629_0_, PV1620_0_, PV1613_1_, PV1613_0_, PV1552_1_, PV1552_0_, PV1539, PV1537, PV1536_0_, PV1512_3_, PV1512_2_, PV1512_1_, PV1495_0_, PV1492_0_, PV1481_0_, PV1480_0_, PV1470, PV1467_0_, PV1459_0_, PV1451_0_, PV1440_0_, PV1439_0_, PV1432, PV1431, PV1429, PV1428, PV1426, PV1423, PV1392_0_, PV1387, PV1386, PV1384, PV1382, PV1380, PV1378, PV1375, PV1374, PV1373, PV1372, PV1371, PV1370, PV1365, PV1297_4_, PV1297_3_, PV1297_2_, PV1297_1_, PV1297_0_, PV1281_0_, PV1274_0_, PV1267, PV1266, PV1265, PV1264, PV1263, PV1262, PV1261, PV1260, PV1259, PV1258, PV1257, PV1256, PV1243_9_, PV1243_8_, PV1243_7_, PV1243_6_, PV1243_5_, PV1243_4_, PV1243_3_, PV1243_2_, PV1243_1_, PV1243_0_, PV1213_11_, PV1213_10_, PV1213_9_, PV1213_8_, PV1213_7_, PV1213_6_, PV1213_5_, PV1213_4_, PV1213_3_, PV1213_2_, PV1213_1_, PV1213_0_, PV986, PV966, PV826_0_, PV821_0_, PV802_0_, PV801, PV798_0_, PV789, PV787, PV784, PV783, PV782, PV781, PV780, PV779, PV778, PV775, PV763, PV707, PV657, PV656, PV655, PV654, PV653, PV652, PV651, PV650, PV640_0_, PV634_0_, PV630, PV621, PV620, PV609_0_, PV603_0_, PV597_0_, PV591_0_, PV587, PV585_0_, PV572_9_, PV572_8_, PV572_7_, PV572_6_, PV572_5_, PV572_4_, PV572_3_, PV572_2_, PV572_1_, PV572_0_, PV548, PV547, PV546, PV545, PV544, PV543, PV542, PV541, PV540, PV539, PV538, PV537, PV527, PV512, PV511_0_, PV508_0_, PV500_0_, PV435_0_, PV432, PV423_0_, PV410_0_, PV398_0_, PV393_0_, PV377, PV375_0_, PV373, PV357, PV356, PV321_2_;

wire n4, n5, n6, n7, n8, n3, n9, n10, n11, n12, n13, n14, n15, n20, n18, n23, n22, n25, n27, n28, n32, n31, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n69, n66, n68, n70, n73, n71, n75, n74, n76, n78, n82, n84, n85, n87, n88, n89, n90, n86, n92, n93, n95, n91, n97, n98, n100, n96, n102, n103, n104, n105, n101, n107, n110, n106, n112, n113, n114, n115, n111, n117, n121, n120, n119, n122, n124, n129, n130, n131, n132, n133, n134, n135, n136, n142, n141, n145, n143, n147, n148, n149, n150, n151, n155, n153, n154, n152, n156, n157, n158, n159, n160, n163, n162, n164, n166, n167, n170, n169, n168, n172, n176, n173, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n191, n193, n195, n196, n194, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n218, n219, n222, n223, n224, n225, n226, n229, n230, n228, n231, n234, n235, n236, n238, n239, n240, n242, n243, n247, n248, n250, n249, n253, n251, n257, n256, n255, n254, n258, n262, n261, n259, n265, n263, n267, n268, n269, n271, n270, n274, n272, n276, n278, n279, n283, n281, n280, n287, n285, n289, n288, n293, n291, n290, n295, n294, n298, n296, n300, n302, n304, n307, n305, n308, n313, n312, n310, n317, n315, n314, n320, n321, n319, n322, n324, n330, n327, n326, n332, n333, n331, n337, n336, n335, n339, n344, n342, n348, n346, n350, n351, n349, n355, n354, n353, n357, n360, n361, n364, n366, n370, n371, n372, n373, n374, n375, n380, n379, n376, n382, n381, n385, n384, n387, n386, n393, n392, n390, n394, n396, n395, n397, n399, n400, n401, n402, n403, n405, n409, n408, n411, n410, n414, n416, n419, n420, n418, n417, n423, n425, n426, n427, n429, n428, n431, n432, n433, n435, n436, n437, n441, n442, n439, n438, n444, n447, n448, n445, n450, n453, n454, n451, n456, n457, n460, n461, n465, n466, n463, n462, n470, n471, n468, n476, n477, n474, n473, n481, n482, n479, n486, n487, n484, n490, n491, n492, n493, n495, n496, n494, n497, n498, n499, n501, n503, n502, n506, n507, n505, n510, n508, n511, n522, n524, n523, n531, n532, n529, n534, n535, n538, n540, n544, n543, n542, n545, n554, n553, n556, n555, n558, n559, n563, n568, n567, n570, n571, n569, n575, n576, n574, n578, n579, n577, n581, n582, n580, n584, n585, n583, n586, n588, n600, n604, n603, n605, n606, n611, n610, n616, n614, n617, n621, n623, n622, n625, n624, n626, n627, n628, n629, n631, n630, n632, n633, n634, n637, n636, n638, n639, n642, n641, n643, n644, n646, n647, n645, n648, n649, n653, n651, n654, n655, n657, n658, n656, n660, n661, n662, n665, n664, n666, n667, n670, n669, n672, n673, n674, n675, n676, n678, n682, n685, n684, n688, n687, n691, n690, n694, n693, n695, n696, n699, n703, n704, n707, n710, n711, n714, n715, n717, n718, n720, n721, n722, n723, n725, n731, n730, n735, n736, n732, n739, n740, n744, n750, n748, n752, n754, n762, n763, n764, n765, n766, n775, n776, n777, n783, n787, n788, n791, n790, n792, n794, n795, n797, n801, n815, n824, n825, n826, n830, n831, n832, n833, n835, n839, n847, n849, n853, n854, n857, n859, n858, n861, n860, n863, n862, n864, n865, n866, n867, n869, n868, n871, n870, n873, n872, n874, n876, n875, n878, n879, n882, n881, n884, n883, n885, n887, n886, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n918, n917, n919, n920, n921, n922, n923, n924, n925, n926, n928, n930, n931, n932, n933, n934, n935, n936, n937, n939, n940, n943, n944, n946, n948, n949, n950, n951, n952, n953, n954, n955, n957, n959, n958, n961, n962, n963, n964, n965, n966, n971, n972, n974, n973, n976, n978, n980, n981, n982, n985, n986, n988, n987, n990, n992, n997, n1001, n1003, n1005, n1006, n1008, n1010, n1011, n1014, n1016, n1020, n1022, n1024, n1025, n1026, n1028, n1027, n1030, n1029, n1033;

assign PV1992_1_ = ( (~ n214) ) ;
 assign PV1992_0_ = ( (~ n920) ) ;
 assign PV1968_0_ = ( (~ n919) ) ;
 assign PV1960_1_ = ( (~ n628) ) ;
 assign PV1960_0_ = ( (~ n629) ) ;
 assign PV1953_7_ = ( (~ n207) ) ;
 assign PV1953_6_ = ( (~ n208) ) ;
 assign PV1953_5_ = ( (~ n209) ) ;
 assign PV1953_4_ = ( (~ n210) ) ;
 assign PV1953_3_ = ( (~ n211) ) ;
 assign PV1953_2_ = ( (~ n212) ) ;
 assign PV1953_1_ = ( PV132_1_  &  (~ n588) ) ;
 assign PV1953_0_ = ( (~ n213) ) ;
 assign PV1921_5_ = ( (~ n206) ) ;
 assign PV1921_4_ = ( (~ n569) ) ;
 assign PV1921_3_ = ( (~ n574) ) ;
 assign PV1921_2_ = ( (~ n577) ) ;
 assign PV1921_1_ = ( (~ n580) ) ;
 assign PV1921_0_ = ( (~ n583) ) ;
 assign PV1901_0_ = ( (~ n205) ) ;
 assign PV1900_0_ = ( (~ n204) ) ;
 assign PV1899_0_ = ( (~ n203) ) ;
 assign PV1898_0_ = ( (~ n202) ) ;
 assign PV1897_0_ = ( (~ n201) ) ;
 assign PV1896_0_ = ( (~ n200) ) ;
 assign PV1864_0_ = ( (~ PV302_0_) ) ;
 assign PV1863_0_ = ( (~ PV301_0_) ) ;
 assign PV1833_0_ = ( (~ PV261_0_) ) ;
 assign PV1832 = ( PV14_0_  &  n198 ) | ( PV14_0_  &  n199 ) ;
 assign PV1829_9_ = ( (~ n907) ) ;
 assign PV1829_8_ = ( (~ n908) ) ;
 assign PV1829_7_ = ( (~ n909) ) ;
 assign PV1829_6_ = ( (~ n910) ) ;
 assign PV1829_5_ = ( (~ n911) ) ;
 assign PV1829_4_ = ( (~ n912) ) ;
 assign PV1829_3_ = ( (~ n913) ) ;
 assign PV1829_2_ = ( (~ n914) ) ;
 assign PV1829_1_ = ( (~ n915) ) ;
 assign PV1829_0_ = ( (~ n916) ) ;
 assign PV1781_1_ = ( (~ n905) ) ;
 assign PV1781_0_ = ( (~ n906) ) ;
 assign PV1771_1_ = ( (~ n903) ) ;
 assign PV1771_0_ = ( (~ n904) ) ;
 assign PV1760_0_ = ( (~ PV101_0_) ) ;
 assign PV1759_0_ = ( (~ n197) ) ;
 assign PV1758_0_ = ( (~ n194) ) ;
 assign PV1745_0_ = ( (~ n228) ) ;
 assign PV1741_0_ = ( n191 ) | ( n193 ) | ( (~ n826) ) ;
 assign PV1736 = ( (~ PV290_0_)  &  (~ n177)  &  (~ n263) ) ;
 assign PV1726_0_ = ( (~ n187) ) ;
 assign PV1719 = ( PV240_0_  &  (~ PV172_0_)  &  (~ n239) ) ;
 assign PV1717_0_ = ( (~ n186) ) ;
 assign PV1709_4_ = ( (~ n181) ) ;
 assign PV1709_3_ = ( (~ n182) ) ;
 assign PV1709_2_ = ( (~ n183) ) ;
 assign PV1709_1_ = ( (~ n184) ) ;
 assign PV1709_0_ = ( (~ n185) ) ;
 assign PV1693_0_ = ( (~ n902) ) ;
 assign PV1679_0_ = ( n180 ) | ( n76 ) ;
 assign PV1671_0_ = ( (~ PV205_0_) ) ;
 assign PV1669 = ( n177  &  n178  &  n179 ) ;
 assign PV1652_0_ = ( (~ PV295_0_) ) | ( PV290_0_ ) | ( PV289_0_ ) | ( PV249_0_ ) | ( n122 ) | ( n231 ) ;
 assign PV1645_0_ = ( (~ n172) ) ;
 assign PV1629_0_ = ( (~ n167) ) ;
 assign PV1620_0_ = ( (~ n166) ) ;
 assign PV1613_1_ = ( (~ n703)  &  n704 ) | ( n703  &  (~ n704) ) ;
 assign PV1613_0_ = ( (~ n890)  &  n891 ) | ( n890  &  (~ n891) ) ;
 assign PV1552_1_ = ( (~ n626) ) ;
 assign PV1552_0_ = ( (~ n627) ) ;
 assign PV1539 = ( PV69_0_  &  (~ n824) ) | ( PV50_0_  &  (~ n824) ) ;
 assign PV1537 = ( PV68_0_  &  (~ n824) ) ;
 assign PV1536_0_ = ( n31 ) | ( n160 ) | ( (~ n732) ) ;
 assign PV1512_3_ = ( (~ n899) ) ;
 assign PV1512_2_ = ( (~ n900) ) ;
 assign PV1512_1_ = ( (~ n901) ) ;
 assign PV1495_0_ = ( (~ PV175_0_) ) ;
 assign PV1492_0_ = ( (~ n159) ) ;
 assign PV1481_0_ = ( (~ PV214_0_) ) ;
 assign PV1480_0_ = ( (~ n156) ) ;
 assign PV1470 = ( PV67_0_  &  n151  &  (~ n824) ) ;
 assign PV1467_0_ = ( PV14_0_  &  n150 ) ;
 assign PV1459_0_ = ( PV14_0_  &  n149 ) ;
 assign PV1451_0_ = ( n148  &  PV14_0_ ) ;
 assign PV1440_0_ = ( (~ PV14_0_) ) | ( n71 ) ;
 assign PV1439_0_ = ( (~ n147) ) ;
 assign PV1432 = ( PV66_0_  &  (~ n824) ) ;
 assign PV1431 = ( (~ PV109_0_)  &  PV1423 ) | ( PV13_0_  &  PV1423 ) ;
 assign PV1429 = ( PV12_0_  &  PV1_0_ ) ;
 assign PV1428 = ( PV11_0_  &  PV1_0_ ) ;
 assign PV1426 = ( n78  &  PV1_0_ ) ;
 assign PV1423 = ( PV9_0_  &  PV1_0_ ) ;
 assign PV1392_0_ = ( n142  &  (~ n824) ) | ( n141  &  (~ n253)  &  (~ n824) ) ;
 assign PV1387 = ( PV8_0_  &  PV9_0_ ) ;
 assign PV1386 = ( PV782  &  (~ n524) ) ;
 assign PV1384 = ( PV56_0_  &  PV782  &  (~ n152)  &  (~ n239)  &  (~ n721) ) ;
 assign PV1382 = ( PV782  &  n136 ) | ( PV782  &  (~ n390) ) ;
 assign PV1380 = ( (~ n135) ) ;
 assign PV1378 = ( PV782  &  n847 ) ;
 assign PV1375 = ( (~ PV268_5_) ) ;
 assign PV1374 = ( (~ PV268_5_)  &  PV268_4_ ) | ( PV268_5_  &  (~ PV268_4_) ) ;
 assign PV1373 = ( (~ PV268_3_)  &  n830 ) | ( PV268_3_  &  (~ n830) ) ;
 assign PV1372 = ( (~ PV268_2_)  &  n623 ) | ( PV268_2_  &  (~ n623) ) ;
 assign PV1371 = ( (~ PV268_1_)  &  n622 ) | ( PV268_1_  &  (~ n622) ) ;
 assign PV1370 = ( (~ n831)  &  PV268_0_ ) | ( n831  &  (~ PV268_0_) ) ;
 assign PV1365 = ( PV62_0_  &  (~ n122)  &  n223  &  n224  &  n225  &  n226  &  (~ n382)  &  (~ n824) ) ;
 assign PV1297_4_ = ( (~ n130) ) ;
 assign PV1297_3_ = ( (~ n131) ) ;
 assign PV1297_2_ = ( (~ n132) ) ;
 assign PV1297_1_ = ( (~ n133) ) ;
 assign PV1297_0_ = ( (~ n134) ) ;
 assign PV1281_0_ = ( (~ n898) ) ;
 assign PV1274_0_ = ( n129  &  (~ n824) ) | ( PV62_0_  &  (~ n410)  &  (~ n824) ) ;
 assign PV1267 = ( PV11_0_  &  PV2_0_ ) ;
 assign PV1266 = ( PV11_0_  &  PV4_0_ ) ;
 assign PV1265 = ( PV52_0_  &  PV1264 ) ;
 assign PV1264 = ( PV4_0_  &  PV12_0_ ) ;
 assign PV1263 = ( PV9_0_  &  PV4_0_ ) ;
 assign PV1262 = ( n78  &  PV4_0_ ) ;
 assign PV1261 = ( (~ PV62_0_)  &  PV1260 ) ;
 assign PV1260 = ( PV3_0_  &  PV11_0_ ) ;
 assign PV1259 = ( PV9_0_  &  PV3_0_ ) ;
 assign PV1258 = ( PV9_0_  &  PV2_0_ ) ;
 assign PV1257 = ( (~ PV174_0_)  &  (~ PV35_0_)  &  PV12_0_  &  PV2_0_  &  n124  &  (~ n164) ) ;
 assign PV1256 = ( n78  &  PV2_0_ ) ;
 assign PV1243_9_ = ( (~ n12) ) ;
 assign PV1243_8_ = ( (~ n10) ) ;
 assign PV1243_7_ = ( (~ n11) ) ;
 assign PV1243_6_ = ( (~ n56) ) ;
 assign PV1243_5_ = ( (~ n57) ) ;
 assign PV1243_4_ = ( (~ n58) ) ;
 assign PV1243_3_ = ( (~ n59) ) ;
 assign PV1243_2_ = ( (~ n60) ) ;
 assign PV1243_1_ = ( (~ n61) ) ;
 assign PV1243_0_ = ( (~ PV321_2_) ) ;
 assign PV1213_11_ = ( (~ n45) ) ;
 assign PV1213_10_ = ( (~ n44) ) ;
 assign PV1213_9_ = ( (~ n43) ) ;
 assign PV1213_8_ = ( (~ n42) ) ;
 assign PV1213_7_ = ( (~ n41) ) ;
 assign PV1213_6_ = ( (~ n40) ) ;
 assign PV1213_5_ = ( (~ n39) ) ;
 assign PV1213_4_ = ( (~ n494) ) ;
 assign PV1213_3_ = ( (~ n38) ) ;
 assign PV1213_2_ = ( (~ n37) ) ;
 assign PV1213_1_ = ( (~ n36) ) ;
 assign PV1213_0_ = ( (~ n35) ) ;
 assign PV986 = ( (~ n824)  &  (~ n955) ) | ( PV62_0_  &  n122  &  (~ n824) ) ;
 assign PV966 = ( n117  &  (~ n824) ) | ( (~ n824)  &  (~ n957) ) | ( (~ n824)  &  (~ n1010) ) ;
 assign PV826_0_ = ( (~ n897) ) ;
 assign PV821_0_ = ( (~ n896) ) ;
 assign PV802_0_ = ( PV51_0_ ) | ( PV52_0_ ) ;
 assign PV801 = ( n84  &  n85 ) ;
 assign PV798_0_ = ( PV302_0_ ) | ( PV289_0_ ) | ( PV214_0_ ) | ( n82 ) | ( n234 ) | ( n235 ) | ( n236 ) | ( (~ n923) ) ;
 assign PV789 = ( (~ PV202_0_)  &  PV1263 ) | ( (~ PV71_0_)  &  PV1263 ) | ( PV13_0_  &  PV1263 ) ;
 assign PV787 = ( PV9_0_  &  PV7_0_ ) ;
 assign PV784 = ( PV11_0_  &  PV7_0_ ) ;
 assign PV783 = ( PV11_0_  &  PV5_0_ ) ;
 assign PV782 = ( PV7_0_  &  n78 ) ;
 assign PV781 = ( PV12_0_  &  PV6_0_  &  (~ n606) ) ;
 assign PV780 = ( PV9_0_  &  PV6_0_ ) ;
 assign PV779 = ( n78  &  PV6_0_ ) ;
 assign PV778 = ( PV9_0_  &  PV5_0_ ) ;
 assign PV775 = ( PV70_0_  &  n76  &  (~ n253)  &  (~ n824) ) ;
 assign PV763 = ( (~ n253) ) ;
 assign PV707 = ( (~ n744) ) ;
 assign PV657 = ( (~ PV257_7_) ) ;
 assign PV656 = ( (~ PV257_7_)  &  PV257_6_ ) | ( PV257_7_  &  (~ PV257_6_) ) ;
 assign PV655 = ( (~ PV257_5_)  &  n853 ) | ( PV257_5_  &  (~ n853) ) ;
 assign PV654 = ( (~ PV257_4_)  &  n611 ) | ( PV257_4_  &  (~ n611) ) ;
 assign PV653 = ( (~ PV257_3_)  &  n610 ) | ( PV257_3_  &  (~ n610) ) ;
 assign PV652 = ( (~ PV257_2_)  &  n854 ) | ( PV257_2_  &  (~ n854) ) ;
 assign PV651 = ( (~ PV257_1_)  &  n75 ) | ( PV257_1_  &  (~ n75) ) ;
 assign PV650 = ( (~ n74)  &  PV257_0_ ) | ( n74  &  (~ PV257_0_) ) ;
 assign PV640_0_ = ( (~ n238) ) ;
 assign PV634_0_ = ( (~ n921) ) ;
 assign PV630 = ( (~ PV302_0_)  &  (~ PV62_0_)  &  (~ n405) ) | ( (~ PV302_0_)  &  n25  &  (~ n405) ) ;
 assign PV621 = ( n70  &  PV293_0_ ) ;
 assign PV620 = ( (~ PV56_0_)  &  n69 ) | ( n69  &  n66 ) | ( n69  &  n68 ) ;
 assign PV609_0_ = ( n65  &  n64 ) ;
 assign PV603_0_ = ( n63  &  n64 ) ;
 assign PV597_0_ = ( (~ n62) ) ;
 assign PV591_0_ = ( (~ n894) ) ;
 assign PV587 = ( (~ n460) ) ;
 assign PV585_0_ = ( (~ PV34_0_) ) ;
 assign PV572_9_ = ( (~ n46) ) ;
 assign PV572_8_ = ( (~ n47) ) ;
 assign PV572_7_ = ( (~ n48) ) ;
 assign PV572_6_ = ( (~ n49) ) ;
 assign PV572_5_ = ( (~ n50) ) ;
 assign PV572_4_ = ( (~ n51) ) ;
 assign PV572_3_ = ( (~ n52) ) ;
 assign PV572_2_ = ( (~ n53) ) ;
 assign PV572_1_ = ( (~ n54) ) ;
 assign PV572_0_ = ( (~ n55) ) ;
 assign PV548 = ( (~ n45)  &  (~ n73) ) ;
 assign PV547 = ( (~ n44)  &  (~ n73) ) ;
 assign PV546 = ( (~ n43)  &  (~ n73) ) ;
 assign PV545 = ( (~ n42)  &  (~ n73) ) ;
 assign PV544 = ( (~ n41)  &  (~ n73) ) ;
 assign PV543 = ( (~ n40)  &  (~ n73) ) ;
 assign PV542 = ( (~ n39)  &  (~ n73) ) ;
 assign PV541 = ( (~ n73)  &  (~ n494) ) ;
 assign PV540 = ( (~ n38)  &  (~ n73) ) ;
 assign PV539 = ( (~ n37)  &  (~ n73) ) ;
 assign PV538 = ( (~ n36)  &  (~ n73) ) ;
 assign PV537 = ( (~ n35)  &  (~ n73) ) ;
 assign PV527 = ( (~ n239)  &  (~ n240)  &  (~ n783) ) ;
 assign PV512 = ( (~ n1008) ) ;
 assign PV511_0_ = ( (~ n28) ) ;
 assign PV508_0_ = ( (~ n27) ) ;
 assign PV500_0_ = ( PV271_0_ ) | ( (~ PV14_0_) ) ;
 assign PV435_0_ = ( PV630 ) | ( (~ n1006) ) ;
 assign PV432 = ( (~ n1006) ) ;
 assign PV423_0_ = ( PV1719 ) | ( n13 ) | ( n14 ) | ( n15 ) | ( (~ n240) ) | ( (~ n930) ) ;
 assign PV410_0_ = ( n239 ) | ( PV15_0_ ) | ( n240 ) ;
 assign PV398_0_ = ( PV214_0_ ) | ( PV43_0_ ) | ( (~ PV423_0_) ) | ( n242 ) ;
 assign PV393_0_ = ( (~ n1005) ) ;
 assign PV377 = ( PV203_0_  &  PV35_0_ ) | ( PV203_0_  &  n9 ) ;
 assign PV375_0_ = ( PV1387 ) | ( PV1423 ) | ( PV1259 ) | ( PV1263 ) | ( PV787 ) | ( PV1258 ) | ( PV778 ) | ( PV780 ) ;
 assign PV373 = ( PV13_0_  &  PV10_0_ ) ;
 assign PV357 = ( n8  &  (~ n86)  &  (~ n96)  &  (~ n122)  &  n219  &  n222 ) ;
 assign PV356 = ( n6  &  n91  &  (~ n122)  &  n215  &  n216  &  n218  &  (~ n642) ) ;
 assign PV321_2_ = ( (~ PV78_4_)  &  n295 ) | ( n295  &  (~ n294) ) | ( (~ PV78_4_)  &  n417 ) | ( (~ n294)  &  n417 ) ;
 assign n4 = ( (~ n638) ) | ( n641 ) | ( n644 ) | ( n764 ) | ( n867 ) ;
 assign n5 = ( n638 ) | ( n641 ) | ( n643 ) | ( n764 ) | ( n866 ) ;
 assign n6 = ( (~ n38) ) | ( n763 ) ;
 assign n7 = ( n91  &  (~ n96)  &  n106  &  (~ n111) ) ;
 assign n8 = ( n38 ) | ( n763 ) ;
 assign n3 = ( n4  &  n5  &  n6  &  n7  &  n8 ) ;
 assign n9 = ( PV203_0_  &  PV165_2_  &  PV165_1_  &  (~ PV165_0_) ) ;
 assign n10 = ( n370  &  n371 ) ;
 assign n11 = ( n372  &  n373 ) ;
 assign n12 = ( n374  &  n375 ) ;
 assign n13 = ( PV174_0_  &  PV56_0_ ) | ( PV56_0_  &  (~ n291) ) ;
 assign n14 = ( n122  &  PV802_0_ ) | ( n122  &  PV59_0_ ) | ( n122  &  PV70_0_ ) ;
 assign n15 = ( (~ PV215_0_)  &  PV66_0_  &  (~ n239)  &  (~ n253) ) ;
 assign n20 = ( (~ PV88_3_) ) | ( (~ PV88_2_) ) ;
 assign n18 = ( (~ n744)  &  (~ n924) ) | ( n20  &  (~ n718)  &  (~ n744) ) ;
 assign n23 = ( n163  &  PV169_1_ ) ;
 assign n22 = ( PV802_0_  &  n23 ) | ( PV802_0_  &  (~ n253) ) ;
 assign n25 = ( n248 ) | ( n720 ) ;
 assign n27 = ( (~ PV59_0_)  &  n411 ) | ( n411  &  n410 ) ;
 assign n28 = ( (~ PV45_0_)  &  (~ PV40_0_) ) | ( PV43_0_  &  (~ PV40_0_) ) ;
 assign n32 = ( n723  &  PV207_0_ ) ;
 assign n31 = ( n32  &  (~ n267) ) | ( PV149_7_  &  PV56_0_  &  (~ n267) ) ;
 assign n35 = ( (~ PV183_0_)  &  n304 ) | ( n296  &  n304 ) ;
 assign n36 = ( (~ PV183_1_)  &  n298 ) | ( n298  &  n296 ) ;
 assign n37 = ( (~ PV183_2_)  &  n300 ) | ( n296  &  n300 ) ;
 assign n38 = ( (~ PV183_3_)  &  n302 ) | ( n296  &  n302 ) ;
 assign n39 = ( (~ PV32_5_)  &  n492  &  n493 ) | ( (~ n294)  &  n492  &  n493 ) ;
 assign n40 = ( (~ PV32_6_)  &  n490  &  n491 ) | ( (~ n294)  &  n490  &  n491 ) ;
 assign n41 = ( (~ PV32_7_)  &  n295 ) | ( n295  &  (~ n294) ) | ( (~ PV32_7_)  &  n484 ) | ( (~ n294)  &  n484 ) ;
 assign n42 = ( (~ PV32_8_)  &  n295 ) | ( n295  &  (~ n294) ) | ( (~ PV32_8_)  &  n479 ) | ( (~ n294)  &  n479 ) ;
 assign n43 = ( (~ PV32_9_)  &  n295 ) | ( n295  &  (~ n294) ) | ( (~ PV32_9_)  &  n473 ) | ( (~ n294)  &  n473 ) ;
 assign n44 = ( (~ PV32_10_)  &  n295 ) | ( n295  &  (~ n294) ) | ( (~ PV32_10_)  &  n468 ) | ( (~ n294)  &  n468 ) ;
 assign n45 = ( (~ PV32_11_)  &  n295 ) | ( n295  &  (~ n294) ) | ( (~ PV32_11_)  &  n462 ) | ( (~ n294)  &  n462 ) ;
 assign n46 = ( PV199_4_  &  n12 ) | ( PV199_4_  &  n414 ) | ( n12  &  (~ n790) ) | ( n414  &  (~ n790) ) ;
 assign n47 = ( n10  &  n416 ) | ( n414  &  n416 ) | ( n10  &  (~ n790) ) | ( n414  &  (~ n790) ) ;
 assign n48 = ( n11  &  n423 ) | ( n414  &  n423 ) | ( n11  &  (~ n790) ) | ( n414  &  (~ n790) ) ;
 assign n49 = ( n56  &  n427 ) | ( n414  &  n427 ) | ( n56  &  (~ n790) ) | ( n414  &  (~ n790) ) ;
 assign n50 = ( n57  &  n433 ) | ( n414  &  n433 ) | ( n57  &  (~ n790) ) | ( n414  &  (~ n790) ) ;
 assign n51 = ( n58  &  n437 ) | ( n414  &  n437 ) | ( n58  &  (~ n790) ) | ( n414  &  (~ n790) ) ;
 assign n52 = ( n444  &  n59 ) | ( n444  &  n414 ) ;
 assign n53 = ( n450  &  n60 ) | ( n450  &  n414 ) ;
 assign n54 = ( n456  &  n61 ) | ( n456  &  n414 ) ;
 assign n55 = ( n457  &  PV321_2_ ) | ( n457  &  n414 ) ;
 assign n56 = ( (~ PV84_4_)  &  n425  &  n426 ) | ( (~ n294)  &  n425  &  n426 ) ;
 assign n57 = ( (~ PV84_3_)  &  n431  &  n432 ) | ( (~ n294)  &  n431  &  n432 ) ;
 assign n58 = ( (~ PV84_2_)  &  n435  &  n436 ) | ( (~ n294)  &  n435  &  n436 ) ;
 assign n59 = ( (~ PV84_1_)  &  n295 ) | ( n295  &  (~ n294) ) | ( (~ PV84_1_)  &  n438 ) | ( (~ n294)  &  n438 ) ;
 assign n60 = ( (~ PV84_0_)  &  n295 ) | ( n295  &  (~ n294) ) | ( (~ PV84_0_)  &  n445 ) | ( (~ n294)  &  n445 ) ;
 assign n61 = ( (~ PV78_5_)  &  n295 ) | ( n295  &  (~ n294) ) | ( (~ PV78_5_)  &  n451 ) | ( (~ n294)  &  n451 ) ;
 assign n62 = ( (~ PV245_0_)  &  (~ n64) ) | ( (~ n64)  &  n460 ) | ( (~ PV245_0_)  &  (~ n895) ) | ( n460  &  (~ n895) ) ;
 assign n63 = ( PV246_0_  &  n379 ) | ( (~ PV246_0_)  &  (~ n379) ) ;
 assign n64 = ( (~ PV802_0_) ) | ( (~ n265) ) ;
 assign n65 = ( PV247_0_  &  n461 ) | ( (~ PV247_0_)  &  (~ n461) ) ;
 assign n69 = ( PV214_0_  &  n961 ) | ( n239  &  n961 ) | ( (~ n958)  &  n961 ) ;
 assign n66 = ( n408  &  (~ n725)  &  (~ n959) ) ;
 assign n68 = ( n32 ) | ( n239 ) | ( PV214_0_ ) ;
 assign n70 = ( PV45_0_  &  PV41_0_ ) | ( (~ PV45_0_)  &  (~ PV41_0_) ) ;
 assign n73 = ( PV174_0_ ) | ( n229 ) ;
 assign n71 = ( PV278_0_  &  (~ PV277_0_) ) | ( PV278_0_  &  n73 ) ;
 assign n75 = ( PV257_2_  &  n854 ) ;
 assign n74 = ( n75  &  PV257_1_ ) ;
 assign n76 = ( PV261_0_  &  PV165_7_  &  PV165_6_  &  PV165_2_  &  PV165_1_  &  PV165_0_  &  (~ n251)  &  (~ n922) ) ;
 assign n78 = ( (~ PV13_0_)  &  PV10_0_ ) ;
 assign n82 = ( PV149_2_  &  PV149_0_  &  (~ n122) ) | ( PV149_1_  &  PV149_0_  &  (~ n122) ) ;
 assign n84 = ( n230  &  n247 ) | ( n230  &  n248 ) ;
 assign n85 = ( (~ PV165_6_)  &  n141 ) ;
 assign n87 = ( n37  &  n354 ) | ( (~ n37)  &  (~ n354) ) ;
 assign n88 = ( n36  &  n355 ) | ( (~ n36)  &  (~ n355) ) ;
 assign n89 = ( (~ n641)  &  n656 ) | ( (~ n641)  &  n974 ) | ( (~ n656)  &  n974 ) ;
 assign n90 = ( (~ n38)  &  n351 ) | ( n38  &  (~ n351) ) ;
 assign n86 = ( n87  &  n88  &  PV288_2_  &  n89  &  n90 ) ;
 assign n92 = ( (~ n37)  &  n350 ) | ( n37  &  (~ n350) ) ;
 assign n93 = ( (~ PV288_3_) ) | ( (~ PV288_2_) ) ;
 assign n95 = ( (~ n36)  &  n346 ) | ( n36  &  (~ n346) ) ;
 assign n91 = ( n90 ) | ( n92 ) | ( n93 ) | ( n95 ) | ( (~ n973) ) ;
 assign n97 = ( (~ n37)  &  n666 ) | ( n37  &  (~ n666) ) ;
 assign n98 = ( (~ n36)  &  n655 ) | ( n36  &  (~ n655) ) ;
 assign n100 = ( (~ n641)  &  n657 ) | ( (~ n641)  &  n974 ) | ( (~ n657)  &  n974 ) ;
 assign n96 = ( n90  &  (~ n93)  &  n97  &  n98  &  n100 ) ;
 assign n102 = ( n37  &  n336 ) | ( (~ n37)  &  (~ n336) ) ;
 assign n103 = ( n36  &  n337 ) | ( (~ n36)  &  (~ n337) ) ;
 assign n104 = ( (~ n641)  &  n669 ) | ( (~ n641)  &  n974 ) | ( (~ n669)  &  n974 ) ;
 assign n105 = ( (~ n38)  &  n333 ) | ( n38  &  (~ n333) ) ;
 assign n101 = ( n102  &  n103  &  PV288_0_  &  n104  &  n105 ) ;
 assign n107 = ( (~ n37)  &  n332 ) | ( n37  &  (~ n332) ) ;
 assign n110 = ( (~ n36)  &  n326 ) | ( n36  &  (~ n326) ) ;
 assign n106 = ( n105 ) | ( n107 ) | ( n110 ) | ( (~ n112) ) | ( (~ n978) ) ;
 assign n112 = ( PV288_1_  &  PV288_0_ ) ;
 assign n113 = ( n37  &  n327 ) | ( (~ n37)  &  (~ n327) ) ;
 assign n114 = ( n169  &  (~ n641) ) | ( (~ n169)  &  n974 ) | ( (~ n641)  &  n974 ) ;
 assign n115 = ( (~ n36)  &  n662 ) | ( n36  &  (~ n662) ) ;
 assign n111 = ( n112  &  n113  &  n105  &  n114  &  n115 ) ;
 assign n117 = ( (~ n84)  &  n85 ) ;
 assign n121 = ( n588  &  n586  &  n522  &  n721  &  n567  &  n722 ) ;
 assign n120 = ( PV260_0_ ) | ( PV259_0_ ) | ( (~ PV258_0_) ) | ( PV59_0_ ) ;
 assign n119 = ( n121  &  n120 ) | ( n121  &  (~ n122) ) ;
 assign n122 = ( PV262_0_ ) | ( n76 ) ;
 assign n124 = ( (~ PV57_0_)  &  n224 ) | ( PV57_0_  &  n624 ) | ( n224  &  n624 ) ;
 assign n129 = ( PV59_0_  &  (~ PV1719)  &  n497  &  n498  &  n499  &  n501 ) ;
 assign n130 = ( (~ PV213_5_)  &  (~ PV165_7_) ) | ( (~ PV213_5_)  &  n510 ) | ( (~ PV165_7_)  &  n511 ) | ( n510  &  n511 ) ;
 assign n131 = ( (~ PV213_4_)  &  (~ PV165_6_) ) | ( (~ PV213_4_)  &  n510 ) | ( (~ PV165_6_)  &  n511 ) | ( n510  &  n511 ) ;
 assign n132 = ( (~ PV213_3_)  &  (~ PV165_5_) ) | ( (~ PV213_3_)  &  n510 ) | ( (~ PV165_5_)  &  n511 ) | ( n510  &  n511 ) ;
 assign n133 = ( (~ PV213_2_)  &  (~ PV165_4_) ) | ( (~ PV213_2_)  &  n510 ) | ( (~ PV165_4_)  &  n511 ) | ( n510  &  n511 ) ;
 assign n134 = ( (~ PV213_1_)  &  (~ PV165_3_) ) | ( (~ PV213_1_)  &  n510 ) | ( (~ PV165_3_)  &  n511 ) | ( n510  &  n511 ) ;
 assign n135 = ( (~ PV782)  &  n617 ) | ( n617  &  n621 ) | ( (~ PV782)  &  (~ n963) ) | ( n621  &  (~ n963) ) ;
 assign n136 = ( PV149_3_  &  (~ n267) ) ;
 assign n142 = ( n385  &  n261  &  PV65_0_ ) ;
 assign n141 = ( (~ PV165_5_)  &  (~ PV165_4_)  &  PV165_3_  &  PV70_0_ ) ;
 assign n145 = ( (~ PV60_0_)  &  (~ PV56_0_) ) ;
 assign n143 = ( (~ PV59_0_)  &  n145 ) ;
 assign n147 = ( (~ PV277_0_)  &  n522 ) | ( (~ PV14_0_)  &  n522 ) | ( (~ n73)  &  n522 ) ;
 assign n148 = ( PV258_0_  &  n523 ) | ( (~ PV258_0_)  &  (~ n523) ) ;
 assign n149 = ( PV259_0_  &  n986 ) | ( (~ PV259_0_)  &  (~ n986) ) ;
 assign n150 = ( PV260_0_  &  n987 ) | ( (~ PV260_0_)  &  (~ n987) ) ;
 assign n151 = ( n248 ) | ( n255 ) ;
 assign n155 = ( (~ n390) ) | ( n394 ) | ( (~ n396) ) ;
 assign n153 = ( (~ n673)  &  n674 ) | ( n673  &  (~ n674) ) ;
 assign n154 = ( (~ n675)  &  n676 ) | ( n675  &  (~ n676) ) ;
 assign n152 = ( n155  &  n153 ) | ( n155  &  n154 ) ;
 assign n156 = ( (~ PV15_0_)  &  (~ n152) ) | ( (~ PV802_0_)  &  (~ n152)  &  (~ n267) ) ;
 assign n157 = ( PV69_0_ ) | ( PV68_0_ ) | ( PV70_0_ ) | ( PV66_0_ ) ;
 assign n158 = ( PV66_0_  &  PV215_0_ ) ;
 assign n159 = ( (~ PV216_0_)  &  (~ n1025) ) | ( PV214_0_  &  (~ n1025) ) ;
 assign n160 = ( n531  &  n532  &  n529 ) | ( n531  &  n532  &  (~ n943) ) ;
 assign n163 = ( (~ n267) ) | ( (~ n563) ) ;
 assign n162 = ( PV56_0_  &  n163  &  PV171_0_ ) ;
 assign n164 = ( PV63_0_  &  (~ n25) ) | ( PV60_0_  &  (~ n25) ) ;
 assign n166 = ( PV302_0_  &  n534 ) | ( (~ PV292_0_)  &  n534 ) ;
 assign n167 = ( n538  &  n70  &  n535 ) | ( n538  &  n70  &  n224 ) ;
 assign n170 = ( n401  &  PV32_0_ ) | ( n402  &  PV32_0_ ) | ( n401  &  n169 ) | ( n402  &  n169 ) ;
 assign n169 = ( n322  &  n657 ) | ( (~ n322)  &  (~ n657) ) ;
 assign n168 = ( n170  &  (~ n1022) ) | ( PV32_0_  &  n169  &  (~ n1022) ) ;
 assign n172 = ( (~ PV149_7_)  &  (~ n168)  &  n540 ) | ( (~ n168)  &  n393  &  n540 ) ;
 assign n176 = ( n76 ) | ( (~ n121) ) | ( n180 ) ;
 assign n173 = ( n176 ) | ( (~ n224) ) | ( (~ n699) ) ;
 assign n177 = ( PV802_0_ ) | ( PV289_0_ ) | ( n276 ) ;
 assign n178 = ( PV289_0_ ) | ( (~ n173) ) | ( n234 ) | ( (~ n259) ) | ( (~ n732) ) ;
 assign n179 = ( PV289_0_  &  n962 ) | ( (~ PV1741_0_)  &  n962 ) | ( n176  &  n962 ) ;
 assign n180 = ( n120  &  PV14_0_  &  PV262_0_ ) ;
 assign n181 = ( (~ PV165_7_)  &  (~ PV100_5_) ) | ( (~ PV100_5_)  &  n544 ) | ( (~ PV165_7_)  &  n545 ) | ( n544  &  n545 ) ;
 assign n182 = ( (~ PV165_6_)  &  (~ PV100_4_) ) | ( (~ PV100_4_)  &  n544 ) | ( (~ PV165_6_)  &  n545 ) | ( n544  &  n545 ) ;
 assign n183 = ( (~ PV165_5_)  &  (~ PV100_3_) ) | ( (~ PV100_3_)  &  n544 ) | ( (~ PV165_5_)  &  n545 ) | ( n544  &  n545 ) ;
 assign n184 = ( (~ PV165_4_)  &  (~ PV100_2_) ) | ( (~ PV100_2_)  &  n544 ) | ( (~ PV165_4_)  &  n545 ) | ( n544  &  n545 ) ;
 assign n185 = ( (~ PV165_3_)  &  (~ PV100_1_) ) | ( (~ PV100_1_)  &  n544 ) | ( (~ PV165_3_)  &  n545 ) | ( n544  &  n545 ) ;
 assign n186 = ( (~ PV1719)  &  n386 ) | ( n278  &  n386 ) | ( n386  &  (~ n946) ) ;
 assign n187 = ( PV1536_0_  &  n554 ) | ( (~ n265)  &  n554 ) | ( n554  &  n553 ) ;
 assign n191 = ( PV62_0_  &  n32  &  (~ n223) ) ;
 assign n193 = ( n267  &  n268  &  (~ n966) ) ;
 assign n195 = ( PV16_0_ ) | ( (~ PV15_0_) ) ;
 assign n196 = ( (~ PV16_0_) ) | ( PV15_0_ ) ;
 assign n194 = ( n195  &  n196 ) ;
 assign n197 = ( (~ PV101_0_)  &  n556 ) | ( (~ PV14_0_)  &  n556 ) | ( n556  &  n555 ) ;
 assign n198 = ( (~ PV262_0_)  &  PV261_0_ ) | ( PV261_0_  &  n180 ) | ( PV261_0_  &  (~ n1024) ) ;
 assign n199 = ( PV268_0_  &  n831 ) ;
 assign n200 = ( (~ PV16_0_)  &  (~ n152)  &  n558 ) | ( (~ PV15_0_)  &  (~ n152)  &  n558 ) ;
 assign n201 = ( (~ PV108_1_)  &  n73 ) | ( (~ PV108_1_)  &  (~ n152) ) | ( n73  &  n559 ) | ( (~ n152)  &  n559 ) ;
 assign n202 = ( (~ PV108_2_)  &  n229 ) | ( n229  &  n559 ) | ( (~ PV108_2_)  &  (~ n731) ) | ( n559  &  (~ n731) ) ;
 assign n203 = ( (~ PV108_3_)  &  n563 ) | ( n559  &  n563 ) | ( (~ PV108_3_)  &  (~ n731) ) | ( n559  &  (~ n731) ) ;
 assign n204 = ( (~ PV108_4_)  &  n195 ) | ( n195  &  n559 ) ;
 assign n205 = ( (~ PV108_5_)  &  n196 ) | ( n196  &  n555 ) ;
 assign n206 = ( (~ PV213_5_)  &  n568 ) | ( n568  &  n567 ) ;
 assign n207 = ( (~ PV132_7_)  &  (~ PV118_5_) ) | ( (~ PV132_7_)  &  n586 ) | ( (~ PV118_5_)  &  n588 ) | ( n586  &  n588 ) ;
 assign n208 = ( (~ PV132_6_)  &  (~ PV118_4_) ) | ( (~ PV132_6_)  &  n586 ) | ( (~ PV118_4_)  &  n588 ) | ( n586  &  n588 ) ;
 assign n209 = ( (~ PV132_5_)  &  (~ PV118_3_) ) | ( (~ PV132_5_)  &  n586 ) | ( (~ PV118_3_)  &  n588 ) | ( n586  &  n588 ) ;
 assign n210 = ( (~ PV132_4_)  &  (~ PV118_2_) ) | ( (~ PV132_4_)  &  n586 ) | ( (~ PV118_2_)  &  n588 ) | ( n586  &  n588 ) ;
 assign n211 = ( (~ PV132_3_)  &  (~ PV118_1_) ) | ( (~ PV132_3_)  &  n586 ) | ( (~ PV118_1_)  &  n588 ) | ( n586  &  n588 ) ;
 assign n212 = ( (~ PV132_2_)  &  (~ PV118_0_) ) | ( (~ PV132_2_)  &  n586 ) | ( (~ PV118_0_)  &  n588 ) | ( n586  &  n588 ) ;
 assign n213 = ( (~ PV132_0_)  &  (~ PV108_5_) ) | ( (~ PV108_5_)  &  n588 ) | ( (~ PV132_0_)  &  n600 ) | ( n588  &  n600 ) ;
 assign n214 = ( (~ PV134_1_)  &  n604 ) | ( n604  &  n603 ) ;
 assign n215 = ( (~ n36) ) | ( (~ n37) ) | ( (~ n38) ) | ( n639 ) | ( n641 ) ;
 assign n216 = ( n660 ) | ( n872 ) | ( n875 ) | ( n642 ) | ( n357 ) | ( n870 ) ;
 assign n218 = ( n344  &  n106  &  n833  &  n5 ) ;
 assign n219 = ( n4  &  (~ n101)  &  (~ n111)  &  n832 ) ;
 assign n222 = ( (~ n37) ) | ( n38 ) | ( n762 ) ;
 assign n223 = ( n718 ) | ( n256 ) ;
 assign n224 = ( n717 ) | ( n718 ) ;
 assign n225 = ( n715 ) | ( n718 ) ;
 assign n226 = ( n777  &  n964 ) ;
 assign n229 = ( (~ PV149_4_) ) | ( PV149_3_ ) | ( n707 ) ;
 assign n230 = ( n247 ) | ( n715 ) ;
 assign n228 = ( PV33_0_  &  PV289_0_  &  n229  &  n230 ) ;
 assign n231 = ( n71  &  n265 ) ;
 assign n234 = ( (~ PV290_0_)  &  PV165_7_  &  n239 ) ;
 assign n235 = ( (~ PV1741_0_)  &  (~ n259)  &  n276 ) ;
 assign n236 = ( n263  &  n9 ) | ( n263  &  n278 ) ;
 assign n238 = ( (~ PV274_0_)  &  (~ PV271_0_) ) | ( (~ PV271_0_)  &  PV202_0_ ) ;
 assign n239 = ( (~ PV165_2_)  &  PV165_1_  &  PV165_0_ ) ;
 assign n240 = ( (~ n243)  &  (~ n381)  &  n384  &  n531 ) ;
 assign n242 = ( n22 ) | ( (~ n937) ) | ( (~ n1005) ) ;
 assign n243 = ( PV56_0_  &  (~ n499) ) | ( PV56_0_  &  (~ n23)  &  (~ n625) ) ;
 assign n247 = ( (~ PV149_5_) ) | ( (~ PV149_4_) ) ;
 assign n248 = ( (~ PV149_6_) ) | ( n711 ) ;
 assign n250 = ( n229  &  n563 ) ;
 assign n249 = ( n250  &  PV802_0_ ) | ( n250  &  PV55_0_ ) | ( n250  &  n84 ) ;
 assign n253 = ( PV292_0_ ) | ( PV291_0_ ) | ( (~ PV169_0_) ) | ( n85 ) | ( n249 ) ;
 assign n251 = ( PV204_0_  &  (~ PV70_0_) ) | ( PV204_0_  &  n253 ) ;
 assign n257 = ( (~ PV149_3_) ) | ( (~ n600) ) | ( n710 ) | ( n740 ) | ( n839 ) ;
 assign n256 = ( PV149_6_ ) | ( n714 ) ;
 assign n255 = ( PV149_5_ ) | ( PV149_4_ ) ;
 assign n254 = ( n257  &  n256 ) | ( n257  &  n247  &  n255 ) ;
 assign n258 = ( n225  &  n224 ) ;
 assign n262 = ( (~ PV62_0_)  &  (~ PV56_0_) ) | ( (~ PV62_0_)  &  n119 ) | ( (~ PV56_0_)  &  n258 ) | ( n119  &  n258 ) ;
 assign n261 = ( n248 ) | ( n718 ) ;
 assign n259 = ( (~ PV65_0_)  &  n262 ) | ( n262  &  n261 ) ;
 assign n265 = ( (~ n289) ) | ( n725 ) ;
 assign n263 = ( PV241_0_  &  n265 ) | ( n265  &  (~ n289) ) ;
 assign n267 = ( (~ PV149_2_) ) | ( PV149_1_ ) | ( PV149_0_ ) ;
 assign n268 = ( n32  &  (~ n239) ) ;
 assign n269 = ( n32  &  n267  &  (~ n966) ) ;
 assign n271 = ( (~ PV242_0_) ) | ( (~ PV134_1_) ) | ( (~ PV134_0_) ) ;
 assign n270 = ( (~ PV261_0_)  &  n271 ) | ( (~ n263)  &  n271 ) ;
 assign n274 = ( (~ PV802_0_)  &  (~ n71)  &  n265 ) ;
 assign n272 = ( PV242_0_  &  (~ PV56_0_)  &  n274 ) | ( PV242_0_  &  n274  &  (~ n725) ) ;
 assign n276 = ( PV165_7_ ) | ( (~ n239) ) ;
 assign n278 = ( PV302_0_ ) | ( n234 ) | ( (~ n276) ) | ( (~ n732) ) ;
 assign n279 = ( (~ PV174_0_)  &  (~ n73) ) | ( (~ PV174_0_)  &  n163 ) | ( (~ PV174_0_)  &  (~ n289) ) ;
 assign n283 = ( (~ PV149_3_) ) | ( n707 ) ;
 assign n281 = ( (~ PV59_0_)  &  (~ n71) ) ;
 assign n280 = ( (~ n279)  &  n283 ) | ( (~ PV60_0_)  &  (~ n279)  &  n281 ) ;
 assign n287 = ( (~ n18)  &  (~ n382)  &  n409 ) ;
 assign n285 = ( n73  &  (~ n136)  &  n287 ) | ( n71  &  (~ n136)  &  n287 ) ;
 assign n289 = ( PV149_4_ ) | ( PV149_3_ ) | ( n707 ) ;
 assign n288 = ( (~ PV56_0_)  &  PV53_0_  &  (~ n122)  &  n283  &  n289 ) ;
 assign n293 = ( PV56_0_ ) | ( PV57_0_ ) | ( PV53_0_ ) ;
 assign n291 = ( n385  &  n410 ) ;
 assign n290 = ( n145  &  (~ n285)  &  n293 ) | ( (~ n285)  &  n293  &  n291 ) ;
 assign n295 = ( (~ n25) ) | ( n288 ) | ( n290 ) ;
 assign n294 = ( (~ PV60_0_)  &  n295 ) | ( n73  &  (~ n136)  &  n295 ) ;
 assign n298 = ( (~ PV223_1_)  &  (~ PV32_1_) ) | ( (~ PV223_1_)  &  (~ n294) ) | ( (~ PV32_1_)  &  n754 ) | ( (~ n294)  &  n754 ) ;
 assign n296 = ( n163 ) | ( n752 ) ;
 assign n300 = ( (~ PV223_2_)  &  (~ PV32_2_) ) | ( (~ PV223_2_)  &  (~ n294) ) | ( (~ PV32_2_)  &  n754 ) | ( (~ n294)  &  n754 ) ;
 assign n302 = ( (~ PV223_3_)  &  (~ PV32_3_) ) | ( (~ PV223_3_)  &  (~ n294) ) | ( (~ PV32_3_)  &  n754 ) | ( (~ n294)  &  n754 ) ;
 assign n304 = ( (~ PV223_0_)  &  (~ PV32_0_) ) | ( (~ PV223_0_)  &  (~ n294) ) | ( (~ PV32_0_)  &  n754 ) | ( (~ n294)  &  n754 ) ;
 assign n307 = ( (~ PV288_7_) ) | ( PV288_6_ ) ;
 assign n305 = ( PV288_7_  &  n307 ) | ( (~ PV288_6_)  &  n307 ) ;
 assign n308 = ( n307  &  (~ n320) ) ;
 assign n313 = ( (~ n351) ) | ( n665 ) | ( (~ n666) ) ;
 assign n312 = ( PV288_1_ ) | ( (~ PV288_0_) ) ;
 assign n310 = ( n313  &  n312 ) | ( n313  &  (~ n666) ) ;
 assign n317 = ( n315 ) | ( (~ n632) ) | ( n653 ) ;
 assign n315 = ( (~ n308)  &  n633 ) | ( n308  &  (~ n633) ) ;
 assign n314 = ( n317  &  n315 ) | ( n317  &  (~ n765) ) ;
 assign n320 = ( (~ PV288_5_) ) | ( PV288_4_ ) ;
 assign n321 = ( PV288_5_ ) | ( (~ PV288_4_) ) ;
 assign n319 = ( (~ n305) ) | ( n320  &  n321 ) ;
 assign n322 = ( (~ n655) ) | ( (~ n112)  &  n310 ) ;
 assign n324 = ( (~ n630) ) | ( n93  &  n314 ) ;
 assign n330 = ( (~ n327) ) | ( n333 ) | ( n662 ) ;
 assign n327 = ( (~ n664)  &  n666 ) | ( n664  &  (~ n666) ) ;
 assign n326 = ( n330  &  (~ n662) ) | ( n330  &  n327  &  (~ n333) ) ;
 assign n332 = ( n327  &  n333 ) | ( (~ n327)  &  (~ n333) ) ;
 assign n333 = ( n351  &  n665 ) | ( (~ n351)  &  (~ n665) ) ;
 assign n331 = ( n326  &  (~ n670) ) | ( n332  &  n333  &  (~ n670) ) ;
 assign n337 = ( n312  &  n331 ) | ( (~ n312)  &  (~ n662) ) | ( n331  &  (~ n662) ) ;
 assign n336 = ( (~ n312)  &  n327 ) | ( n312  &  n878 ) | ( n327  &  n878 ) ;
 assign n335 = ( n337  &  (~ n1016) ) | ( (~ n333)  &  n336  &  (~ n1016) ) ;
 assign n339 = ( (~ PV288_1_)  &  (~ PV288_0_) ) ;
 assign n344 = ( n672 ) | ( n883 ) | ( n886 ) | ( n642 ) | ( n339 ) | ( n881 ) ;
 assign n342 = ( (~ n101)  &  n106  &  (~ n111)  &  (~ n122)  &  n344 ) ;
 assign n348 = ( n351 ) | ( n666 ) | ( n655 ) ;
 assign n346 = ( n348  &  (~ n655) ) | ( n348  &  (~ n351)  &  (~ n666) ) ;
 assign n350 = ( (~ n351)  &  n666 ) | ( n351  &  (~ n666) ) ;
 assign n351 = ( n632  &  n653 ) | ( (~ n632)  &  (~ n653) ) ;
 assign n349 = ( n346  &  (~ n658) ) | ( n350  &  n351  &  (~ n658) ) ;
 assign n355 = ( n349  &  (~ n655) ) | ( (~ n655)  &  n765 ) | ( n349  &  (~ n765) ) ;
 assign n354 = ( (~ n666)  &  n765 ) | ( (~ n666)  &  n976 ) | ( (~ n765)  &  n976 ) ;
 assign n353 = ( n355  &  (~ n869) ) | ( (~ n351)  &  n354  &  (~ n869) ) ;
 assign n357 = ( (~ PV288_3_)  &  (~ PV288_2_) ) ;
 assign n360 = ( (~ n86)  &  n91  &  (~ n96)  &  (~ n122)  &  n216 ) ;
 assign n361 = ( (~ PV288_5_)  &  (~ PV288_4_) ) ;
 assign n364 = ( PV288_7_  &  PV288_6_  &  (~ n1020) ) ;
 assign n366 = ( (~ n4)  &  (~ n764) ) | ( n122  &  (~ n764) ) | ( (~ n764)  &  (~ n925) ) ;
 assign n370 = ( (~ PV239_3_)  &  (~ PV199_3_) ) | ( (~ PV239_3_)  &  n296 ) | ( (~ PV199_3_)  &  n754 ) | ( n296  &  n754 ) ;
 assign n371 = ( (~ PV88_0_)  &  (~ PV32_10_) ) | ( (~ PV32_10_)  &  (~ n294) ) | ( (~ PV88_0_)  &  n766 ) | ( (~ n294)  &  n766 ) ;
 assign n372 = ( (~ PV239_2_)  &  (~ PV199_2_) ) | ( (~ PV239_2_)  &  n296 ) | ( (~ PV199_2_)  &  n754 ) | ( n296  &  n754 ) ;
 assign n373 = ( (~ PV84_5_)  &  (~ PV32_9_) ) | ( (~ PV32_9_)  &  (~ n294) ) | ( (~ PV84_5_)  &  n766 ) | ( (~ n294)  &  n766 ) ;
 assign n374 = ( (~ PV239_4_)  &  (~ PV199_4_) ) | ( (~ PV239_4_)  &  n296 ) | ( (~ PV199_4_)  &  n754 ) | ( n296  &  n754 ) ;
 assign n375 = ( (~ PV88_1_)  &  (~ PV32_11_) ) | ( (~ PV32_11_)  &  (~ n294) ) | ( (~ PV88_1_)  &  n766 ) | ( (~ n294)  &  n766 ) ;
 assign n380 = ( n11  &  n694 ) | ( n12  &  n694 ) | ( n694  &  (~ n928) ) ;
 assign n379 = ( (~ PV245_0_) ) | ( (~ PV244_0_) ) | ( (~ PV243_0_) ) ;
 assign n376 = ( (~ PV247_0_)  &  n380 ) | ( (~ PV246_0_)  &  n380 ) | ( n380  &  n379 ) ;
 assign n382 = ( (~ PV149_3_)  &  n247  &  (~ n267) ) ;
 assign n381 = ( PV59_0_  &  n382 ) | ( PV59_0_  &  (~ n964) ) ;
 assign n385 = ( (~ n18) ) | ( (~ n23) ) ;
 assign n384 = ( (~ PV62_0_) ) | ( n385 ) ;
 assign n387 = ( (~ PV802_0_) ) | ( (~ n136) ) ;
 assign n386 = ( n387  &  n71 ) | ( n387  &  n64 ) ;
 assign n393 = ( (~ PV802_0_) ) | ( n267 ) ;
 assign n392 = ( PV174_0_ ) | ( n563 ) ;
 assign n390 = ( (~ PV802_0_)  &  n393 ) | ( n393  &  n392 ) ;
 assign n394 = ( PV56_0_  &  (~ n25) ) | ( PV56_0_  &  (~ n224) ) | ( PV56_0_  &  (~ n721) ) ;
 assign n396 = ( (~ PV802_0_) ) | ( n73 ) ;
 assign n395 = ( (~ PV802_0_)  &  n396 ) | ( n392  &  n396 ) ;
 assign n397 = ( PV56_0_  &  (~ n224) ) | ( PV56_0_  &  (~ n506) ) | ( PV56_0_  &  (~ n699) ) ;
 assign n399 = ( PV32_3_  &  PV32_2_  &  (~ n333) ) | ( PV32_3_  &  n327  &  (~ n333) ) ;
 assign n400 = ( n327  &  PV32_2_ ) ;
 assign n401 = ( PV32_1_  &  n399 ) | ( PV32_1_  &  n400 ) | ( n399  &  (~ n662) ) | ( n400  &  (~ n662) ) ;
 assign n402 = ( PV32_1_  &  (~ n662) ) ;
 assign n403 = ( (~ n64)  &  n71 ) | ( PV59_0_  &  n71  &  n263 ) ;
 assign n405 = ( (~ PV270_0_)  &  (~ PV56_0_)  &  (~ n403) ) | ( (~ PV270_0_)  &  n25  &  (~ n403) ) ;
 assign n409 = ( (~ PV149_3_) ) | ( n392 ) ;
 assign n408 = ( n23  &  (~ n136) ) | ( (~ n136)  &  n409 ) ;
 assign n411 = ( (~ PV56_0_)  &  n939 ) | ( n66  &  n699  &  n939 ) ;
 assign n410 = ( (~ n23) ) | ( n409 ) ;
 assign n414 = ( n788 ) | ( n396 ) ;
 assign n416 = ( PV199_4_  &  PV199_3_ ) | ( (~ PV199_4_)  &  (~ PV199_3_) ) ;
 assign n419 = ( (~ PV234_0_)  &  (~ PV194_0_) ) | ( (~ PV194_0_)  &  n463 ) | ( (~ PV234_0_)  &  n474 ) | ( n463  &  n474 ) ;
 assign n420 = ( (~ PV32_2_)  &  n940 ) | ( n439  &  n940 ) ;
 assign n418 = ( (~ n122) ) | ( (~ n280) ) | ( n794 ) ;
 assign n417 = ( (~ PV257_7_)  &  n419  &  n420 ) | ( n419  &  n420  &  n418 ) ;
 assign n423 = ( PV199_2_  &  n678 ) | ( (~ PV199_2_)  &  (~ n678) ) ;
 assign n425 = ( (~ PV32_11_)  &  (~ PV32_8_) ) | ( (~ PV32_11_)  &  n766 ) | ( (~ PV32_8_)  &  n797 ) | ( n766  &  n797 ) ;
 assign n426 = ( (~ PV239_1_)  &  (~ PV199_1_) ) | ( (~ PV239_1_)  &  n296 ) | ( (~ PV199_1_)  &  n754 ) | ( n296  &  n754 ) ;
 assign n427 = ( PV199_1_  &  n429 ) | ( (~ PV199_1_)  &  (~ n429) ) ;
 assign n429 = ( n678  &  PV199_2_ ) ;
 assign n428 = ( PV199_1_  &  n429 ) ;
 assign n431 = ( (~ PV32_10_)  &  (~ PV32_7_) ) | ( (~ PV32_10_)  &  n766 ) | ( (~ PV32_7_)  &  n797 ) | ( n766  &  n797 ) ;
 assign n432 = ( (~ PV239_0_)  &  (~ PV199_0_) ) | ( (~ PV239_0_)  &  n296 ) | ( (~ PV199_0_)  &  n754 ) | ( n296  &  n754 ) ;
 assign n433 = ( PV199_0_  &  n428 ) | ( (~ PV199_0_)  &  (~ n428) ) ;
 assign n435 = ( (~ PV32_9_)  &  (~ PV32_6_) ) | ( (~ PV32_9_)  &  n766 ) | ( (~ PV32_6_)  &  n797 ) | ( n766  &  n797 ) ;
 assign n436 = ( (~ PV234_4_)  &  (~ PV194_4_) ) | ( (~ PV234_4_)  &  n296 ) | ( (~ PV194_4_)  &  n754 ) | ( n296  &  n754 ) ;
 assign n437 = ( PV194_4_  &  n682 ) | ( (~ PV194_4_)  &  (~ n682) ) ;
 assign n441 = ( (~ PV149_7_)  &  (~ PV32_8_) ) | ( (~ PV149_7_)  &  n792 ) | ( (~ PV32_8_)  &  n795 ) | ( n792  &  n795 ) ;
 assign n442 = ( (~ PV234_3_)  &  (~ PV194_3_) ) | ( (~ PV194_3_)  &  n463 ) | ( (~ PV234_3_)  &  n474 ) | ( n463  &  n474 ) ;
 assign n439 = ( n143 ) | ( n750 ) ;
 assign n438 = ( (~ PV32_5_)  &  n441  &  n442 ) | ( n441  &  n442  &  n439 ) ;
 assign n444 = ( (~ PV149_7_)  &  n684 ) | ( (~ PV149_7_)  &  (~ n790) ) | ( n684  &  n801 ) | ( (~ n790)  &  n801 ) ;
 assign n447 = ( (~ PV149_6_)  &  (~ PV32_7_) ) | ( (~ PV149_6_)  &  n792 ) | ( (~ PV32_7_)  &  n795 ) | ( n792  &  n795 ) ;
 assign n448 = ( (~ PV234_2_)  &  (~ PV194_2_) ) | ( (~ PV194_2_)  &  n463 ) | ( (~ PV234_2_)  &  n474 ) | ( n463  &  n474 ) ;
 assign n445 = ( (~ PV32_4_)  &  n447  &  n448 ) | ( n439  &  n447  &  n448 ) ;
 assign n450 = ( (~ PV149_6_)  &  n687 ) | ( (~ PV149_6_)  &  (~ n790) ) | ( n687  &  n801 ) | ( (~ n790)  &  n801 ) ;
 assign n453 = ( (~ PV149_5_)  &  (~ PV32_6_) ) | ( (~ PV149_5_)  &  n792 ) | ( (~ PV32_6_)  &  n795 ) | ( n792  &  n795 ) ;
 assign n454 = ( (~ PV234_1_)  &  (~ PV194_1_) ) | ( (~ PV194_1_)  &  n463 ) | ( (~ PV234_1_)  &  n474 ) | ( n463  &  n474 ) ;
 assign n451 = ( (~ PV32_3_)  &  n453  &  n454 ) | ( n439  &  n453  &  n454 ) ;
 assign n456 = ( (~ PV149_5_)  &  n690 ) | ( (~ PV149_5_)  &  (~ n790) ) | ( n690  &  n801 ) | ( (~ n790)  &  n801 ) ;
 assign n457 = ( (~ PV149_4_)  &  n693 ) | ( (~ PV149_4_)  &  (~ n790) ) | ( n693  &  n801 ) | ( (~ n790)  &  n801 ) ;
 assign n460 = ( PV243_0_ ) | ( (~ n64) ) ;
 assign n461 = ( (~ PV246_0_) ) | ( n379 ) ;
 assign n465 = ( (~ PV32_4_)  &  (~ PV32_1_) ) | ( (~ PV32_4_)  &  n439 ) | ( (~ PV32_1_)  &  n792 ) | ( n439  &  n792 ) ;
 assign n466 = ( (~ PV257_6_)  &  (~ PV189_5_) ) | ( (~ PV189_5_)  &  n418 ) | ( (~ PV257_6_)  &  n474 ) | ( n418  &  n474 ) ;
 assign n463 = ( n265 ) | ( (~ n748) ) ;
 assign n462 = ( (~ PV229_5_)  &  n465  &  n466 ) | ( n465  &  n466  &  n463 ) ;
 assign n470 = ( (~ PV32_3_)  &  (~ PV32_0_) ) | ( (~ PV32_3_)  &  n439 ) | ( (~ PV32_0_)  &  n792 ) | ( n439  &  n792 ) ;
 assign n471 = ( (~ PV257_5_)  &  (~ PV189_4_) ) | ( (~ PV189_4_)  &  n418 ) | ( (~ PV257_5_)  &  n474 ) | ( n418  &  n474 ) ;
 assign n468 = ( (~ PV229_4_)  &  n470  &  n471 ) | ( n463  &  n470  &  n471 ) ;
 assign n476 = ( (~ PV229_3_)  &  n439 ) | ( n439  &  n463 ) ;
 assign n477 = ( (~ PV257_4_)  &  (~ PV32_2_) ) | ( (~ PV32_2_)  &  n418 ) | ( (~ PV257_4_)  &  n750 ) | ( n418  &  n750 ) ;
 assign n474 = ( n163 ) | ( (~ n748) ) ;
 assign n473 = ( (~ PV189_3_)  &  n476  &  n477 ) | ( n476  &  n477  &  n474 ) ;
 assign n481 = ( (~ PV229_2_)  &  n439 ) | ( n439  &  n463 ) ;
 assign n482 = ( (~ PV257_3_)  &  (~ PV32_1_) ) | ( (~ PV32_1_)  &  n418 ) | ( (~ PV257_3_)  &  n750 ) | ( n418  &  n750 ) ;
 assign n479 = ( (~ PV189_2_)  &  n481  &  n482 ) | ( n474  &  n481  &  n482 ) ;
 assign n486 = ( (~ PV229_1_)  &  n439 ) | ( n439  &  n463 ) ;
 assign n487 = ( (~ PV257_2_)  &  (~ PV32_0_) ) | ( (~ PV32_0_)  &  n418 ) | ( (~ PV257_2_)  &  n750 ) | ( n418  &  n750 ) ;
 assign n484 = ( (~ PV189_1_)  &  n486  &  n487 ) | ( n474  &  n486  &  n487 ) ;
 assign n490 = ( (~ PV257_1_)  &  n766 ) | ( n766  &  n815 ) ;
 assign n491 = ( (~ PV229_0_)  &  (~ PV189_0_) ) | ( (~ PV229_0_)  &  n296 ) | ( (~ PV189_0_)  &  n754 ) | ( n296  &  n754 ) ;
 assign n492 = ( (~ PV257_0_)  &  n797 ) | ( n797  &  n815 ) ;
 assign n493 = ( (~ PV223_5_)  &  (~ PV183_5_) ) | ( (~ PV223_5_)  &  n296 ) | ( (~ PV183_5_)  &  n754 ) | ( n296  &  n754 ) ;
 assign n495 = ( (~ PV223_4_)  &  (~ PV183_4_) ) | ( (~ PV223_4_)  &  n296 ) | ( (~ PV183_4_)  &  n754 ) | ( n296  &  n754 ) ;
 assign n496 = ( (~ PV257_6_)  &  (~ PV32_4_) ) | ( (~ PV257_6_)  &  (~ n294) ) | ( (~ PV32_4_)  &  n815 ) | ( (~ n294)  &  n815 ) ;
 assign n494 = ( n495  &  n496 ) ;
 assign n497 = ( (~ n265)  &  n408 ) ;
 assign n498 = ( n506  &  n23 ) | ( n506  &  n625 ) ;
 assign n499 = ( PV149_3_ ) | ( n247 ) | ( n267 ) ;
 assign n501 = ( PV174_0_  &  (~ n740) ) | ( n230  &  (~ n740) ) ;
 assign n503 = ( PV165_7_ ) | ( PV165_3_ ) | ( PV165_6_ ) ;
 assign n502 = ( PV165_5_  &  (~ n32) ) | ( PV165_4_  &  (~ n32) ) | ( (~ n32)  &  n503 ) ;
 assign n506 = ( PV174_0_ ) | ( n247 ) | ( n248 ) ;
 assign n507 = ( PV302_0_  &  (~ n23) ) | ( (~ n23)  &  n267 ) | ( PV302_0_  &  n392 ) | ( n267  &  n392 ) ;
 assign n505 = ( n506  &  n223  &  n507 ) ;
 assign n510 = ( n229 ) | ( n826 ) ;
 assign n508 = ( n229  &  n510 ) | ( n510  &  (~ n825) ) ;
 assign n511 = ( (~ PV14_0_) ) | ( (~ n510) ) | ( (~ n1011) ) ;
 assign n522 = ( n247 ) | ( n717 ) ;
 assign n524 = ( (~ n122) ) | ( (~ n1024) ) ;
 assign n523 = ( (~ n199)  &  n524 ) ;
 assign n531 = ( (~ PV59_0_) ) | ( n777 ) ;
 assign n532 = ( PV274_0_  &  PV172_0_ ) | ( PV271_0_  &  PV172_0_ ) | ( PV274_0_  &  (~ n243) ) | ( PV271_0_  &  (~ n243) ) ;
 assign n529 = ( PV248_0_ ) | ( n162 ) | ( (~ n723) ) ;
 assign n534 = ( (~ PV174_0_)  &  (~ n85) ) | ( (~ n85)  &  (~ n239)  &  n732 ) ;
 assign n535 = ( (~ PV91_1_)  &  (~ PV91_0_) ) | ( (~ PV91_0_)  &  (~ PV62_0_) ) | ( (~ PV91_1_)  &  (~ PV59_0_) ) | ( (~ PV62_0_)  &  (~ PV59_0_) ) ;
 assign n538 = ( PV294_0_ ) | ( (~ n261) ) | ( n959 ) ;
 assign n540 = ( PV289_0_ ) | ( (~ PV14_0_) ) | ( (~ n268) ) | ( n505 ) ;
 assign n544 = ( n543 ) | ( n826 ) ;
 assign n543 = ( n710  &  n563 ) ;
 assign n542 = ( n544  &  n543 ) | ( n544  &  (~ n825) ) ;
 assign n545 = ( (~ PV14_0_) ) | ( (~ n544) ) | ( (~ n1014) ) ;
 assign n554 = ( (~ PV242_0_) ) | ( (~ PV14_0_) ) | ( n725 ) ;
 assign n553 = ( (~ PV194_0_) ) | ( n694 ) ;
 assign n556 = ( n250 ) | ( n196 ) ;
 assign n555 = ( PV56_0_  &  (~ n600) ) ;
 assign n558 = ( (~ PV108_0_) ) | ( n559 ) ;
 assign n559 = ( PV56_0_  &  n839 ) ;
 assign n563 = ( PV149_2_ ) | ( PV149_1_ ) | ( PV149_0_ ) ;
 assign n568 = ( (~ PV124_5_)  &  (~ PV100_5_) ) | ( (~ PV100_5_)  &  n588 ) | ( (~ PV124_5_)  &  n722 ) | ( n588  &  n722 ) ;
 assign n567 = ( n717 ) | ( n255 ) ;
 assign n570 = ( (~ PV213_4_)  &  (~ PV100_4_) ) | ( (~ PV100_4_)  &  n567 ) | ( (~ PV213_4_)  &  n722 ) | ( n567  &  n722 ) ;
 assign n571 = ( (~ PV124_4_)  &  (~ PV108_4_) ) | ( (~ PV108_4_)  &  n588 ) | ( (~ PV124_4_)  &  (~ n839) ) | ( n588  &  (~ n839) ) ;
 assign n569 = ( n570  &  n571 ) ;
 assign n575 = ( (~ PV213_3_)  &  (~ PV100_3_) ) | ( (~ PV100_3_)  &  n567 ) | ( (~ PV213_3_)  &  n722 ) | ( n567  &  n722 ) ;
 assign n576 = ( (~ PV124_3_)  &  (~ PV108_3_) ) | ( (~ PV108_3_)  &  n588 ) | ( (~ PV124_3_)  &  (~ n839) ) | ( n588  &  (~ n839) ) ;
 assign n574 = ( n575  &  n576 ) ;
 assign n578 = ( (~ PV213_2_)  &  (~ PV100_2_) ) | ( (~ PV100_2_)  &  n567 ) | ( (~ PV213_2_)  &  n722 ) | ( n567  &  n722 ) ;
 assign n579 = ( (~ PV124_2_)  &  (~ PV108_2_) ) | ( (~ PV108_2_)  &  n588 ) | ( (~ PV124_2_)  &  (~ n839) ) | ( n588  &  (~ n839) ) ;
 assign n577 = ( n578  &  n579 ) ;
 assign n581 = ( (~ PV213_1_)  &  (~ PV100_1_) ) | ( (~ PV100_1_)  &  n567 ) | ( (~ PV213_1_)  &  n722 ) | ( n567  &  n722 ) ;
 assign n582 = ( (~ PV124_1_)  &  (~ PV108_1_) ) | ( (~ PV108_1_)  &  n588 ) | ( (~ PV124_1_)  &  (~ n839) ) | ( n588  &  (~ n839) ) ;
 assign n580 = ( n581  &  n582 ) ;
 assign n584 = ( (~ PV213_0_)  &  (~ PV100_0_) ) | ( (~ PV100_0_)  &  n567 ) | ( (~ PV213_0_)  &  n722 ) | ( n567  &  n722 ) ;
 assign n585 = ( (~ PV124_0_)  &  (~ PV108_0_) ) | ( (~ PV108_0_)  &  n588 ) | ( (~ PV124_0_)  &  (~ n839) ) | ( n588  &  (~ n839) ) ;
 assign n583 = ( n584  &  n585 ) ;
 assign n586 = ( n717 ) | ( n720 ) ;
 assign n588 = ( n720 ) | ( n256 ) ;
 assign n600 = ( PV149_7_ ) | ( (~ PV149_6_) ) | ( n739 ) ;
 assign n604 = ( PV134_1_ ) | ( n849 ) ;
 assign n603 = ( (~ n787) ) | ( n847 ) ;
 assign n605 = ( PV202_0_  &  PV274_0_ ) ;
 assign n606 = ( PV174_0_  &  (~ PV52_0_) ) | ( (~ PV52_0_)  &  (~ n835) ) ;
 assign n611 = ( PV257_5_  &  n853 ) ;
 assign n610 = ( n611  &  PV257_4_ ) ;
 assign n616 = ( PV802_0_ ) | ( n289 ) | ( (~ n553) ) ;
 assign n614 = ( (~ n553)  &  n616 ) | ( n616  &  (~ n725) ) ;
 assign n617 = ( (~ PV1378)  &  (~ PV782) ) | ( (~ PV1378)  &  n71 ) | ( (~ PV1378)  &  n614 ) ;
 assign n621 = ( (~ PV134_1_) ) | ( (~ PV134_0_) ) | ( (~ n71) ) | ( (~ n553) ) | ( n787 ) ;
 assign n623 = ( n830  &  PV268_3_ ) ;
 assign n622 = ( PV268_2_  &  n623 ) ;
 assign n625 = ( PV149_4_ ) | ( n744 ) | ( n775 ) | ( n776 ) ;
 assign n624 = ( n73  &  (~ n136)  &  n287  &  n625 ) ;
 assign n626 = ( PV239_4_  &  n12 ) | ( n695  &  n12 ) | ( PV239_4_  &  n390 ) | ( n695  &  n390 ) ;
 assign n627 = ( n696  &  n10 ) | ( n695  &  n10 ) | ( n696  &  n390 ) | ( n695  &  n390 ) ;
 assign n628 = ( (~ PV118_7_)  &  (~ PV46_0_) ) | ( (~ PV46_0_)  &  n586 ) | ( (~ PV118_7_)  &  n699 ) | ( n586  &  n699 ) ;
 assign n629 = ( (~ PV118_6_)  &  (~ PV48_0_) ) | ( (~ PV48_0_)  &  n586 ) | ( (~ PV118_6_)  &  n699 ) | ( n586  &  n699 ) ;
 assign n631 = ( (~ n764)  &  n639 ) | ( n764  &  (~ n639) ) ;
 assign n630 = ( (~ n319)  &  n631 ) | ( n319  &  (~ n631) ) ;
 assign n632 = ( n307  &  n320 ) | ( (~ n307)  &  (~ n320) ) ;
 assign n633 = ( (~ n305)  &  n321 ) | ( n305  &  (~ n321) ) ;
 assign n634 = ( n315  &  n632 ) | ( (~ n315)  &  (~ n632) ) ;
 assign n637 = ( (~ n315)  &  (~ n630) ) | ( (~ n315)  &  (~ n632) ) | ( n630  &  (~ n632) ) ;
 assign n636 = ( n321  &  n634 ) | ( (~ n630)  &  n634 ) | ( n321  &  n637 ) | ( (~ n630)  &  n637 ) ;
 assign n638 = ( (~ n38)  &  n632 ) | ( n38  &  (~ n632) ) ;
 assign n639 = ( (~ PV288_7_)  &  (~ PV288_6_) ) ;
 assign n642 = ( (~ PV802_0_)  &  n740 ) ;
 assign n641 = ( (~ n35) ) | ( n642 ) ;
 assign n643 = ( (~ n37)  &  n634 ) | ( n37  &  (~ n634) ) ;
 assign n644 = ( (~ n37)  &  n315 ) | ( n37  &  (~ n315) ) ;
 assign n646 = ( (~ n632)  &  n861 ) ;
 assign n647 = ( n764  &  n319  &  n639 ) ;
 assign n645 = ( n320  &  n646 ) | ( n320  &  n647 ) ;
 assign n648 = ( n35  &  n645 ) | ( (~ n35)  &  (~ n645) ) ;
 assign n649 = ( n320  &  n638 ) | ( (~ n320)  &  (~ n638) ) ;
 assign n653 = ( (~ PV288_3_) ) | ( PV288_2_ ) ;
 assign n651 = ( (~ n632)  &  (~ n765) ) | ( n653  &  (~ n765) ) ;
 assign n654 = ( n314  &  n93 ) ;
 assign n655 = ( n630  &  n654 ) | ( (~ n630)  &  (~ n654) ) ;
 assign n657 = ( (~ n324)  &  n647 ) | ( n324  &  (~ n647) ) ;
 assign n658 = ( n350  &  n346 ) ;
 assign n656 = ( n657  &  n658 ) | ( n658  &  (~ n765) ) | ( n657  &  (~ n972) ) | ( (~ n765)  &  (~ n972) ) ;
 assign n660 = ( n90  &  n653 ) | ( (~ n90)  &  (~ n653) ) ;
 assign n661 = ( (~ n112)  &  n310 ) ;
 assign n662 = ( n655  &  n661 ) | ( (~ n655)  &  (~ n661) ) ;
 assign n665 = ( (~ PV288_1_) ) | ( PV288_0_ ) ;
 assign n664 = ( n312  &  (~ n351) ) | ( n312  &  n665 ) ;
 assign n666 = ( (~ n651)  &  n315 ) | ( n651  &  (~ n315) ) ;
 assign n667 = ( (~ n169)  &  n330 ) ;
 assign n670 = ( n333  &  n332  &  n326 ) ;
 assign n669 = ( n169  &  (~ n667) ) | ( n312  &  (~ n667) ) | ( n169  &  n670 ) | ( n312  &  n670 ) ;
 assign n672 = ( n105  &  n665 ) | ( (~ n105)  &  (~ n665) ) ;
 assign n673 = ( (~ PV84_5_)  &  PV84_4_ ) | ( PV84_5_  &  (~ PV84_4_) ) ;
 assign n674 = ( (~ PV84_3_)  &  n1027 ) | ( PV84_3_  &  (~ n1027) ) ;
 assign n675 = ( (~ PV78_1_)  &  PV78_0_ ) | ( PV78_1_  &  (~ PV78_0_) ) ;
 assign n676 = ( (~ PV78_3_)  &  n1029 ) | ( PV78_3_  &  (~ n1029) ) ;
 assign n678 = ( PV199_3_  &  PV199_4_ ) ;
 assign n682 = ( n429  &  PV199_0_  &  PV199_1_ ) ;
 assign n685 = ( n682  &  PV194_4_ ) ;
 assign n684 = ( PV194_3_  &  n685 ) | ( (~ PV194_3_)  &  (~ n685) ) ;
 assign n688 = ( n685  &  PV194_3_ ) ;
 assign n687 = ( PV194_2_  &  n688 ) | ( (~ PV194_2_)  &  (~ n688) ) ;
 assign n691 = ( n688  &  PV194_2_ ) ;
 assign n690 = ( PV194_1_  &  n691 ) | ( (~ PV194_1_)  &  (~ n691) ) ;
 assign n694 = ( (~ PV194_1_) ) | ( (~ n691) ) ;
 assign n693 = ( (~ n694)  &  PV194_0_ ) | ( n694  &  (~ PV194_0_) ) ;
 assign n695 = ( PV802_0_ ) | ( (~ n136) ) ;
 assign n696 = ( PV239_4_  &  PV239_3_ ) | ( (~ PV239_4_)  &  (~ PV239_3_) ) ;
 assign n699 = ( n261  &  n225 ) ;
 assign n703 = ( (~ n948)  &  n949 ) | ( n948  &  (~ n949) ) ;
 assign n704 = ( (~ n950)  &  n1033 ) | ( n950  &  (~ n1033) ) ;
 assign n707 = ( (~ PV149_2_) ) | ( (~ PV149_1_) ) | ( PV149_0_ ) ;
 assign n710 = ( PV149_2_ ) | ( (~ PV149_1_) ) | ( PV149_0_ ) ;
 assign n711 = ( (~ PV149_7_) ) | ( PV149_3_ ) | ( n710 ) ;
 assign n714 = ( PV149_7_ ) | ( PV149_3_ ) | ( n710 ) ;
 assign n715 = ( (~ PV149_6_) ) | ( n714 ) ;
 assign n717 = ( PV149_6_ ) | ( n711 ) ;
 assign n718 = ( (~ PV149_5_) ) | ( PV149_4_ ) ;
 assign n720 = ( PV149_5_ ) | ( (~ PV149_4_) ) ;
 assign n721 = ( n715 ) | ( n720 ) ;
 assign n722 = ( n715 ) | ( n255 ) ;
 assign n723 = ( (~ PV172_0_) ) | ( (~ PV56_0_) ) ;
 assign n725 = ( (~ n73) ) | ( (~ n283) ) ;
 assign n731 = ( PV172_0_  &  PV215_0_  &  PV67_0_ ) ;
 assign n730 = ( n731 ) | ( n269 ) | ( PV214_0_ ) | ( n191 ) ;
 assign n735 = ( (~ PV261_0_) ) | ( PV802_0_ ) | ( n71 ) | ( (~ n263) ) ;
 assign n736 = ( PV275_0_ ) | ( (~ PV272_0_) ) | ( PV802_0_ ) | ( (~ n71) ) | ( n270 ) ;
 assign n732 = ( (~ n272)  &  (~ n730)  &  n735  &  n736 ) ;
 assign n739 = ( (~ PV149_3_) ) | ( n255 ) | ( n710 ) ;
 assign n740 = ( (~ PV149_7_)  &  (~ PV149_6_)  &  (~ n739) ) ;
 assign n744 = ( PV149_3_ ) | ( n392 ) ;
 assign n750 = ( n253 ) | ( n122 ) ;
 assign n748 = ( (~ n122)  &  (~ n280)  &  n750  &  (~ n794) ) ;
 assign n752 = ( n295 ) | ( (~ n748) ) ;
 assign n754 = ( (~ n163) ) | ( n752 ) ;
 assign n762 = ( (~ PV288_6_) ) | ( (~ n36) ) | ( n641 ) ;
 assign n763 = ( (~ PV288_7_) ) | ( n37 ) | ( n762 ) ;
 assign n764 = ( (~ PV288_5_) ) | ( (~ PV288_4_) ) ;
 assign n765 = ( (~ PV288_3_)  &  PV288_2_ ) ;
 assign n766 = ( n295 ) | ( n439 ) ;
 assign n775 = ( PV149_5_  &  n20 ) ;
 assign n776 = ( (~ PV149_5_)  &  PV88_3_ ) | ( (~ PV149_5_)  &  PV88_2_ ) ;
 assign n777 = ( (~ n23) ) | ( n625 ) ;
 assign n783 = ( n32 ) | ( PV214_0_ ) | ( PV43_0_ ) ;
 assign n787 = ( PV274_0_ ) | ( (~ PV271_0_) ) | ( (~ n25) ) ;
 assign n788 = ( n274 ) | ( (~ n621) ) ;
 assign n791 = ( (~ PV802_0_) ) | ( n283 ) ;
 assign n790 = ( n396  &  n791  &  n788 ) ;
 assign n792 = ( (~ n143) ) | ( n750 ) ;
 assign n794 = ( (~ n283)  &  n281 ) ;
 assign n795 = ( n122 ) | ( (~ n280) ) | ( (~ n794) ) ;
 assign n797 = ( n295 ) | ( n792 ) ;
 assign n801 = ( n788 ) | ( n791 ) ;
 assign n815 = ( n295 ) | ( n418 ) ;
 assign n824 = ( (~ PV14_0_) ) | ( n278 ) ;
 assign n825 = ( n230  &  n540  &  n268 ) ;
 assign n826 = ( (~ PV290_0_) ) | ( (~ n239) ) ;
 assign n830 = ( PV268_5_  &  PV268_4_ ) ;
 assign n831 = ( n623  &  PV268_2_  &  PV268_1_ ) ;
 assign n832 = ( (~ PV288_4_) ) | ( (~ n638) ) | ( n641 ) | ( n864 ) | ( n865 ) ;
 assign n833 = ( n649 ) | ( n858 ) | ( n862 ) | ( n642 ) | ( n361 ) | ( n648 ) ;
 assign n835 = ( PV56_0_  &  (~ n84) ) ;
 assign n839 = ( PV149_7_  &  (~ PV149_6_)  &  (~ n739) ) ;
 assign n847 = ( PV802_0_  &  n725 ) ;
 assign n849 = ( n847 ) | ( n787 ) ;
 assign n853 = ( PV257_7_  &  PV257_6_ ) ;
 assign n854 = ( PV257_4_  &  PV257_3_  &  n611 ) ;
 assign n857 = ( (~ n632)  &  n634 ) | ( n632  &  (~ n634) ) ;
 assign n859 = ( (~ n320)  &  n971 ) | ( n636  &  (~ n646)  &  n971 ) ;
 assign n858 = ( (~ n36)  &  n859 ) | ( n36  &  (~ n859) ) ;
 assign n861 = ( n315  &  (~ n321) ) | ( n315  &  n857 ) | ( n321  &  n857 ) ;
 assign n860 = ( n632  &  n861 ) | ( (~ n632)  &  (~ n861) ) ;
 assign n863 = ( n315  &  (~ n320) ) | ( n315  &  n860 ) | ( n320  &  n860 ) ;
 assign n862 = ( (~ n37)  &  n863 ) | ( n37  &  (~ n863) ) ;
 assign n864 = ( (~ n36)  &  n636 ) | ( n36  &  (~ n636) ) ;
 assign n865 = ( (~ n37)  &  n861 ) | ( n37  &  (~ n861) ) ;
 assign n866 = ( (~ n36)  &  n637 ) | ( n36  &  (~ n637) ) ;
 assign n867 = ( n36  &  n630 ) | ( (~ n36)  &  (~ n630) ) ;
 assign n869 = ( (~ n351)  &  n355  &  n354 ) ;
 assign n868 = ( (~ n869)  &  n656 ) | ( n869  &  (~ n656) ) ;
 assign n871 = ( (~ n653)  &  n657 ) | ( n653  &  n868 ) | ( n657  &  n868 ) ;
 assign n870 = ( (~ n35)  &  n871 ) | ( n35  &  (~ n871) ) ;
 assign n873 = ( n353  &  n653 ) | ( n353  &  (~ n655) ) | ( (~ n653)  &  (~ n655) ) ;
 assign n872 = ( (~ n36)  &  n873 ) | ( n36  &  (~ n873) ) ;
 assign n874 = ( n351  &  n354 ) | ( (~ n351)  &  (~ n354) ) ;
 assign n876 = ( (~ n653)  &  (~ n666) ) | ( n653  &  n874 ) | ( (~ n666)  &  n874 ) ;
 assign n875 = ( (~ n37)  &  n876 ) | ( n37  &  (~ n876) ) ;
 assign n878 = ( (~ n333)  &  n332 ) | ( n333  &  (~ n332) ) ;
 assign n879 = ( (~ n669)  &  n1016 ) | ( n669  &  (~ n1016) ) ;
 assign n882 = ( n169  &  (~ n665) ) | ( n169  &  n879 ) | ( n665  &  n879 ) ;
 assign n881 = ( (~ n35)  &  n882 ) | ( n35  &  (~ n882) ) ;
 assign n884 = ( n335  &  (~ n662) ) | ( n335  &  n665 ) | ( (~ n662)  &  (~ n665) ) ;
 assign n883 = ( (~ n36)  &  n884 ) | ( n36  &  (~ n884) ) ;
 assign n885 = ( n333  &  n336 ) | ( (~ n333)  &  (~ n336) ) ;
 assign n887 = ( n327  &  (~ n665) ) | ( n327  &  n885 ) | ( n665  &  n885 ) ;
 assign n886 = ( (~ n37)  &  n887 ) | ( n37  &  (~ n887) ) ;
 assign n889 = ( (~ PV280_0_)  &  PV279_0_ ) | ( PV280_0_  &  (~ PV279_0_) ) ;
 assign n890 = ( (~ n951)  &  n952 ) | ( n951  &  (~ n952) ) ;
 assign n891 = ( (~ n953)  &  n954 ) | ( n953  &  (~ n954) ) ;
 assign n892 = ( (~ PV39_0_)  &  PV38_0_ ) | ( PV39_0_  &  (~ PV38_0_) ) ;
 assign n893 = ( (~ PV42_0_)  &  PV44_0_ ) | ( PV42_0_  &  (~ PV44_0_) ) ;
 assign n894 = ( (~ PV244_0_)  &  n981 ) | ( n460  &  n981 ) ;
 assign n895 = ( (~ PV244_0_)  &  n982 ) | ( (~ PV245_0_)  &  PV243_0_  &  n982 ) ;
 assign n896 = ( PV279_0_  &  (~ PV149_5_) ) | ( PV279_0_  &  n387 ) | ( (~ PV149_5_)  &  (~ n387) ) ;
 assign n897 = ( (~ PV149_4_)  &  (~ n387) ) | ( (~ PV149_4_)  &  n889 ) | ( n387  &  n889 ) ;
 assign n898 = ( n502  &  (~ n508) ) | ( n502  &  n985 ) | ( n508  &  n985 ) ;
 assign n899 = ( (~ PV1536_0_)  &  n3 ) | ( PV1536_0_  &  (~ n732) ) | ( n3  &  (~ n732) ) ;
 assign n900 = ( PV1536_0_  &  (~ n990) ) | ( n218  &  n219  &  (~ n990) ) ;
 assign n901 = ( (~ PV1536_0_)  &  (~ n992) ) | ( n732  &  n835  &  (~ n992) ) ;
 assign n902 = ( n502  &  (~ n542) ) | ( n502  &  n997 ) | ( n542  &  n997 ) ;
 assign n903 = ( PV134_1_  &  PV88_3_ ) | ( PV134_1_  &  n25 ) | ( PV88_3_  &  (~ n25) ) ;
 assign n904 = ( PV134_0_  &  PV88_2_ ) | ( PV134_0_  &  n25 ) | ( PV88_2_  &  (~ n25) ) ;
 assign n905 = ( PV78_3_  &  (~ n25) ) | ( PV78_3_  &  (~ n45) ) | ( n25  &  (~ n45) ) ;
 assign n906 = ( PV78_2_  &  (~ n25) ) | ( PV78_2_  &  (~ n44) ) | ( n25  &  (~ n44) ) ;
 assign n907 = ( (~ PV37_0_)  &  (~ PV321_2_) ) | ( PV37_0_  &  (~ n12) ) | ( (~ PV321_2_)  &  (~ n12) ) ;
 assign n908 = ( PV37_0_  &  (~ n10) ) | ( (~ PV37_0_)  &  (~ n45) ) | ( (~ n10)  &  (~ n45) ) ;
 assign n909 = ( PV37_0_  &  (~ n11) ) | ( (~ PV37_0_)  &  (~ n44) ) | ( (~ n11)  &  (~ n44) ) ;
 assign n910 = ( (~ PV37_0_)  &  (~ n43) ) | ( PV37_0_  &  (~ n56) ) | ( (~ n43)  &  (~ n56) ) ;
 assign n911 = ( (~ PV37_0_)  &  (~ n42) ) | ( PV37_0_  &  (~ n57) ) | ( (~ n42)  &  (~ n57) ) ;
 assign n912 = ( (~ PV37_0_)  &  (~ n41) ) | ( PV37_0_  &  (~ n58) ) | ( (~ n41)  &  (~ n58) ) ;
 assign n913 = ( (~ PV37_0_)  &  (~ n40) ) | ( PV37_0_  &  (~ n59) ) | ( (~ n40)  &  (~ n59) ) ;
 assign n914 = ( (~ PV37_0_)  &  (~ n39) ) | ( PV37_0_  &  (~ n60) ) | ( (~ n39)  &  (~ n60) ) ;
 assign n915 = ( PV37_0_  &  (~ n61) ) | ( (~ PV37_0_)  &  (~ n494) ) | ( (~ n61)  &  (~ n494) ) ;
 assign n916 = ( (~ PV37_0_)  &  (~ PV321_2_) ) | ( PV37_0_  &  (~ n37) ) | ( (~ PV321_2_)  &  (~ n37) ) ;
 assign n918 = ( PV108_4_ ) | ( (~ PV101_0_) ) | ( n195 ) ;
 assign n917 = ( (~ PV56_0_)  &  PV14_0_  &  n918 ) | ( PV14_0_  &  n586  &  n918 ) ;
 assign n919 = ( (~ PV110_0_)  &  (~ n1001) ) | ( (~ n917)  &  (~ n1001) ) ;
 assign n920 = ( (~ PV134_0_)  &  n1003 ) | ( n604  &  n603  &  n1003 ) ;
 assign n921 = ( PV271_0_  &  PV269_0_ ) | ( (~ PV271_0_)  &  n605 ) | ( PV269_0_  &  n605 ) ;
 assign n922 = ( (~ PV165_5_) ) | ( (~ PV165_4_) ) | ( (~ PV165_3_) ) ;
 assign n923 = ( (~ PV290_0_)  &  PV14_0_ ) | ( PV14_0_  &  n239 ) ;
 assign n924 = ( PV149_5_  &  (~ PV149_4_) ) | ( (~ PV149_4_)  &  (~ PV88_3_)  &  (~ PV88_2_) ) ;
 assign n925 = ( n833  &  n832  &  n5 ) ;
 assign n926 = ( n93  &  (~ n112) ) | ( n93  &  n342 ) | ( (~ n112)  &  n360 ) | ( n342  &  n360 ) ;
 assign n928 = ( (~ n10)  &  n364 ) | ( (~ n10)  &  n366 ) | ( (~ n10)  &  (~ n926) ) ;
 assign n930 = ( (~ PV802_0_)  &  n386 ) | ( n287  &  n386 ) ;
 assign n931 = ( (~ PV88_3_)  &  PV88_2_ ) | ( PV88_3_  &  (~ PV88_2_) ) ;
 assign n932 = ( (~ PV88_0_)  &  PV84_2_ ) | ( PV88_0_  &  (~ PV84_2_) ) ;
 assign n933 = ( (~ PV94_1_)  &  n932 ) | ( PV94_1_  &  (~ n932) ) ;
 assign n934 = ( (~ PV84_1_)  &  PV84_0_ ) | ( PV84_1_  &  (~ PV84_0_) ) ;
 assign n935 = ( (~ PV78_4_)  &  PV78_2_ ) | ( PV78_4_  &  (~ PV78_2_) ) ;
 assign n936 = ( (~ PV94_0_)  &  n935 ) | ( PV94_0_  &  (~ n935) ) ;
 assign n937 = ( (~ PV1719) ) | ( (~ PV302_0_)  &  (~ n9) ) ;
 assign n939 = ( (~ PV62_0_) ) | ( n261 ) ;
 assign n940 = ( (~ PV149_4_)  &  (~ PV32_5_) ) | ( (~ PV149_4_)  &  n792 ) | ( (~ PV32_5_)  &  n795 ) | ( n792  &  n795 ) ;
 assign n943 = ( (~ PV278_0_)  &  PV177_0_ ) | ( PV177_0_  &  (~ n265) ) ;
 assign n944 = ( (~ n86)  &  n216  &  n344 ) ;
 assign n946 = ( PV280_0_  &  (~ n9) ) | ( (~ n9)  &  (~ n136) ) ;
 assign n948 = ( (~ n207)  &  n208 ) | ( n207  &  (~ n208) ) ;
 assign n949 = ( (~ n209)  &  n210 ) | ( n209  &  (~ n210) ) ;
 assign n950 = ( (~ n628)  &  n629 ) | ( n628  &  (~ n629) ) ;
 assign n951 = ( (~ PV1953_1_)  &  n206 ) | ( PV1953_1_  &  (~ n206) ) ;
 assign n952 = ( (~ n569)  &  n574 ) | ( n569  &  (~ n574) ) ;
 assign n953 = ( (~ n577)  &  n580 ) | ( n577  &  (~ n580) ) ;
 assign n954 = ( (~ n213)  &  n583 ) | ( n213  &  (~ n583) ) ;
 assign n955 = ( (~ PV59_0_)  &  (~ n1026) ) | ( n497  &  (~ n1026) ) ;
 assign n957 = ( (~ PV56_0_)  &  (~ PV802_0_) ) | ( (~ PV56_0_)  &  n82 ) | ( (~ PV802_0_)  &  n254 ) | ( n82  &  n254 ) ;
 assign n959 = ( (~ n152)  &  (~ n224) ) ;
 assign n958 = ( PV59_0_  &  (~ n410) ) | ( PV59_0_  &  n959 ) ;
 assign n961 = ( PV214_0_ ) | ( (~ PV62_0_) ) | ( n239 ) | ( n261 ) ;
 assign n962 = ( (~ PV66_0_) ) | ( n151 ) ;
 assign n963 = ( (~ PV248_0_)  &  n735 ) | ( PV802_0_  &  n735 ) ;
 assign n964 = ( (~ n18) ) | ( n23 ) ;
 assign n965 = ( n23 ) | ( (~ n506) ) ;
 assign n966 = ( (~ PV59_0_)  &  (~ n223) ) | ( (~ PV59_0_)  &  n965 ) | ( (~ n223)  &  (~ n965) ) ;
 assign n971 = ( n320 ) | ( (~ n630) ) ;
 assign n972 = ( (~ n348)  &  n657 ) | ( n348  &  (~ n657) ) ;
 assign n974 = ( (~ n35)  &  (~ n642) ) ;
 assign n973 = ( (~ n641)  &  (~ n972) ) | ( (~ n641)  &  n974 ) | ( n972  &  n974 ) ;
 assign n976 = ( (~ n351)  &  n350 ) | ( n351  &  (~ n350) ) ;
 assign n978 = ( (~ n641)  &  (~ n667) ) | ( (~ n641)  &  n974 ) | ( n667  &  n974 ) ;
 assign n980 = ( (~ PV66_0_)  &  (~ n253) ) | ( (~ PV66_0_)  &  n395 ) | ( n253  &  n395 ) ;
 assign n981 = ( PV244_0_ ) | ( (~ PV243_0_) ) | ( (~ n64) ) ;
 assign n982 = ( PV244_0_ ) | ( PV245_0_ ) ;
 assign n985 = ( (~ PV213_0_) ) | ( (~ PV14_0_) ) | ( (~ n1011) ) ;
 assign n986 = ( PV258_0_  &  (~ n199) ) | ( (~ PV258_0_)  &  n524 ) | ( (~ n199)  &  n524 ) ;
 assign n988 = ( (~ PV259_0_) ) | ( (~ PV258_0_) ) | ( (~ n199) ) ;
 assign n987 = ( n988  &  PV259_0_ ) | ( n988  &  n524 ) | ( n988  &  PV258_0_ ) ;
 assign n990 = ( PV1536_0_  &  (~ n31) ) | ( PV1536_0_  &  (~ n732) ) ;
 assign n992 = ( (~ PV1536_0_)  &  (~ n7) ) | ( (~ PV1536_0_)  &  n101 ) | ( (~ PV1536_0_)  &  (~ n944) ) ;
 assign n997 = ( (~ PV100_0_) ) | ( (~ PV14_0_) ) | ( (~ n1014) ) ;
 assign n1001 = ( (~ PV110_0_)  &  PV102_0_  &  (~ n563) ) | ( (~ PV110_0_)  &  (~ n194)  &  (~ n563) ) ;
 assign n1003 = ( (~ PV134_1_) ) | ( PV134_0_ ) | ( n849 ) ;
 assign n1005 = ( PV248_0_ ) | ( (~ PV1719) ) | ( n376 ) ;
 assign n1006 = ( PV15_0_ ) | ( (~ PV423_0_) ) | ( n122 ) | ( n152 ) | ( n158 ) | ( n168 ) | ( n242 ) | ( n783 ) ;
 assign n1008 = ( n892 ) | ( n893 ) ;
 assign n1010 = ( n253 ) | ( n606 ) | ( (~ n835) ) ;
 assign n1011 = ( (~ PV56_0_) ) | ( n567 ) ;
 assign n1014 = ( (~ PV56_0_) ) | ( n722 ) ;
 assign n1016 = ( (~ n333)  &  n337  &  n336 ) ;
 assign n1020 = ( n6  &  n8  &  (~ n122)  &  n215  &  n222 ) ;
 assign n1022 = ( n393  &  (~ n397)  &  n962  &  n980 ) ;
 assign n1024 = ( PV56_0_ ) | ( PV62_0_ ) | ( PV50_0_ ) ;
 assign n1025 = ( PV215_0_  &  PV14_0_  &  n157  &  (~ n730) ) ;
 assign n1026 = ( n254  &  n119  &  n1010  &  PV56_0_ ) ;
 assign n1028 = ( PV88_1_  &  n931 ) | ( (~ PV88_1_)  &  (~ n931) ) ;
 assign n1027 = ( (~ n933)  &  n1028 ) | ( n933  &  (~ n1028) ) ;
 assign n1030 = ( PV78_5_  &  n934 ) | ( (~ PV78_5_)  &  (~ n934) ) ;
 assign n1029 = ( (~ n936)  &  n1030 ) | ( n936  &  (~ n1030) ) ;
 assign n1033 = ( n211  &  n212 ) | ( (~ n211)  &  (~ n212) ) ;
 assign PV1757_0_ = ( PV15_0_ ) ;


endmodule

