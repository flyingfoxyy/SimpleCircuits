module apex4_mapped (
	i_7_, i_8_, i_5_, i_6_, i_3_, i_4_, i_1_, i_2_, 
	i_0_, o_1_, o_2_, o_0_, o_12_, o_11_, o_14_, o_13_, o_16_, o_15_, 
	o_18_, o_17_, o_10_, o_9_, o_7_, o_8_, o_5_, o_6_, o_3_, o_4_);

input i_7_, i_8_, i_5_, i_6_, i_3_, i_4_, i_1_, i_2_, i_0_;

output o_1_, o_2_, o_0_, o_12_, o_11_, o_14_, o_13_, o_16_, o_15_, o_18_, o_17_, o_10_, o_9_, o_7_, o_8_, o_5_, o_6_, o_3_, o_4_;

wire n_n110, wire4865, wire4866, wire4867, wire4989, wire4990, wire4991, wire5046, wire5047, wire5049, wire5066, wire5067, wire5108, wire5111, wire5125, wire5126, wire5166, wire5169, wire5218, wire5219, wire5221, wire5228, wire5229, wire5233, wire5249, wire5250, wire5260, wire5261, wire5265, wire5268, wire5269, wire5270, n_n655, wire5369, wire5370, wire5373, n_n586, wire5487, wire5488, wire5489, wire5540, wire5590, wire5658, wire5684, wire5733, wire5780, wire5821, wire5822, wire5875, wire5876, wire5934, wire5935, wire5940, wire5941, n_n243, wire6024, wire6025, wire6028, n_n80, n_n75, n_n81, n_n58, n_n101, n_n93, n_n78, n_n91, n_n99, n_n103, n_n1281, n_n100, n_n84, n_n1185, n_n1164, n_n1021, wire4837, wire4838, n_n97, n_n1174, wire172, wire192, n_n96, wire235, n_n92, wire252, wire329, n_n74, n_n1077, n_n82, n_n95, n_n90, n_n1172, n_n1078, n_n54, wire245, n_n1081, n_n1279, n_n1181, wire243, wire295, wire4923, n_n137, wire231, wire1512, wire1513, wire4936, n_n135, n_n102, n_n1153, wire308, wire304, wire4942, n_n136, n_n1297, n_n1324, n_n1092, n_n1108, n_n1105, wire4949, wire4950, n_n139, wire127, n_n83, wire35, wire1477, wire1479, wire232, n_n63, n_n77, wire251, wire321, n_n1254, n_n1259, n_n1204, wire4994, n_n1369, wire1516, wire1518, wire1519, wire1408, wire1409, wire1410, wire301, n_n85, wire314, wire349, n_n1022, n_n1134, n_n94, n_n1039, wire241, n_n87, n_n1091, wire322, n_n1093, n_n1103, n_n1120, n_n1052, n_n1331, n_n38, n_n40, wire177, n_n1109, wire1345, wire1348, wire257, n_n1193, n_n1330, n_n1267, wire342, wire346, wire323, wire352, wire357, n_n1176, n_n1074, n_n1032, n_n1294, n_n1312, wire326, wire5222, wire310, n_n1169, n_n942, n_n1057, n_n1125, n_n1128, wire248, n_n1046, n_n1042, n_n1047, wire302, n_n1286, n_n79, n_n937, wire351, wire189, n_n1283, n_n1087, n_n663, wire5312, wire5313, wire5314, n_n71, n_n968, n_n958, n_n66, n_n974, n_n973, n_n989, n_n64, n_n938, n_n944, n_n70, n_n982, n_n967, n_n956, n_n1121, n_n53, wire4880, wire4881, wire70, n_n962, n_n961, n_n964, wire168, wire236, n_n941, n_n949, n_n943, wire291, n_n954, n_n952, n_n951, wire297, n_n960, n_n959, n_n957, wire298, wire319, n_n1082, n_n324, n_n397, wire5403, n_n1045, n_n1043, n_n1122, n_n1036, n_n1118, n_n1030, wire5442, n_n1083, n_n1101, n_n1156, wire5448, wire5449, n_n593, n_n1060, wire1104, wire5452, wire5453, n_n597, wire355, n_n1100, n_n969, n_n939, wire131, n_n971, n_n1035, n_n1037, wire334, wire345, wire903, n_n421, n_n1058, n_n947, wire831, wire5541, n_n241, n_n1059, n_n975, wire292, n_n1184, n_n1145, wire356, wire1384, wire1386, n_n554, n_n1188, wire694, wire868, wire869, n_n211, n_n1132, n_n1048, n_n980, n_n981, n_n1130, n_n983, wire354, n_n1117, wire303, n_n67, wire103, n_n76, n_n1177, wire5825, wire5826, n_n385, wire335, wire340, wire344, n_n1158, wire125, wire5903, n_n208, wire5338, n_n970, wire174, n_n966, wire1017, wire1018, wire464, wire465, wire466, wire307, wire5686, n_n1147, n_n950, wire1020, n_n652, n_n1173, n_n1088, wire5985, wire5986, wire5987, wire5990, wire5991, n_n261, n_n940, wire242, wire246, wire336, n_n995, wire1557, wire1558, n_n882, n_n986, wire296, n_n999, n_n1004, n_n1216, wire194, wire1311, wire306, n_n1055, n_n1009, wire4871, n_n1011, n_n1217, n_n1144, wire290, wire1146, wire5273, wire1501, wire1502, wire1503, wire332, wire333, n_n1001, n_n994, n_n1025, n_n976, n_n987, n_n953, wire5400, n_n990, n_n991, n_n1095, n_n1013, n_n1014, n_n1028, n_n1002, wire752, wire753, wire167, n_n1040, wire299, n_n1006, n_n1068, wire613, wire615, n_n296, n_n1146, n_n1010, n_n1020, wire249, n_n984, n_n978, wire4902, wire203, n_n1163, n_n1079, wire106, n_n1085, n_n1170, wire343, wire305, n_n1018, wire1005, wire1007, wire1008, wire289, wire1151, wire1153, wire1154, wire1001, wire1002, wire1003, wire309, n_n993, wire5396, wire4873, n_n1026, wire1102, wire286, wire1529, wire1531, n_n1070, n_n977, n_n1160, wire861, wire862, wire863, wire300, wire730, wire809, wire810, wire287, n_n1215, wire350, wire1504, wire5012, n_n955, wire353, wire5542, n_n1019, wire130, wire135, wire348, wire5993, wire60, wire69, wire165, wire382, wire383, wire384, wire385, wire386, wire387, wire388, wire389, wire390, wire391, wire392, wire393, wire394, wire395, wire5943, wire413, wire430, wire431, wire432, wire433, wire434, wire435, wire436, wire437, wire438, wire439, wire467, wire468, wire469, wire5847, wire475, wire476, wire477, wire478, wire479, wire480, wire481, wire482, wire483, wire484, wire485, wire5828, wire507, wire508, wire526, wire532, wire5783, wire559, wire562, wire596, wire611, wire5734, wire5709, wire617, wire618, wire619, wire620, wire621, wire5688, wire641, wire642, wire643, wire644, wire645, wire646, wire647, wire648, wire649, wire662, wire663, wire664, wire5661, wire666, wire668, wire669, wire670, wire671, wire690, wire692, wire693, wire696, wire5626, wire697, wire732, wire734, wire736, wire755, wire756, wire757, wire758, wire759, wire805, wire5558, wire807, wire808, wire812, wire5544, wire825, wire827, wire833, wire834, wire835, wire836, wire839, wire840, wire864, wire866, wire867, wire870, wire871, wire872, wire873, wire874, wire876, wire877, wire5498, wire878, wire895, wire897, wire899, wire900, wire901, wire5457, wire906, wire5458, wire907, wire5459, wire908, wire909, wire910, wire911, wire940, wire942, wire944, wire946, wire948, wire5444, wire950, wire957, wire958, wire959, wire960, wire961, wire962, wire963, wire5423, wire978, wire979, wire980, wire981, wire982, wire983, wire984, wire985, wire986, wire989, wire1009, wire1011, wire1012, wire5398, wire1013, wire1024, wire1039, wire5375, wire1041, wire1043, wire1046, wire1048, wire1080, wire1082, wire5319, wire1085, wire5318, wire5276, wire1106, wire5277, wire1107, wire5279, wire1108, wire1109, wire5281, wire1110, wire1111, wire1112, wire1113, wire1114, wire1115, wire1116, wire1117, wire1118, wire1119, wire1120, wire1123, wire1142, wire1143, wire1144, wire1145, wire1155, wire1156, wire1293, wire1294, wire5251, wire1157, wire1173, wire1175, wire1177, wire1179, wire1191, wire1192, wire1193, wire1194, wire1197, wire1213, wire1214, wire1215, wire1234, wire1235, wire5143, wire1253, wire1254, wire1255, wire1256, wire1257, wire1281, wire1283, wire1285, wire1286, wire1287, wire1288, wire5141, wire1289, wire1290, wire1291, wire1292, wire1295, wire1313, wire1317, wire1318, wire1319, wire1320, wire1350, wire1351, wire1352, wire1354, wire1356, wire1357, wire1358, wire1359, wire1360, wire1361, wire1362, wire1380, wire1381, wire1382, wire1383, wire1388, wire1389, wire1411, wire1413, wire1414, wire1415, wire1417, wire1421, wire1440, wire1443, wire4958, wire1445, wire4959, wire1446, wire1447, wire1448, wire1449, wire1450, wire1451, wire1452, wire4952, wire1483, wire1484, wire1485, wire1486, wire1487, wire1489, wire1490, wire1491, wire1499, wire1507, wire1508, wire4931, wire1509, wire1510, wire1511, wire4930, wire1520, wire1521, wire1522, wire1523, wire1524, wire1525, wire1527, wire4921, wire1533, wire1534, wire1535, wire1536, wire1559, wire1560, wire1562, wire1583, wire4841, wire1589, wire1590, wire1591, wire1592, wire1595, wire1596, wire1599, wire1600, wire1601, wire1602, wire1617, wire1618, wire1619, wire1620, wire1621, wire1622, wire1623, wire1624, wire4840, wire1625, wire1627, wire1628, wire1629, wire1631, wire4849, wire4851, wire4854, wire4855, wire4856, wire4857, wire4858, wire4859, wire4861, wire4875, wire4876, wire4877, wire4878, wire4887, wire4890, wire4891, wire4892, wire4893, wire4894, wire4895, wire4899, wire4900, wire4904, wire4910, wire4911, wire4912, wire4913, wire4914, wire4919, wire4920, wire4928, wire4929, wire4954, wire4955, wire4957, wire4960, wire4971, wire4972, wire4973, wire4974, wire4975, wire4976, wire4977, wire4978, wire4983, wire4984, wire4985, wire4997, wire5001, wire5002, wire5003, wire5004, wire5005, wire5006, wire5010, wire5011, wire5015, wire5020, wire5021, wire5022, wire5023, wire5024, wire5025, wire5029, wire5030, wire5036, wire5037, wire5038, wire5039, wire5040, wire5041, wire5057, wire5058, wire5059, wire5060, wire5061, wire5062, wire5072, wire5073, wire5074, wire5075, wire5076, wire5080, wire5081, wire5093, wire5094, wire5095, wire5096, wire5097, wire5098, wire5099, wire5100, wire5101, wire5106, wire5107, wire5117, wire5118, wire5119, wire5120, wire5121, wire5130, wire5131, wire5132, wire5133, wire5134, wire5139, wire5140, wire5150, wire5151, wire5152, wire5153, wire5154, wire5155, wire5156, wire5157, wire5158, wire5159, wire5164, wire5165, wire5176, wire5177, wire5178, wire5179, wire5180, wire5181, wire5185, wire5186, wire5191, wire5193, wire5194, wire5195, wire5196, wire5197, wire5198, wire5202, wire5203, wire5207, wire5208, wire5209, wire5210, wire5211, wire5212, wire5213, wire5214, wire5227, wire5230, wire5237, wire5239, wire5240, wire5241, wire5242, wire5243, wire5244, wire5257, wire5258, wire5259, wire5295, wire5296, wire5297, wire5298, wire5299, wire5300, wire5301, wire5302, wire5303, wire5304, wire5305, wire5326, wire5327, wire5328, wire5329, wire5330, wire5331, wire5335, wire5336, wire5340, wire5342, wire5353, wire5354, wire5355, wire5356, wire5357, wire5358, wire5359, wire5360, wire5367, wire5368, wire5379, wire5380, wire5381, wire5382, wire5383, wire5388, wire5389, wire5401, wire5412, wire5413, wire5414, wire5415, wire5416, wire5421, wire5422, wire5431, wire5432, wire5433, wire5434, wire5435, wire5436, wire5440, wire5441, wire5445, wire5470, wire5471, wire5472, wire5473, wire5474, wire5475, wire5476, wire5477, wire5478, wire5482, wire5483, wire5484, wire5502, wire5503, wire5504, wire5505, wire5506, wire5507, wire5508, wire5512, wire5513, wire5521, wire5523, wire5524, wire5525, wire5526, wire5527, wire5528, wire5529, wire5530, wire5537, wire5538, wire5547, wire5548, wire5549, wire5550, wire5551, wire5556, wire5557, wire5569, wire5570, wire5571, wire5572, wire5573, wire5574, wire5575, wire5576, wire5584, wire5585, wire5586, wire5587, wire5597, wire5598, wire5599, wire5600, wire5601, wire5605, wire5606, wire5613, wire5614, wire5615, wire5616, wire5617, wire5622, wire5623, wire5634, wire5635, wire5636, wire5637, wire5638, wire5639, wire5640, wire5641, wire5642, wire5643, wire5644, wire5645, wire5652, wire5653, wire5654, wire5655, wire5662, wire5668, wire5671, wire5672, wire5673, wire5674, wire5675, wire5676, wire5681, wire5682, wire5698, wire5699, wire5700, wire5701, wire5702, wire5703, wire5707, wire5708, wire5719, wire5720, wire5721, wire5722, wire5723, wire5724, wire5725, wire5730, wire5731, wire5741, wire5742, wire5743, wire5744, wire5748, wire5749, wire5750, wire5756, wire5758, wire5759, wire5760, wire5761, wire5762, wire5763, wire5764, wire5765, wire5766, wire5767, wire5768, wire5775, wire5776, wire5777, wire5787, wire5788, wire5789, wire5790, wire5791, wire5795, wire5796, wire5803, wire5804, wire5805, wire5806, wire5807, wire5808, wire5809, wire5815, wire5816, wire5817, wire5818, wire5833, wire5836, wire5837, wire5838, wire5839, wire5840, wire5841, wire5845, wire5846, wire5848, wire5858, wire5859, wire5860, wire5861, wire5862, wire5863, wire5864, wire5865, wire5866, wire5871, wire5872, wire5873, wire5886, wire5887, wire5888, wire5889, wire5890, wire5891, wire5892, wire5896, wire5897, wire5901, wire5902, wire5905, wire5907, wire5908, wire5919, wire5920, wire5921, wire5922, wire5923, wire5924, wire5925, wire5926, wire5927, wire5936, wire5937, wire5947, wire5948, wire5949, wire5950, wire5951, wire5952, wire5957, wire5958, wire5971, wire5972, wire5973, wire5974, wire5975, wire5976, wire5977, wire5978, wire5979, wire5989, wire5995, wire6006, wire6007, wire6008, wire6009, wire6010, wire6011, wire6012, wire6013, wire6014, wire6015, wire6016, wire6023, _19, _39, _41, _46, _48, _50, _57, _69, _83, _4857, _4863, _4865, _4879, _4881, _4906, _5158, _5183, _5226, _5523, _5553, _5615, _5644, _5645, _5668, _5724, _5729, _5732, _5733, _5783, _5786, _5980, _6026, _6079, _6088, _6101, _6140, _6161, _6190, _6228, _6248, _6319, _6325, _6345, _6353, _6357, _6358, _6359, _6377, _6430;

assign o_1_ = ( n_n110 ) | ( wire4865 ) | ( wire4866 ) | ( wire4867 ) ;
 assign o_2_ = ( wire4989 ) | ( wire4990 ) | ( wire4991 ) ;
 assign o_0_ =((~ i_7_) & i_7_);
 assign o_12_ = ( wire5046 ) | ( wire5047 ) | ( wire5049 ) ;
 assign o_11_ = ( wire5066 ) | ( wire5067 ) | ( wire5108 ) | ( wire5111 ) ;
 assign o_14_ = ( wire5125 ) | ( wire5126 ) | ( wire5166 ) | ( wire5169 ) ;
 assign o_13_ = ( wire5218 ) | ( wire5219 ) | ( wire5221 ) ;
 assign o_16_ = ( wire5228 ) | ( wire5229 ) | ( wire5233 ) ;
 assign o_15_ = ( wire5249 ) | ( wire5250 ) ;
 assign o_18_ = ( wire5260 ) | ( wire5261 ) | ( wire5265 ) ;
 assign o_17_ = ( wire5268 ) | ( wire5269 ) | ( wire5270 ) ;
 assign o_10_ = ( n_n655 ) | ( wire5369 ) | ( wire5370 ) | ( wire5373 ) ;
 assign o_9_ = ( n_n586 ) | ( wire5487 ) | ( wire5488 ) | ( wire5489 ) ;
 assign o_7_ = ( wire5540 ) | ( wire5590 ) | ( _6101 ) ;
 assign o_8_ = ( wire5658 ) | ( wire5684 ) | ( _6228 ) ;
 assign o_5_ = ( wire5733 ) | ( wire5780 ) | ( _6345 ) ;
 assign o_6_ = ( wire5821 ) | ( wire5822 ) | ( wire5875 ) | ( wire5876 ) ;
 assign o_3_ = ( wire5934 ) | ( wire5935 ) | ( wire5940 ) | ( wire5941 ) ;
 assign o_4_ = ( n_n243 ) | ( wire6024 ) | ( wire6025 ) | ( wire6028 ) ;
 assign n_n110 = ( n_n1164 ) | ( n_n1021 ) | ( wire4837 ) | ( wire4838 ) ;
 assign wire4865 = ( wire1595 ) | ( wire1596 ) | ( wire4849 ) | ( wire4859 ) ;
 assign wire4866 = ( wire1601 ) | ( wire1602 ) | ( wire4854 ) | ( wire4861 ) ;
 assign wire4867 = ( wire4855 ) | ( wire4856 ) | ( wire4857 ) | ( wire4858 ) ;
 assign wire4989 = ( wire4899 ) | ( wire4900 ) | ( wire4985 ) ;
 assign wire4990 = ( n_n137 ) | ( n_n135 ) | ( wire4919 ) | ( wire4920 ) ;
 assign wire4991 = ( n_n136 ) | ( n_n139 ) | ( wire4983 ) | ( wire4984 ) ;
 assign wire5046 = ( wire231 ) | ( wire301 ) | ( wire5036 ) | ( wire5037 ) ;
 assign wire5047 = ( wire5038 ) | ( wire5039 ) | ( wire5040 ) | ( wire5041 ) ;
 assign wire5049 = ( wire5010 ) | ( wire5011 ) | ( wire5029 ) | ( wire5030 ) ;
 assign wire5066 = ( n_n554 ) | ( wire5057 ) | ( wire5062 ) ;
 assign wire5067 = ( wire5058 ) | ( wire5059 ) | ( wire5060 ) | ( wire5061 ) ;
 assign wire5108 = ( wire5096 ) | ( wire5097 ) | ( wire5098 ) | ( wire5099 ) ;
 assign wire5111 = ( wire5080 ) | ( wire5081 ) | ( wire5106 ) | ( wire5107 ) ;
 assign wire5125 = ( n_n882 ) | ( wire296 ) | ( wire5121 ) ;
 assign wire5126 = ( wire5117 ) | ( wire5118 ) | ( wire5119 ) | ( wire5120 ) ;
 assign wire5166 = ( wire5154 ) | ( wire5155 ) | ( wire5156 ) | ( wire5157 ) ;
 assign wire5169 = ( wire5139 ) | ( wire5140 ) | ( wire5164 ) | ( wire5165 ) ;
 assign wire5218 = ( wire5208 ) | ( wire5209 ) | ( wire5214 ) ;
 assign wire5219 = ( wire5210 ) | ( wire5211 ) | ( wire5212 ) | ( wire5213 ) ;
 assign wire5221 = ( wire5185 ) | ( wire5186 ) | ( wire5202 ) | ( wire5203 ) ;
 assign wire5228 = ( n_n1109 ) | ( n_n1132 ) | ( wire1191 ) | ( wire1192 ) ;
 assign wire5229 = ( n_n1176 ) | ( wire135 ) | ( _5523 ) ;
 assign wire5233 = ( wire310 ) | ( wire5227 ) | ( wire5230 ) ;
 assign wire5249 = ( wire310 ) | ( wire302 ) | ( wire5239 ) | ( wire5240 ) ;
 assign wire5250 = ( wire5241 ) | ( wire5242 ) | ( wire5243 ) | ( wire5244 ) ;
 assign wire5260 = ( n_n1294 ) | ( n_n1169 ) | ( n_n942 ) | ( n_n1057 ) ;
 assign wire5261 = ( n_n1109 ) | ( n_n1125 ) | ( n_n1128 ) | ( n_n1286 ) ;
 assign wire5265 = ( wire302 ) | ( wire5257 ) | ( wire5258 ) | ( wire5259 ) ;
 assign wire5268 = ( n_n1109 ) | ( n_n1132 ) | ( wire1191 ) | ( wire1192 ) ;
 assign wire5269 = ( n_n941 ) | ( n_n955 ) | ( wire135 ) | ( wire1173 ) ;
 assign wire5270 = ( n_n1259 ) | ( n_n1176 ) | ( wire248 ) | ( n_n1283 ) ;
 assign n_n655 = ( n_n663 ) | ( wire5312 ) | ( wire5313 ) | ( wire5314 ) ;
 assign wire5369 = ( wire298 ) | ( wire5353 ) | ( wire5354 ) | ( wire5355 ) ;
 assign wire5370 = ( wire5356 ) | ( wire5357 ) | ( wire5358 ) | ( wire5359 ) ;
 assign wire5373 = ( wire5335 ) | ( wire5336 ) | ( wire5367 ) | ( wire5368 ) ;
 assign n_n586 = ( n_n324 ) | ( n_n397 ) | ( wire5403 ) ;
 assign wire5487 = ( wire5388 ) | ( wire5389 ) | ( wire5484 ) ;
 assign wire5488 = ( wire5421 ) | ( wire5422 ) | ( wire5440 ) | ( wire5441 ) ;
 assign wire5489 = ( n_n593 ) | ( n_n597 ) | ( wire5482 ) | ( wire5483 ) ;
 assign wire5540 = ( wire5512 ) | ( wire5513 ) | ( wire5538 ) ;
 assign wire5590 = ( wire5556 ) | ( wire5557 ) | ( wire5584 ) | ( wire5585 ) ;
 assign wire5658 = ( wire5622 ) | ( wire5623 ) | ( wire5652 ) | ( wire5653 ) ;
 assign wire5684 = ( wire5605 ) | ( wire5606 ) | ( wire5682 ) ;
 assign wire5733 = ( wire5707 ) | ( wire5708 ) | ( wire5731 ) ;
 assign wire5780 = ( n_n324 ) | ( wire5748 ) | ( wire5749 ) | ( wire5775 ) ;
 assign wire5821 = ( wire5795 ) | ( wire5796 ) | ( wire5818 ) ;
 assign wire5822 = ( n_n397 ) | ( wire5815 ) | ( wire5816 ) | ( wire5817 ) ;
 assign wire5875 = ( wire5872 ) | ( wire5873 ) ;
 assign wire5876 = ( n_n385 ) | ( wire5845 ) | ( wire5846 ) | ( wire5871 ) ;
 assign wire5934 = ( wire168 ) | ( n_n211 ) | ( wire5927 ) ;
 assign wire5935 = ( wire303 ) | ( wire307 ) | ( wire5919 ) | ( wire5920 ) ;
 assign wire5940 = ( wire5896 ) | ( wire5897 ) | ( wire5936 ) ;
 assign wire5941 = ( n_n208 ) | ( wire5907 ) | ( wire5908 ) | ( wire5937 ) ;
 assign n_n243 = ( wire5985 ) | ( wire5986 ) | ( wire5987 ) ;
 assign wire6024 = ( wire6009 ) | ( wire6010 ) | ( wire6011 ) | ( wire6012 ) ;
 assign wire6025 = ( wire6013 ) | ( wire6014 ) | ( wire6015 ) | ( wire6016 ) ;
 assign wire6028 = ( n_n261 ) | ( wire5957 ) | ( wire5958 ) | ( wire6023 ) ;
 assign n_n80 = ( (~ i_3_)  &  (~ i_2_)  &  i_0_ ) ;
 assign n_n75 = ( (~ i_7_)  &  i_8_ ) ;
 assign n_n81 = ( i_5_  &  i_3_  &  i_4_ ) ;
 assign n_n58 = ( i_7_  &  i_8_  &  (~ i_6_) ) ;
 assign n_n101 = ( i_7_  &  (~ i_8_)  &  i_6_ ) ;
 assign n_n93 = ( (~ i_7_)  &  (~ i_8_)  &  i_6_ ) ;
 assign n_n78 = ( (~ i_7_)  &  (~ i_8_)  &  (~ i_6_) ) ;
 assign n_n91 = ( (~ i_7_)  &  i_8_  &  i_6_ ) ;
 assign n_n99 = ( (~ i_5_)  &  (~ i_3_)  &  (~ i_4_) ) ;
 assign n_n103 = ( i_1_  &  i_2_  &  (~ i_0_) ) ;
 assign n_n1281 = ( n_n91  &  n_n99  &  n_n103 ) ;
 assign n_n100 = ( (~ i_1_)  &  (~ i_2_)  &  i_0_ ) ;
 assign n_n84 = ( (~ i_5_)  &  i_3_  &  (~ i_4_) ) ;
 assign n_n1185 = ( n_n78  &  n_n100  &  n_n84 ) ;
 assign n_n1164 = ( n_n93  &  n_n97  &  n_n96 ) ;
 assign n_n1021 = ( n_n96  &  n_n82  &  n_n85 ) ;
 assign wire4837 = ( n_n1134 ) | ( n_n1091 ) | ( wire1631 ) ;
 assign wire4838 = ( n_n1120 ) | ( n_n956 ) | ( n_n1156 ) | ( wire355 ) ;
 assign n_n97 = ( i_1_  &  i_2_  &  i_0_ ) ;
 assign n_n1174 = ( n_n93  &  n_n99  &  n_n97 ) ;
 assign wire172 = ( i_7_  &  (~ i_8_)  &  i_4_ ) ;
 assign wire192 = ( i_7_  &  (~ i_8_)  &  i_6_ ) | ( (~ i_7_)  &  i_8_  &  (~ i_6_) ) ;
 assign n_n96 = ( i_5_  &  (~ i_3_)  &  (~ i_4_) ) ;
 assign wire235 = ( n_n91  &  n_n97  &  n_n96 ) ;
 assign n_n92 = ( i_5_  &  i_3_  &  (~ i_4_) ) ;
 assign wire252 = ( n_n93  &  n_n103  &  n_n92 ) ;
 assign wire329 = ( n_n81  &  n_n101  &  n_n103 ) ;
 assign n_n74 = ( (~ i_5_)  &  (~ i_3_)  &  i_4_ ) ;
 assign n_n1077 = ( n_n91  &  n_n100  &  n_n74 ) ;
 assign n_n82 = ( i_7_  &  (~ i_8_)  &  (~ i_6_) ) ;
 assign n_n95 = ( i_7_  &  i_8_  &  i_6_ ) ;
 assign n_n90 = ( (~ i_1_)  &  i_2_  &  (~ i_0_) ) ;
 assign n_n1172 = ( n_n81  &  n_n95  &  n_n90 ) ;
 assign n_n1078 = ( n_n78  &  n_n99  &  n_n97 ) ;
 assign n_n54 = ( i_5_  &  (~ i_6_)  &  (~ i_4_) ) ;
 assign wire245 = ( i_3_  &  i_2_  &  i_0_ ) ;
 assign n_n1081 = ( i_7_  &  i_8_  &  n_n54  &  wire245 ) ;
 assign n_n1279 = ( n_n78  &  n_n74  &  n_n90 ) ;
 assign n_n1181 = ( n_n78  &  n_n96  &  n_n94 ) ;
 assign wire243 = ( n_n78  &  n_n103  &  n_n84 ) ;
 assign wire295 = ( n_n1204 ) | ( wire1529 ) | ( wire1531 ) ;
 assign wire4923 = ( wire1533 ) | ( wire1534 ) | ( wire1535 ) | ( wire1536 ) ;
 assign n_n137 = ( n_n1181 ) | ( wire243 ) | ( wire295 ) | ( wire4923 ) ;
 assign wire231 = ( wire1516 ) | ( wire1518 ) | ( wire1519 ) ;
 assign wire1512 = ( (~ i_7_)  &  i_8_  &  n_n81  &  n_n103 ) ;
 assign wire1513 = ( n_n93  &  n_n103  &  n_n77 ) ;
 assign wire4936 = ( wire340 ) | ( wire1509 ) | ( wire1510 ) | ( wire1511 ) ;
 assign n_n135 = ( wire231 ) | ( wire1512 ) | ( wire1513 ) | ( wire4936 ) ;
 assign n_n102 = ( (~ i_5_)  &  i_3_  &  i_4_ ) ;
 assign n_n1153 = ( n_n58  &  n_n90  &  n_n102 ) ;
 assign wire308 = ( wire1501 ) | ( wire1502 ) | ( wire1503 ) ;
 assign wire304 = ( wire349 ) | ( wire350 ) | ( wire1504 ) ;
 assign wire4942 = ( n_n1215 ) | ( wire1507 ) | ( wire1508 ) ;
 assign n_n136 = ( wire308 ) | ( wire304 ) | ( wire4942 ) ;
 assign n_n1297 = ( n_n96  &  n_n95  &  n_n90 ) ;
 assign n_n1324 = ( n_n93  &  n_n90  &  n_n102 ) ;
 assign n_n1092 = ( n_n91  &  n_n100  &  n_n84 ) ;
 assign n_n1108 = ( n_n81  &  n_n93  &  n_n90 ) ;
 assign n_n1105 = ( n_n81  &  n_n58  &  n_n94 ) ;
 assign wire4949 = ( n_n1100 ) | ( wire1491 ) | ( wire1499 ) ;
 assign wire4950 = ( n_n1103 ) | ( wire319 ) | ( n_n1130 ) | ( n_n1117 ) ;
 assign n_n139 = ( n_n1108 ) | ( n_n1105 ) | ( wire4949 ) | ( wire4950 ) ;
 assign wire127 = ( i_6_  &  (~ i_3_)  &  i_4_ ) ;
 assign n_n83 = ( (~ i_1_)  &  i_2_  &  i_0_ ) ;
 assign wire35 = ( n_n96  &  n_n38 ) | ( n_n75  &  n_n40 ) ;
 assign wire1477 = ( (~ i_3_)  &  (~ i_1_)  &  i_0_  &  wire4952 ) ;
 assign wire1479 = ( i_7_  &  (~ i_6_)  &  n_n103  &  n_n102 ) ;
 assign wire232 = ( wire1477 ) | ( wire1479 ) | ( n_n83  &  wire35 ) ;
 assign n_n63 = ( (~ i_7_)  &  i_8_  &  (~ i_6_) ) ;
 assign n_n77 = ( i_5_  &  (~ i_3_)  &  i_4_ ) ;
 assign wire251 = ( n_n103  &  n_n63  &  n_n77 ) ;
 assign wire321 = ( n_n101  &  n_n97  &  n_n74 ) ;
 assign n_n1254 = ( n_n78  &  n_n92  &  n_n90 ) ;
 assign n_n1259 = ( n_n92  &  n_n90  &  n_n63 ) ;
 assign n_n1204 = ( n_n100  &  n_n96  &  n_n95 ) ;
 assign wire4994 = ( (~ i_7_)  &  i_8_  &  (~ i_5_)  &  (~ i_6_) ) ;
 assign n_n1369 = ( (~ i_3_)  &  (~ i_1_)  &  (~ i_0_)  &  wire4994 ) ;
 assign wire1516 = ( i_7_  &  i_8_  &  n_n54  &  wire4930 ) ;
 assign wire1518 = ( n_n99  &  n_n82  &  n_n85 ) ;
 assign wire1519 = ( n_n58  &  n_n100  &  n_n77 ) ;
 assign wire1408 = ( n_n92  &  n_n95  &  n_n85 ) ;
 assign wire1409 = ( n_n93  &  n_n100  &  n_n102 ) ;
 assign wire1410 = ( n_n91  &  n_n99  &  n_n83 ) ;
 assign wire301 = ( wire1408 ) | ( wire1409 ) | ( wire1410 ) ;
 assign n_n85 = ( i_1_  &  (~ i_2_)  &  i_0_ ) ;
 assign wire314 = ( n_n78  &  n_n102  &  n_n85 ) ;
 assign wire349 = ( n_n81  &  n_n58  &  n_n103 ) ;
 assign n_n1022 = ( n_n58  &  n_n102  &  n_n85 ) ;
 assign n_n1134 = ( n_n58  &  n_n100  &  n_n74 ) ;
 assign n_n94 = ( i_1_  &  (~ i_2_)  &  (~ i_0_) ) ;
 assign n_n1039 = ( n_n78  &  n_n102  &  n_n94 ) ;
 assign wire241 = ( i_3_  &  (~ i_2_)  &  i_0_ ) ;
 assign n_n87 = ( i_5_  &  (~ i_6_)  &  i_4_ ) ;
 assign n_n1091 = ( i_7_  &  i_8_  &  wire241  &  n_n87 ) ;
 assign wire322 = ( (~ i_3_)  &  i_2_  &  (~ i_0_) ) ;
 assign n_n1093 = ( (~ i_7_)  &  i_8_  &  n_n54  &  wire322 ) ;
 assign n_n1103 = ( n_n95  &  n_n102  &  n_n83 ) ;
 assign n_n1120 = ( n_n92  &  n_n95  &  n_n83 ) ;
 assign n_n1052 = ( n_n74  &  n_n63  &  n_n94 ) ;
 assign n_n1331 = ( n_n91  &  n_n74  &  n_n90 ) ;
 assign n_n38 = ( i_7_  &  (~ i_6_) ) ;
 assign n_n40 = ( (~ i_5_)  &  (~ i_6_)  &  i_4_ ) ;
 assign wire177 = ( (~ i_7_)  &  i_8_  &  i_6_ ) | ( i_7_  &  (~ i_8_)  &  i_6_ ) ;
 assign n_n1109 = ( n_n101  &  n_n74  &  n_n90 ) ;
 assign wire1345 = ( i_7_  &  i_6_  &  n_n97  &  n_n77 ) ;
 assign wire1348 = ( (~ i_7_)  &  (~ i_6_)  &  n_n99  &  n_n100 ) ;
 assign wire257 = ( n_n1078 ) | ( n_n1109 ) | ( wire1345 ) | ( wire1348 ) ;
 assign n_n1193 = ( n_n58  &  n_n84  &  n_n94 ) ;
 assign n_n1330 = ( n_n95  &  n_n90  &  n_n102 ) ;
 assign n_n1267 = ( n_n101  &  n_n100  &  n_n84 ) ;
 assign wire342 = ( (~ i_7_)  &  (~ i_6_)  &  n_n77  &  n_n94 ) ;
 assign wire346 = ( n_n100  &  n_n74  &  n_n82 ) ;
 assign wire323 = ( n_n99  &  n_n82  &  n_n94 ) ;
 assign wire352 = ( n_n78  &  n_n96  &  n_n90 ) ;
 assign wire357 = ( n_n101  &  n_n103  &  n_n96 ) ;
 assign n_n1176 = ( n_n91  &  n_n74  &  n_n94 ) ;
 assign n_n1074 = ( n_n101  &  n_n74  &  n_n94 ) ;
 assign n_n1032 = ( n_n93  &  n_n74  &  n_n90 ) ;
 assign n_n1294 = ( n_n78  &  n_n84  &  n_n90 ) ;
 assign n_n1312 = ( n_n101  &  n_n96  &  n_n90 ) ;
 assign wire326 = ( n_n101  &  n_n77  &  n_n94 ) ;
 assign wire5222 = ( n_n91  &  n_n96  &  n_n90 ) | ( n_n96  &  n_n95  &  n_n90 ) ;
 assign wire310 = ( n_n1312 ) | ( wire326 ) | ( wire5222 ) ;
 assign n_n1169 = ( n_n91  &  n_n90  &  n_n102 ) ;
 assign n_n942 = ( n_n91  &  n_n92  &  n_n94 ) ;
 assign n_n1057 = ( n_n81  &  n_n82  &  n_n90 ) ;
 assign n_n1125 = ( n_n81  &  n_n78  &  n_n90 ) ;
 assign n_n1128 = ( n_n78  &  n_n84  &  n_n94 ) ;
 assign wire248 = ( n_n95  &  n_n77  &  n_n94 ) ;
 assign n_n1046 = ( n_n101  &  n_n90  &  n_n102 ) ;
 assign n_n1042 = ( n_n93  &  n_n92  &  n_n94 ) ;
 assign n_n1047 = ( n_n81  &  n_n90  &  n_n63 ) ;
 assign wire302 = ( n_n1039 ) | ( n_n1046 ) | ( n_n1042 ) | ( n_n1047 ) ;
 assign n_n1286 = ( n_n58  &  n_n92  &  n_n94 ) ;
 assign n_n79 = ( (~ i_5_)  &  (~ i_6_)  &  (~ i_4_) ) ;
 assign n_n937 = ( (~ i_1_)  &  (~ i_2_)  &  (~ i_0_) ) ;
 assign wire351 = ( (~ i_3_)  &  (~ i_1_)  &  (~ i_0_) ) ;
 assign wire189 = ( n_n937 ) | ( n_n79  &  wire351 ) ;
 assign n_n1283 = ( n_n91  &  n_n96  &  n_n90 ) ;
 assign n_n1087 = ( n_n81  &  n_n63  &  n_n94 ) ;
 assign n_n663 = ( n_n1294 ) | ( wire290 ) | ( wire1146 ) | ( wire5273 ) ;
 assign wire5312 = ( wire308 ) | ( wire5295 ) | ( wire5296 ) | ( wire5297 ) ;
 assign wire5313 = ( wire5298 ) | ( wire5299 ) | ( wire5300 ) | ( wire5301 ) ;
 assign wire5314 = ( wire5302 ) | ( wire5303 ) | ( wire5304 ) | ( wire5305 ) ;
 assign n_n71 = ( (~ i_5_)  &  i_6_  &  (~ i_4_) ) ;
 assign n_n968 = ( i_7_  &  (~ i_8_)  &  n_n80  &  n_n71 ) ;
 assign n_n958 = ( n_n95  &  n_n77  &  n_n85 ) ;
 assign n_n66 = ( i_5_  &  i_6_  &  (~ i_4_) ) ;
 assign n_n974 = ( i_7_  &  (~ i_8_)  &  n_n83  &  n_n66 ) ;
 assign n_n973 = ( n_n103  &  n_n74  &  n_n82 ) ;
 assign n_n989 = ( n_n81  &  n_n91  &  n_n94 ) ;
 assign n_n64 = ( i_7_  &  i_8_ ) ;
 assign n_n938 = ( n_n101  &  n_n103  &  n_n102 ) ;
 assign n_n944 = ( n_n91  &  n_n97  &  n_n102 ) ;
 assign n_n70 = ( i_7_  &  (~ i_8_) ) ;
 assign n_n982 = ( n_n81  &  n_n93  &  n_n83 ) ;
 assign n_n967 = ( n_n93  &  n_n100  &  n_n77 ) ;
 assign n_n956 = ( n_n78  &  n_n97  &  n_n96 ) ;
 assign n_n1121 = ( i_5_  &  i_6_  &  wire172  &  n_n90 ) ;
 assign n_n53 = ( (~ i_3_)  &  i_1_  &  i_2_ ) ;
 assign wire4880 = ( (~ i_5_)  &  (~ i_3_) ) ;
 assign wire4881 = ( (~ i_7_)  &  (~ i_6_)  &  i_1_  &  (~ i_2_) ) ;
 assign wire70 = ( n_n80  &  n_n40 ) | ( wire4880  &  wire4881 ) ;
 assign n_n962 = ( n_n78  &  n_n74  &  n_n83 ) ;
 assign n_n961 = ( n_n100  &  n_n95  &  n_n102 ) ;
 assign n_n964 = ( n_n99  &  n_n95  &  n_n94 ) ;
 assign wire168 = ( n_n962 ) | ( n_n961 ) | ( n_n964 ) ;
 assign wire236 = ( i_7_  &  i_8_  &  n_n100  &  n_n87 ) ;
 assign n_n941 = ( n_n93  &  n_n96  &  n_n94 ) ;
 assign n_n949 = ( n_n101  &  n_n84  &  n_n85 ) ;
 assign n_n943 = ( n_n93  &  n_n92  &  n_n90 ) ;
 assign wire291 = ( n_n941 ) | ( n_n949 ) | ( n_n943 ) ;
 assign n_n954 = ( n_n81  &  n_n78  &  n_n94 ) ;
 assign n_n952 = ( n_n81  &  n_n82  &  n_n85 ) ;
 assign n_n951 = ( n_n92  &  n_n82  &  n_n83 ) ;
 assign wire297 = ( n_n954 ) | ( n_n952 ) | ( n_n951 ) ;
 assign n_n960 = ( (~ i_7_)  &  i_8_  &  n_n85  &  n_n76 ) ;
 assign n_n959 = ( n_n91  &  n_n84  &  n_n97 ) ;
 assign n_n957 = ( n_n91  &  n_n100  &  n_n92 ) ;
 assign wire298 = ( n_n960 ) | ( n_n959 ) | ( n_n957 ) ;
 assign wire319 = ( (~ i_7_)  &  (~ i_6_)  &  n_n90  &  n_n77 ) ;
 assign n_n1082 = ( n_n97  &  n_n74  &  n_n63 ) ;
 assign n_n324 = ( wire297 ) | ( n_n960 ) | ( n_n957 ) | ( wire303 ) ;
 assign n_n397 = ( n_n941 ) | ( n_n943 ) | ( wire125 ) | ( wire5400 ) ;
 assign wire5403 = ( wire168 ) | ( n_n652 ) | ( wire5401 ) ;
 assign n_n1045 = ( i_8_  &  (~ i_6_)  &  n_n84  &  n_n94 ) ;
 assign n_n1043 = ( n_n91  &  n_n102  &  n_n85 ) ;
 assign n_n1122 = ( n_n101  &  n_n99  &  n_n94 ) ;
 assign n_n1036 = ( n_n91  &  n_n103  &  n_n74 ) ;
 assign n_n1118 = ( (~ i_7_)  &  i_8_  &  n_n90  &  wire127 ) ;
 assign n_n1030 = ( n_n81  &  n_n82  &  n_n83 ) ;
 assign wire5442 = ( i_6_  &  i_3_  &  (~ i_4_) ) ;
 assign n_n1083 = ( i_7_  &  i_8_  &  n_n103  &  wire5442 ) ;
 assign n_n1101 = ( i_7_  &  (~ i_8_)  &  n_n54  &  wire322 ) ;
 assign n_n1156 = ( n_n91  &  n_n99  &  n_n94 ) ;
 assign wire5448 = ( wire957 ) | ( wire958 ) | ( wire353  &  wire5445 ) ;
 assign wire5449 = ( wire251 ) | ( wire335 ) | ( wire950 ) | ( wire1440 ) ;
 assign n_n593 = ( n_n1128 ) | ( n_n1156 ) | ( wire5448 ) | ( wire5449 ) ;
 assign n_n1060 = ( n_n103  &  n_n74  &  n_n63 ) ;
 assign wire1104 = ( (~ i_5_)  &  (~ i_6_)  &  i_4_  &  wire5318 ) ;
 assign wire5452 = ( n_n1058 ) | ( n_n1059 ) | ( wire1354 ) ;
 assign wire5453 = ( n_n1052 ) | ( n_n1057 ) | ( n_n1055 ) | ( wire948 ) ;
 assign n_n597 = ( n_n1060 ) | ( wire1104 ) | ( wire5452 ) | ( wire5453 ) ;
 assign wire355 = ( (~ i_7_)  &  (~ i_6_)  &  n_n81  &  n_n83 ) ;
 assign n_n1100 = ( n_n100  &  n_n82  &  n_n77 ) ;
 assign n_n969 = ( n_n93  &  n_n83  &  n_n77 ) ;
 assign n_n939 = ( (~ i_8_)  &  (~ i_6_)  &  n_n99  &  n_n100 ) ;
 assign wire131 = ( (~ i_6_)  &  (~ i_3_)  &  (~ i_4_) ) ;
 assign n_n971 = ( (~ i_7_)  &  (~ i_8_)  &  n_n100  &  wire131 ) ;
 assign n_n1035 = ( n_n101  &  n_n74  &  n_n85 ) ;
 assign n_n1037 = ( (~ i_8_)  &  i_6_  &  n_n102  &  n_n94 ) ;
 assign wire334 = ( n_n78  &  n_n99  &  n_n103 ) ;
 assign wire345 = ( n_n99  &  n_n95  &  n_n83 ) ;
 assign wire903 = ( i_7_  &  i_8_  &  n_n103  &  n_n40 ) ;
 assign n_n421 = ( wire334 ) | ( wire345 ) | ( wire903 ) ;
 assign n_n1058 = ( n_n58  &  n_n74  &  n_n94 ) ;
 assign n_n947 = ( (~ i_3_)  &  (~ i_0_)  &  n_n87  &  wire5396 ) ;
 assign wire831 = ( n_n97  &  n_n95  &  n_n102 ) ;
 assign wire5541 = ( (~ i_8_)  &  i_6_  &  i_3_  &  (~ i_4_) ) ;
 assign n_n241 = ( n_n947 ) | ( wire831 ) | ( n_n97  &  wire5541 ) ;
 assign n_n1059 = ( (~ i_7_)  &  (~ i_8_)  &  wire245  &  n_n71 ) ;
 assign n_n975 = ( n_n101  &  n_n84  &  n_n83 ) ;
 assign wire292 = ( n_n968 ) | ( n_n973 ) | ( n_n975 ) ;
 assign n_n1184 = ( n_n84  &  n_n95  &  n_n94 ) ;
 assign n_n1145 = ( (~ i_6_)  &  i_3_  &  wire172  &  n_n94 ) ;
 assign wire356 = ( n_n93  &  n_n102  &  n_n85 ) ;
 assign wire1384 = ( i_8_  &  (~ i_6_)  &  n_n81  &  n_n85 ) ;
 assign wire1386 = ( n_n93  &  n_n84  &  n_n94 ) ;
 assign n_n554 = ( wire356 ) | ( wire1384 ) | ( wire1386 ) ;
 assign n_n1188 = ( n_n81  &  n_n58  &  n_n90 ) ;
 assign wire694 = ( n_n58  &  n_n99  &  n_n94 ) ;
 assign wire868 = ( n_n81  &  n_n100  &  n_n95 ) ;
 assign wire869 = ( n_n82  &  n_n90  &  n_n102 ) ;
 assign n_n211 = ( wire694 ) | ( wire868 ) | ( wire869 ) ;
 assign n_n1132 = ( n_n93  &  n_n96  &  n_n90 ) ;
 assign n_n1048 = ( n_n96  &  n_n95  &  n_n94 ) ;
 assign n_n980 = ( n_n84  &  n_n82  &  n_n83 ) ;
 assign n_n981 = ( n_n84  &  n_n95  &  n_n85 ) ;
 assign n_n1130 = ( n_n58  &  n_n84  &  n_n85 ) ;
 assign n_n983 = ( n_n99  &  n_n100  &  n_n95 ) ;
 assign wire354 = ( (~ i_5_)  &  (~ i_6_)  &  i_3_ ) ;
 assign n_n1117 = ( i_7_  &  (~ i_8_)  &  n_n94  &  wire354 ) ;
 assign wire303 = ( n_n967 ) | ( n_n966 ) | ( wire1017 ) | ( wire1018 ) ;
 assign n_n67 = ( (~ i_3_)  &  (~ i_1_)  &  i_0_ ) ;
 assign wire103 = ( n_n83  &  n_n66  &  n_n70 ) | ( n_n66  &  n_n70  &  n_n67 ) ;
 assign n_n76 = ( i_5_  &  (~ i_6_)  &  i_3_ ) ;
 assign n_n1177 = ( n_n78  &  n_n92  &  n_n94 ) ;
 assign wire5825 = ( n_n1125 ) | ( wire526 ) | ( wire1082 ) ;
 assign wire5826 = ( n_n1121 ) | ( wire734 ) | ( wire1144 ) | ( wire1145 ) ;
 assign n_n385 = ( n_n1153 ) | ( wire251 ) | ( wire5825 ) | ( wire5826 ) ;
 assign wire335 = ( n_n81  &  n_n97  &  n_n82 ) ;
 assign wire340 = ( n_n91  &  n_n92  &  n_n85 ) ;
 assign wire344 = ( n_n93  &  n_n103  &  n_n84 ) ;
 assign n_n1158 = ( n_n78  &  n_n103  &  n_n96 ) ;
 assign wire125 = ( n_n942 ) | ( n_n938 ) | ( n_n940 ) ;
 assign wire5903 = ( n_n958 ) | ( n_n952 ) | ( n_n953 ) ;
 assign n_n208 = ( n_n241 ) | ( wire125 ) | ( wire5903 ) ;
 assign wire5338 = ( i_5_  &  i_6_  &  i_4_ ) ;
 assign n_n970 = ( (~ i_7_)  &  i_8_  &  n_n85  &  wire5338 ) ;
 assign wire174 = ( i_3_  &  (~ i_1_)  &  i_2_ ) ;
 assign n_n966 = ( n_n101  &  n_n97  &  n_n102 ) ;
 assign wire1017 = ( i_8_  &  i_6_  &  n_n103  &  n_n77 ) ;
 assign wire1018 = ( (~ i_7_)  &  (~ i_6_)  &  n_n102  &  n_n85 ) ;
 assign wire464 = ( i_7_  &  i_8_  &  n_n103  &  wire130 ) ;
 assign wire465 = ( n_n93  &  n_n102  &  n_n83 ) ;
 assign wire466 = ( n_n81  &  n_n58  &  n_n97 ) ;
 assign wire307 = ( wire464 ) | ( wire465 ) | ( wire466 ) ;
 assign wire5686 = ( (~ i_7_)  &  (~ i_8_)  &  (~ i_3_) ) ;
 assign n_n1147 = ( i_1_  &  (~ i_2_)  &  n_n87  &  wire5686 ) ;
 assign n_n950 = ( n_n103  &  n_n95  &  n_n102 ) ;
 assign wire1020 = ( n_n97  &  n_n95  &  n_n102 ) ;
 assign n_n652 = ( n_n949 ) | ( n_n950 ) | ( wire1020 ) ;
 assign n_n1173 = ( n_n91  &  n_n103  &  n_n96 ) ;
 assign n_n1088 = ( n_n91  &  n_n97  &  n_n92 ) ;
 assign wire5985 = ( wire307 ) | ( wire300 ) | ( wire5979 ) ;
 assign wire5986 = ( wire5971 ) | ( wire5972 ) | ( wire5973 ) | ( wire5974 ) ;
 assign wire5987 = ( wire5975 ) | ( wire5976 ) | ( wire5977 ) | ( wire5978 ) ;
 assign wire5990 = ( n_n981 ) | ( n_n994 ) | ( n_n978 ) | ( wire1043 ) ;
 assign wire5991 = ( n_n999 ) | ( wire613 ) | ( wire615 ) | ( wire5989 ) ;
 assign n_n261 = ( wire5990 ) | ( wire5991 ) ;
 assign n_n940 = ( n_n97  &  n_n96  &  n_n95 ) ;
 assign wire242 = ( i_3_  &  i_2_  &  (~ i_0_) ) ;
 assign wire246 = ( n_n91  &  n_n103  &  n_n84 ) ;
 assign wire336 = ( n_n84  &  n_n97  &  n_n95 ) ;
 assign n_n995 = ( n_n100  &  n_n74  &  n_n95 ) ;
 assign wire1557 = ( n_n81  &  n_n101  &  n_n90 ) ;
 assign wire1558 = ( n_n78  &  n_n97  &  n_n102 ) ;
 assign n_n882 = ( n_n995 ) | ( wire1557 ) | ( wire1558 ) ;
 assign n_n986 = ( n_n92  &  n_n63  &  n_n94 ) ;
 assign wire296 = ( n_n980 ) | ( n_n983 ) | ( n_n986 ) ;
 assign n_n999 = ( n_n93  &  n_n103  &  n_n96 ) ;
 assign n_n1004 = ( n_n91  &  n_n97  &  n_n74 ) ;
 assign n_n1216 = ( n_n101  &  n_n100  &  n_n74 ) ;
 assign wire194 = ( i_5_  &  (~ i_3_)  &  i_4_ ) | ( (~ i_5_)  &  i_3_  &  (~ i_4_) ) ;
 assign wire1311 = ( n_n97  &  n_n92  &  n_n63 ) ;
 assign wire306 = ( n_n1174 ) | ( n_n1177 ) | ( wire1311 ) ;
 assign n_n1055 = ( n_n58  &  n_n96  &  n_n94 ) ;
 assign n_n1009 = ( n_n81  &  n_n103  &  n_n95 ) ;
 assign wire4871 = ( i_5_  &  i_6_  &  (~ i_3_) ) ;
 assign n_n1011 = ( i_7_  &  i_8_  &  n_n103  &  wire4871 ) ;
 assign n_n1217 = ( n_n101  &  n_n103  &  n_n74 ) ;
 assign n_n1144 = ( (~ i_7_)  &  i_8_  &  n_n79  &  wire174 ) ;
 assign wire290 = ( wire1151 ) | ( wire1153 ) | ( wire1154 ) ;
 assign wire1146 = ( (~ i_7_)  &  (~ i_8_)  &  wire241  &  n_n40 ) ;
 assign wire5273 = ( wire1155 ) | ( wire1156 ) | ( wire1358 ) | ( wire1359 ) ;
 assign wire1501 = ( (~ i_7_)  &  i_8_  &  n_n85  &  n_n87 ) ;
 assign wire1502 = ( i_7_  &  (~ i_8_)  &  n_n92  &  n_n85 ) ;
 assign wire1503 = ( (~ i_7_)  &  (~ i_8_)  &  n_n84  &  n_n85 ) ;
 assign wire332 = ( n_n74  &  n_n95  &  n_n90 ) ;
 assign wire333 = ( i_7_  &  i_6_  &  n_n92  &  n_n94 ) ;
 assign n_n1001 = ( n_n99  &  n_n97  &  n_n63 ) ;
 assign n_n994 = ( n_n91  &  n_n103  &  n_n102 ) ;
 assign n_n1025 = ( n_n74  &  n_n82  &  n_n83 ) ;
 assign n_n976 = ( (~ i_7_)  &  i_6_  &  n_n74  &  n_n85 ) ;
 assign n_n987 = ( n_n93  &  n_n97  &  n_n102 ) ;
 assign n_n953 = ( (~ i_7_)  &  (~ i_8_)  &  n_n80  &  n_n79 ) ;
 assign wire5400 = ( n_n944 ) | ( n_n939 ) | ( n_n947 ) | ( wire1013 ) ;
 assign n_n990 = ( n_n74  &  n_n95  &  n_n83 ) ;
 assign n_n991 = ( n_n81  &  n_n103  &  n_n82 ) ;
 assign n_n1095 = ( n_n91  &  n_n103  &  n_n92 ) ;
 assign n_n1013 = ( n_n93  &  n_n99  &  n_n103 ) ;
 assign n_n1014 = ( n_n81  &  n_n78  &  n_n100 ) ;
 assign n_n1028 = ( n_n97  &  n_n63  &  n_n77 ) ;
 assign n_n1002 = ( (~ i_7_)  &  i_8_  &  wire245  &  n_n79 ) ;
 assign wire752 = ( i_7_  &  i_8_  &  n_n74  &  n_n85 ) ;
 assign wire753 = ( (~ i_7_)  &  (~ i_8_)  &  n_n85  &  n_n76 ) ;
 assign wire167 = ( n_n1002 ) | ( wire752 ) | ( wire753 ) ;
 assign n_n1040 = ( n_n96  &  n_n95  &  n_n85 ) ;
 assign wire299 = ( n_n1039 ) | ( n_n1032 ) | ( n_n1042 ) | ( n_n1040 ) ;
 assign n_n1006 = ( n_n74  &  n_n95  &  n_n94 ) ;
 assign n_n1068 = ( n_n99  &  n_n95  &  n_n85 ) ;
 assign wire613 = ( n_n81  &  n_n101  &  n_n90 ) ;
 assign wire615 = ( n_n83  &  (~ n_n76)  &  wire5734 ) ;
 assign n_n296 = ( n_n999 ) | ( wire613 ) | ( wire615 ) ;
 assign n_n1146 = ( n_n101  &  n_n96  &  n_n85 ) ;
 assign n_n1010 = ( n_n78  &  n_n84  &  n_n97 ) ;
 assign n_n1020 = ( i_6_  &  i_3_  &  wire172  &  n_n94 ) ;
 assign wire249 = ( i_7_  &  i_6_  &  n_n81  &  n_n97 ) ;
 assign n_n984 = ( n_n103  &  n_n102  &  n_n63 ) ;
 assign n_n978 = ( n_n92  &  n_n83  &  n_n63 ) ;
 assign wire4902 = ( (~ i_7_)  &  i_5_  &  (~ i_6_)  &  i_3_ ) ;
 assign wire203 = ( n_n97  &  wire4902 ) | ( n_n91  &  n_n97  &  n_n74 ) ;
 assign n_n1163 = ( n_n91  &  n_n84  &  n_n83 ) ;
 assign n_n1079 = ( n_n81  &  n_n93  &  n_n100 ) ;
 assign wire106 = ( wire1479 ) | ( n_n83  &  wire35 ) ;
 assign n_n1085 = ( n_n102  &  n_n63  &  n_n94 ) ;
 assign n_n1170 = ( n_n93  &  n_n100  &  n_n92 ) ;
 assign wire343 = ( n_n101  &  n_n103  &  n_n92 ) ;
 assign wire305 = ( n_n989 ) | ( n_n987 ) | ( n_n991 ) | ( n_n984 ) ;
 assign n_n1018 = ( n_n100  &  n_n95  &  n_n77 ) ;
 assign wire1005 = ( n_n81  &  n_n93  &  n_n85 ) ;
 assign wire1007 = ( n_n91  &  n_n100  &  n_n102 ) ;
 assign wire1008 = ( n_n93  &  n_n99  &  n_n85 ) ;
 assign wire289 = ( wire1005 ) | ( wire1007 ) | ( wire1008 ) ;
 assign wire1151 = ( n_n100  &  n_n84  &  n_n82 ) ;
 assign wire1153 = ( n_n78  &  n_n90  &  n_n102 ) ;
 assign wire1154 = ( n_n93  &  n_n74  &  n_n94 ) ;
 assign wire1001 = ( n_n93  &  n_n103  &  n_n74 ) ;
 assign wire1002 = ( n_n90  &  n_n102  &  n_n63 ) ;
 assign wire1003 = ( n_n93  &  n_n90  &  n_n77 ) ;
 assign wire309 = ( wire352 ) | ( wire1001 ) | ( wire1002 ) | ( wire1003 ) ;
 assign n_n993 = ( (~ i_7_)  &  i_6_  &  n_n81  &  n_n103 ) ;
 assign wire5396 = ( (~ i_7_)  &  (~ i_8_)  &  i_1_ ) ;
 assign wire4873 = ( (~ i_3_)  &  i_1_  &  (~ i_0_) ) ;
 assign n_n1026 = ( i_7_  &  (~ i_8_)  &  n_n71  &  wire4873 ) ;
 assign wire1102 = ( i_7_  &  (~ i_8_)  &  n_n100  &  n_n54 ) ;
 assign wire286 = ( n_n1011 ) | ( n_n1006 ) | ( wire1102 ) ;
 assign wire1529 = ( n_n91  &  n_n102  &  n_n94 ) ;
 assign wire1531 = ( n_n81  &  n_n95  &  n_n94 ) ;
 assign n_n1070 = ( n_n93  &  n_n99  &  n_n94 ) ;
 assign n_n977 = ( i_7_  &  i_8_  &  n_n79  &  n_n67 ) ;
 assign n_n1160 = ( n_n81  &  n_n101  &  n_n83 ) ;
 assign wire861 = ( n_n91  &  n_n100  &  n_n96 ) ;
 assign wire862 = ( n_n101  &  n_n100  &  n_n92 ) ;
 assign wire863 = ( n_n81  &  n_n91  &  n_n83 ) ;
 assign wire300 = ( wire861 ) | ( wire862 ) | ( wire863 ) ;
 assign wire730 = ( (~ i_8_)  &  i_6_  &  n_n97  &  n_n92 ) ;
 assign wire809 = ( i_7_  &  (~ i_8_)  &  n_n97  &  n_n87 ) ;
 assign wire810 = ( i_7_  &  i_8_  &  n_n54  &  n_n85 ) ;
 assign wire287 = ( wire730 ) | ( wire809 ) | ( wire810 ) ;
 assign n_n1215 = ( n_n58  &  n_n100  &  n_n96 ) ;
 assign wire350 = ( n_n101  &  n_n100  &  n_n77 ) ;
 assign wire1504 = ( n_n101  &  n_n99  &  n_n97 ) ;
 assign wire5012 = ( (~ i_5_)  &  i_6_  &  (~ i_3_)  &  (~ i_4_) ) ;
 assign n_n955 = ( (~ i_1_)  &  i_2_  &  (~ i_0_)  &  wire5012 ) ;
 assign wire353 = ( (~ i_3_)  &  (~ i_1_)  &  i_2_ ) ;
 assign wire5542 = ( i_7_  &  i_8_  &  i_6_ ) ;
 assign n_n1019 = ( (~ i_5_)  &  i_4_  &  n_n85  &  wire5542 ) ;
 assign wire130 = ( (~ i_5_)  &  (~ i_6_)  &  (~ i_3_) ) ;
 assign wire135 = ( (~ i_1_)  &  (~ i_2_)  &  (~ i_0_) ) | ( (~ i_1_)  &  (~ i_0_)  &  wire131 ) ;
 assign wire348 = ( n_n78  &  n_n100  &  n_n77 ) ;
 assign wire5993 = ( i_7_  &  (~ i_8_)  &  (~ i_6_)  &  (~ i_4_) ) ;
 assign wire60 = ( i_3_  &  i_2_  &  (~ i_0_)  &  wire5993 ) ;
 assign wire69 = ( (~ i_7_)  &  i_6_  &  n_n99  &  n_n83 ) ;
 assign wire165 = ( i_7_  &  (~ i_8_)  &  n_n102  &  n_n85 ) ;
 assign wire382 = ( i_7_  &  (~ i_8_)  &  n_n85  &  n_n40 ) ;
 assign wire383 = ( (~ i_7_)  &  i_8_  &  n_n80  &  n_n54 ) ;
 assign wire384 = ( (~ i_7_)  &  (~ i_8_)  &  n_n103  &  wire130 ) ;
 assign wire385 = ( (~ i_7_)  &  (~ i_8_)  &  n_n81  &  n_n103 ) ;
 assign wire386 = ( i_7_  &  i_8_  &  n_n100  &  n_n76 ) ;
 assign wire387 = ( n_n103  &  n_n77  &  wire177 ) ;
 assign wire388 = ( (~ i_7_)  &  i_8_  &  n_n96  &  n_n85 ) ;
 assign wire389 = ( n_n99  &  n_n103  &  n_n63 ) ;
 assign wire390 = ( i_7_  &  i_8_  &  n_n103  &  n_n71 ) ;
 assign wire391 = ( n_n90  &  n_n102  &  n_n63 ) ;
 assign wire392 = ( n_n101  &  n_n100  &  n_n102 ) ;
 assign wire393 = ( n_n81  &  n_n82  &  n_n94 ) ;
 assign wire394 = ( n_n91  &  n_n92  &  n_n83 ) ;
 assign wire395 = ( n_n81  &  n_n93  &  n_n85 ) ;
 assign wire5943 = ( (~ i_5_)  &  (~ i_4_)  &  i_2_  &  i_0_ ) ;
 assign wire413 = ( i_7_  &  i_8_  &  (~ i_6_)  &  wire5943 ) ;
 assign wire430 = ( i_7_  &  i_8_  &  n_n79  &  n_n53 ) ;
 assign wire431 = ( i_7_  &  i_8_  &  n_n87  &  wire174 ) ;
 assign wire432 = ( i_7_  &  i_8_  &  n_n54  &  wire174 ) ;
 assign wire433 = ( n_n93  &  n_n103  &  n_n74 ) ;
 assign wire434 = ( n_n100  &  n_n92  &  n_n95 ) ;
 assign wire435 = ( (~ i_7_)  &  i_8_  &  n_n81  &  n_n103 ) ;
 assign wire436 = ( i_7_  &  i_6_  &  n_n103  &  n_n84 ) ;
 assign wire437 = ( n_n101  &  n_n99  &  n_n83 ) ;
 assign wire438 = ( n_n93  &  n_n92  &  n_n85 ) ;
 assign wire439 = ( n_n58  &  n_n103  &  n_n77 ) ;
 assign wire467 = ( (~ i_7_)  &  i_8_  &  n_n100  &  n_n40 ) ;
 assign wire468 = ( n_n81  &  n_n101  &  n_n85 ) ;
 assign wire469 = ( i_7_  &  i_6_  &  n_n99  &  n_n85 ) ;
 assign wire5847 = ( i_5_  &  i_6_  &  i_3_ ) ;
 assign wire475 = ( i_7_  &  i_8_  &  n_n90  &  wire5847 ) ;
 assign wire476 = ( (~ i_7_)  &  (~ i_8_)  &  n_n103  &  n_n76 ) ;
 assign wire477 = ( i_7_  &  i_8_  &  n_n85  &  n_n76 ) ;
 assign wire478 = ( n_n91  &  n_n100  &  n_n96 ) ;
 assign wire479 = ( n_n100  &  wire192  &  n_n102 ) ;
 assign wire480 = ( n_n92  &  n_n82  &  n_n90 ) ;
 assign wire481 = ( n_n100  &  n_n92  &  n_n63 ) ;
 assign wire482 = ( n_n91  &  n_n102  &  n_n94 ) ;
 assign wire483 = ( n_n91  &  n_n100  &  n_n77 ) ;
 assign wire484 = ( i_7_  &  i_6_  &  n_n103  &  n_n84 ) ;
 assign wire485 = ( n_n99  &  n_n82  &  n_n83 ) ;
 assign wire5828 = ( i_7_  &  (~ i_8_)  &  i_0_ ) ;
 assign wire507 = ( n_n74  &  (~ n_n67)  &  wire5828 ) ;
 assign wire508 = ( (~ i_7_)  &  i_8_  &  n_n103  &  n_n96 ) ;
 assign wire526 = ( (~ i_1_)  &  i_0_  &  n_n58  &  n_n54 ) ;
 assign wire532 = ( (~ i_5_)  &  (~ i_4_)  &  i_1_  &  _6377 ) ;
 assign wire5783 = ( i_7_  &  (~ i_6_)  &  (~ i_3_)  &  (~ i_4_) ) ;
 assign wire559 = ( i_1_  &  i_2_  &  (~ i_0_)  &  wire5783 ) ;
 assign wire562 = ( i_7_  &  (~ i_8_)  &  n_n84  &  n_n94 ) ;
 assign wire596 = ( (~ i_1_)  &  i_2_  &  i_0_  &  _6319 ) ;
 assign wire611 = ( i_7_  &  i_6_  &  n_n96  &  n_n83 ) ;
 assign wire5734 = ( (~ i_7_)  &  i_5_  &  (~ i_6_) ) ;
 assign wire5709 = ( (~ i_4_)  &  (~ i_1_)  &  i_0_ ) ;
 assign wire617 = ( n_n93  &  (~ n_n67)  &  wire5709 ) ;
 assign wire618 = ( i_7_  &  (~ i_8_)  &  n_n85  &  n_n40 ) ;
 assign wire619 = ( n_n74  &  n_n63  &  n_n85 ) ;
 assign wire620 = ( n_n93  &  n_n100  &  n_n74 ) ;
 assign wire621 = ( n_n81  &  n_n82  &  n_n94 ) ;
 assign wire5688 = ( i_5_  &  (~ i_6_)  &  (~ i_3_) ) ;
 assign wire641 = ( i_7_  &  i_8_  &  n_n97  &  wire5688 ) ;
 assign wire642 = ( (~ i_7_)  &  i_8_  &  n_n94  &  wire130 ) ;
 assign wire643 = ( i_7_  &  i_8_  &  n_n54  &  wire174 ) ;
 assign wire644 = ( i_7_  &  i_8_  &  n_n103  &  wire131 ) ;
 assign wire645 = ( n_n81  &  n_n101  &  n_n85 ) ;
 assign wire646 = ( n_n81  &  n_n91  &  n_n100 ) ;
 assign wire647 = ( n_n101  &  n_n84  &  n_n97 ) ;
 assign wire648 = ( n_n91  &  n_n99  &  n_n83 ) ;
 assign wire649 = ( n_n93  &  n_n74  &  n_n85 ) ;
 assign wire662 = ( n_n78  &  n_n92  &  n_n85 ) ;
 assign wire663 = ( n_n101  &  n_n103  &  n_n77 ) ;
 assign wire664 = ( i_7_  &  (~ i_8_)  &  n_n54  &  n_n53 ) ;
 assign wire5661 = ( i_7_  &  i_5_  &  (~ i_6_)  &  (~ i_3_) ) ;
 assign wire666 = ( i_1_  &  (~ i_2_)  &  (~ i_0_)  &  wire5661 ) ;
 assign wire668 = ( n_n93  &  n_n92  &  n_n83 ) ;
 assign wire669 = ( i_7_  &  i_8_  &  n_n103  &  n_n71 ) ;
 assign wire670 = ( n_n101  &  n_n99  &  n_n97 ) ;
 assign wire671 = ( n_n58  &  n_n90  &  n_n77 ) ;
 assign wire690 = ( n_n78  &  n_n103  &  n_n102 ) ;
 assign wire692 = ( (~ i_6_)  &  (~ i_3_)  &  wire172  &  n_n85 ) ;
 assign wire693 = ( n_n97  &  n_n92  &  n_n63 ) ;
 assign wire696 = ( i_7_  &  i_8_  &  n_n94  &  n_n66 ) ;
 assign wire5626 = ( (~ i_7_)  &  i_8_  &  i_6_  &  i_1_ ) ;
 assign wire697 = ( i_5_  &  (~ i_3_)  &  i_4_  &  wire5626 ) ;
 assign wire732 = ( (~ i_7_)  &  i_8_  &  n_n87  &  n_n67 ) ;
 assign wire734 = ( i_7_  &  (~ i_8_)  &  n_n97  &  wire127 ) ;
 assign wire736 = ( n_n78  &  n_n97  &  n_n102 ) ;
 assign wire755 = ( (~ i_7_)  &  i_8_  &  n_n94  &  wire130 ) ;
 assign wire756 = ( (~ i_7_)  &  (~ i_8_)  &  n_n103  &  wire130 ) ;
 assign wire757 = ( i_7_  &  (~ i_8_)  &  n_n71  &  wire242 ) ;
 assign wire758 = ( n_n100  &  n_n102  &  n_n63 ) ;
 assign wire759 = ( (~ i_7_)  &  (~ i_8_)  &  n_n99  &  n_n83 ) ;
 assign wire805 = ( n_n97  &  n_n82  &  n_n102 ) ;
 assign wire5558 = ( (~ i_3_)  &  i_4_  &  i_1_  &  i_0_ ) ;
 assign wire807 = ( (~ i_7_)  &  i_8_  &  i_6_  &  wire5558 ) ;
 assign wire808 = ( (~ i_7_)  &  i_8_  &  n_n87  &  n_n67 ) ;
 assign wire812 = ( (~ i_7_)  &  i_8_  &  n_n71  &  n_n67 ) ;
 assign wire5544 = ( i_7_  &  (~ i_8_)  &  i_6_  &  (~ i_3_) ) ;
 assign wire825 = ( (~ i_1_)  &  i_2_  &  i_0_  &  wire5544 ) ;
 assign wire827 = ( (~ i_7_)  &  (~ i_8_)  &  n_n54  &  n_n83 ) ;
 assign wire833 = ( i_7_  &  i_8_  &  n_n87  &  wire174 ) ;
 assign wire834 = ( (~ i_7_)  &  i_8_  &  n_n96  &  n_n85 ) ;
 assign wire835 = ( n_n81  &  n_n95  &  n_n94 ) ;
 assign wire836 = ( n_n101  &  n_n92  &  n_n90 ) ;
 assign wire839 = ( n_n100  &  n_n102  &  n_n63 ) ;
 assign wire840 = ( n_n58  &  n_n100  &  n_n77 ) ;
 assign wire864 = ( n_n81  &  n_n78  &  n_n97 ) ;
 assign wire866 = ( i_7_  &  (~ i_8_)  &  n_n81  &  n_n100 ) ;
 assign wire867 = ( n_n93  &  n_n74  &  n_n85 ) ;
 assign wire870 = ( n_n82  &  n_n83  &  n_n77 ) ;
 assign wire871 = ( n_n95  &  n_n90  &  n_n77 ) ;
 assign wire872 = ( (~ i_8_)  &  i_6_  &  n_n74  &  n_n83 ) ;
 assign wire873 = ( n_n58  &  n_n84  &  n_n97 ) ;
 assign wire874 = ( i_7_  &  i_8_  &  n_n54  &  wire322 ) ;
 assign wire876 = ( n_n81  &  n_n93  &  n_n103 ) ;
 assign wire877 = ( n_n99  &  n_n82  &  n_n83 ) ;
 assign wire5498 = ( (~ i_5_)  &  (~ i_4_)  &  i_1_  &  (~ i_0_) ) ;
 assign wire878 = ( i_7_  &  (~ i_8_)  &  (~ i_6_)  &  wire5498 ) ;
 assign wire895 = ( (~ i_7_)  &  (~ i_8_)  &  n_n97  &  n_n77 ) ;
 assign wire897 = ( n_n91  &  n_n84  &  n_n85 ) ;
 assign wire899 = ( i_5_  &  i_3_  &  n_n93  &  n_n97 ) ;
 assign wire900 = ( i_7_  &  i_8_  &  n_n94  &  n_n66 ) ;
 assign wire901 = ( n_n74  &  n_n63  &  n_n85 ) ;
 assign wire5457 = ( i_7_  &  i_3_  &  i_1_  &  (~ i_2_) ) ;
 assign wire906 = ( (~ i_5_)  &  (~ i_6_)  &  i_4_  &  wire5457 ) ;
 assign wire5458 = ( i_8_  &  i_3_  &  (~ i_2_)  &  i_0_ ) ;
 assign wire907 = ( i_5_  &  (~ i_6_)  &  (~ i_4_)  &  wire5458 ) ;
 assign wire5459 = ( i_8_  &  i_6_  &  (~ i_3_)  &  i_4_ ) ;
 assign wire908 = ( i_1_  &  (~ i_2_)  &  i_0_  &  wire5459 ) ;
 assign wire909 = ( (~ i_7_)  &  i_6_  &  n_n99  &  n_n83 ) ;
 assign wire910 = ( i_7_  &  i_8_  &  n_n103  &  n_n40 ) ;
 assign wire911 = ( n_n91  &  n_n84  &  n_n85 ) ;
 assign wire940 = ( (~ i_7_)  &  i_8_  &  n_n71  &  n_n67 ) ;
 assign wire942 = ( (~ i_7_)  &  (~ i_6_)  &  n_n103  &  n_n92 ) ;
 assign wire944 = ( n_n97  &  n_n96  &  n_n63 ) ;
 assign wire946 = ( i_7_  &  (~ i_8_)  &  n_n79  &  n_n53 ) ;
 assign wire948 = ( i_7_  &  i_8_  &  n_n40  &  n_n53 ) ;
 assign wire5444 = ( (~ i_7_)  &  i_8_  &  (~ i_5_)  &  i_6_ ) ;
 assign wire950 = ( (~ i_1_)  &  i_2_  &  (~ i_0_)  &  wire5444 ) ;
 assign wire957 = ( n_n82  &  n_n102  &  n_n83 ) ;
 assign wire958 = ( n_n84  &  n_n63  &  n_n85 ) ;
 assign wire959 = ( i_7_  &  (~ i_8_)  &  n_n87  &  wire353 ) ;
 assign wire960 = ( n_n83  &  n_n63  &  wire194 ) ;
 assign wire961 = ( n_n58  &  n_n84  &  n_n97 ) ;
 assign wire962 = ( n_n81  &  n_n78  &  n_n97 ) ;
 assign wire963 = ( n_n101  &  n_n103  &  n_n84 ) ;
 assign wire5423 = ( i_5_  &  (~ i_6_)  &  (~ i_3_) ) ;
 assign wire978 = ( (~ i_7_)  &  (~ i_8_)  &  n_n83  &  wire5423 ) ;
 assign wire979 = ( n_n91  &  n_n84  &  n_n94 ) ;
 assign wire980 = ( (~ i_8_)  &  (~ i_6_)  &  n_n100  &  n_n92 ) ;
 assign wire981 = ( i_7_  &  i_8_  &  n_n99  &  n_n90 ) ;
 assign wire982 = ( i_7_  &  i_8_  &  n_n71  &  wire242 ) ;
 assign wire983 = ( n_n58  &  n_n100  &  n_n84 ) ;
 assign wire984 = ( n_n99  &  n_n97  &  n_n95 ) ;
 assign wire985 = ( n_n78  &  n_n92  &  n_n85 ) ;
 assign wire986 = ( n_n92  &  n_n82  &  n_n94 ) ;
 assign wire989 = ( n_n93  &  n_n100  &  n_n84 ) ;
 assign wire1009 = ( i_7_  &  i_8_  &  n_n100  &  wire131 ) ;
 assign wire1011 = ( n_n91  &  n_n102  &  n_n83 ) ;
 assign wire1012 = ( n_n58  &  n_n103  &  n_n92 ) ;
 assign wire5398 = ( (~ i_8_)  &  i_6_  &  i_3_  &  (~ i_4_) ) ;
 assign wire1013 = ( i_1_  &  i_2_  &  i_0_  &  wire5398 ) ;
 assign wire1024 = ( i_7_  &  i_8_  &  n_n74  &  n_n85 ) ;
 assign wire1039 = ( i_7_  &  (~ i_8_)  &  n_n66  &  n_n67 ) ;
 assign wire5375 = ( i_7_  &  (~ i_3_)  &  i_1_  &  i_2_ ) ;
 assign wire1041 = ( i_5_  &  (~ i_6_)  &  (~ i_4_)  &  wire5375 ) ;
 assign wire1043 = ( i_7_  &  (~ i_8_)  &  n_n84  &  n_n97 ) ;
 assign wire1046 = ( i_7_  &  (~ i_8_)  &  n_n79  &  n_n53 ) ;
 assign wire1048 = ( n_n97  &  n_n96  &  n_n63 ) ;
 assign wire1080 = ( i_7_  &  (~ i_8_)  &  n_n84  &  n_n94 ) ;
 assign wire1082 = ( (~ i_8_)  &  (~ i_6_)  &  n_n96  &  n_n94 ) ;
 assign wire5319 = ( (~ i_8_)  &  (~ i_6_)  &  (~ i_3_) ) ;
 assign wire1085 = ( i_7_  &  i_6_  &  n_n96  &  n_n83 ) ;
 assign wire5318 = ( i_8_  &  i_3_  &  (~ i_1_)  &  i_0_ ) ;
 assign wire5276 = ( i_5_  &  i_4_  &  (~ i_1_)  &  i_2_ ) ;
 assign wire1106 = ( i_7_  &  i_8_  &  i_6_  &  wire5276 ) ;
 assign wire5277 = ( i_7_  &  i_8_  &  i_1_ ) ;
 assign wire1107 = ( i_3_  &  i_2_  &  n_n40  &  wire5277 ) ;
 assign wire5279 = ( i_5_  &  i_6_  &  i_3_ ) ;
 assign wire1108 = ( i_7_  &  i_8_  &  n_n90  &  wire5279 ) ;
 assign wire1109 = ( _5644  &  _5645 ) ;
 assign wire5281 = ( (~ i_7_)  &  i_8_  &  i_4_ ) ;
 assign wire1110 = ( (~ i_6_)  &  i_3_  &  n_n100  &  wire5281 ) ;
 assign wire1111 = ( i_1_  &  (~ i_0_)  &  n_n93  &  n_n102 ) ;
 assign wire1112 = ( i_7_  &  i_8_  &  n_n97  &  wire127 ) ;
 assign wire1113 = ( (~ i_7_)  &  (~ i_8_)  &  n_n103  &  n_n76 ) ;
 assign wire1114 = ( i_7_  &  i_8_  &  n_n100  &  n_n76 ) ;
 assign wire1115 = ( i_7_  &  (~ i_8_)  &  n_n71  &  wire242 ) ;
 assign wire1116 = ( i_7_  &  i_8_  &  n_n103  &  wire131 ) ;
 assign wire1117 = ( n_n93  &  n_n84  &  n_n90 ) ;
 assign wire1118 = ( (~ i_3_)  &  (~ i_1_)  &  i_0_  &  _5668 ) ;
 assign wire1119 = ( n_n91  &  n_n84  &  n_n94 ) ;
 assign wire1120 = ( n_n82  &  n_n102  &  n_n83 ) ;
 assign wire1123 = ( n_n93  &  n_n77  &  n_n85 ) ;
 assign wire1142 = ( n_n101  &  n_n96  &  n_n94 ) ;
 assign wire1143 = ( n_n58  &  n_n100  &  n_n84 ) ;
 assign wire1144 = ( n_n101  &  n_n77  &  n_n85 ) ;
 assign wire1145 = ( n_n103  &  n_n82  &  n_n77 ) ;
 assign wire1155 = ( i_8_  &  (~ i_6_)  &  n_n74  &  n_n90 ) ;
 assign wire1156 = ( n_n81  &  n_n83  &  n_n63 ) ;
 assign wire1293 = ( i_7_  &  (~ i_3_)  &  (~ i_4_)  &  (~ i_0_) ) ;
 assign wire1294 = ( (~ i_5_)  &  (~ i_3_)  &  (~ i_4_)  &  (~ i_0_) ) ;
 assign wire5251 = ( (~ i_7_)  &  (~ i_8_)  &  (~ i_1_) ) ;
 assign wire1157 = ( wire1293  &  wire5251 ) | ( wire1294  &  wire5251 ) ;
 assign wire1173 = ( n_n58  &  n_n102  &  n_n94 ) ;
 assign wire1175 = ( i_7_  &  (~ i_6_)  &  n_n74  &  n_n90 ) ;
 assign wire1177 = ( n_n92  &  n_n82  &  n_n90 ) ;
 assign wire1179 = ( i_7_  &  (~ i_6_)  &  n_n74  &  n_n90 ) ;
 assign wire1191 = ( n_n95  &  n_n90  &  n_n77 ) ;
 assign wire1192 = ( n_n81  &  n_n93  &  n_n94 ) ;
 assign wire1193 = ( (~ i_7_)  &  (~ i_8_)  &  wire241  &  n_n40 ) ;
 assign wire1194 = ( n_n91  &  n_n92  &  n_n90 ) ;
 assign wire1197 = ( n_n93  &  n_n100  &  n_n102 ) ;
 assign wire1213 = ( (~ i_7_)  &  (~ i_8_)  &  n_n83  &  n_n79 ) ;
 assign wire1214 = ( n_n91  &  n_n99  &  n_n85 ) ;
 assign wire1215 = ( i_7_  &  i_8_  &  n_n54  &  n_n85 ) ;
 assign wire1234 = ( n_n83  &  n_n63  &  wire194 ) ;
 assign wire1235 = ( i_7_  &  (~ i_6_)  &  n_n103  &  n_n102 ) ;
 assign wire5143 = ( (~ i_7_)  &  (~ i_8_)  &  (~ i_1_) ) ;
 assign wire1253 = ( wire1293  &  wire5143 ) | ( wire1294  &  wire5143 ) ;
 assign wire1254 = ( i_7_  &  i_8_  &  n_n85  &  n_n76 ) ;
 assign wire1255 = ( n_n101  &  n_n92  &  n_n90 ) ;
 assign wire1256 = ( n_n84  &  n_n83  &  n_n63 ) ;
 assign wire1257 = ( n_n93  &  n_n90  &  n_n77 ) ;
 assign wire1281 = ( i_7_  &  i_6_  &  n_n99  &  n_n85 ) ;
 assign wire1283 = ( n_n58  &  n_n99  &  n_n94 ) ;
 assign wire1285 = ( n_n78  &  n_n97  &  n_n74 ) ;
 assign wire1286 = ( n_n93  &  n_n77  &  n_n94 ) ;
 assign wire1287 = ( n_n93  &  n_n84  &  n_n90 ) ;
 assign wire1288 = ( n_n99  &  n_n103  &  n_n63 ) ;
 assign wire5141 = ( (~ i_3_)  &  i_2_  &  i_0_ ) ;
 assign wire1289 = ( i_7_  &  i_8_  &  n_n54  &  wire5141 ) ;
 assign wire1290 = ( n_n93  &  n_n103  &  n_n77 ) ;
 assign wire1291 = ( n_n101  &  n_n103  &  n_n84 ) ;
 assign wire1292 = ( n_n93  &  n_n92  &  n_n85 ) ;
 assign wire1295 = ( i_8_  &  (~ i_6_)  &  n_n81  &  n_n85 ) ;
 assign wire1313 = ( i_7_  &  i_6_  &  n_n102  &  n_n94 ) ;
 assign wire1317 = ( n_n92  &  n_n90  &  wire177 ) ;
 assign wire1318 = ( (~ i_7_)  &  i_6_  &  n_n99  &  n_n83 ) ;
 assign wire1319 = ( n_n92  &  n_n82  &  n_n85 ) ;
 assign wire1320 = ( i_7_  &  i_6_  &  n_n102  &  n_n94 ) ;
 assign wire1350 = ( n_n58  &  n_n103  &  n_n77 ) | ( n_n58  &  n_n90  &  n_n77 ) ;
 assign wire1351 = ( n_n91  &  n_n103  &  n_n77 ) ;
 assign wire1352 = ( n_n100  &  n_n84  &  n_n95 ) ;
 assign wire1354 = ( i_7_  &  (~ i_6_)  &  n_n103  &  n_n84 ) ;
 assign wire1356 = ( (~ i_7_)  &  (~ i_8_)  &  n_n66  &  wire353 ) ;
 assign wire1357 = ( n_n93  &  n_n77  &  n_n85 ) ;
 assign wire1358 = ( n_n101  &  n_n102  &  n_n83 ) ;
 assign wire1359 = ( n_n74  &  n_n82  &  n_n94 ) ;
 assign wire1360 = ( (~ i_7_)  &  (~ i_8_)  &  n_n83  &  wire354 ) ;
 assign wire1361 = ( n_n93  &  n_n103  &  n_n77 ) | ( n_n93  &  n_n90  &  n_n77 ) ;
 assign wire1362 = ( n_n99  &  n_n82  &  n_n85 ) ;
 assign wire1380 = ( n_n91  &  n_n99  &  n_n85 ) ;
 assign wire1381 = ( n_n91  &  n_n83  &  n_n77 ) ;
 assign wire1382 = ( i_7_  &  i_8_  &  n_n85  &  n_n87 ) ;
 assign wire1383 = ( n_n101  &  n_n84  &  n_n97 ) ;
 assign wire1388 = ( n_n99  &  n_n63  &  n_n85 ) ;
 assign wire1389 = ( (~ i_7_)  &  (~ i_8_)  &  n_n99  &  n_n83 ) ;
 assign wire1411 = ( n_n83  &  n_n63  &  n_n77 ) ;
 assign wire1413 = ( n_n103  &  n_n92  &  n_n82 ) ;
 assign wire1414 = ( n_n81  &  n_n97  &  n_n63 ) ;
 assign wire1415 = ( n_n91  &  n_n83  &  n_n77 ) ;
 assign wire1417 = ( n_n93  &  n_n97  &  n_n74 ) ;
 assign wire1421 = ( (~ i_7_)  &  (~ i_6_)  &  n_n99  &  n_n83 ) ;
 assign wire1440 = ( n_n93  &  n_n84  &  n_n94 ) ;
 assign wire1443 = ( i_1_  &  i_2_  &  n_n58  &  n_n102 ) ;
 assign wire4958 = ( (~ i_7_)  &  (~ i_8_)  &  i_1_  &  i_0_ ) ;
 assign wire1445 = ( i_5_  &  i_3_  &  i_4_  &  wire4958 ) ;
 assign wire4959 = ( (~ i_7_)  &  (~ i_8_)  &  i_5_  &  (~ i_6_) ) ;
 assign wire1446 = ( (~ i_1_)  &  (~ i_2_)  &  i_0_  &  wire4959 ) ;
 assign wire1447 = ( i_7_  &  i_8_  &  n_n97  &  wire127 ) ;
 assign wire1448 = ( n_n74  &  n_n82  &  n_n94 ) ;
 assign wire1449 = ( n_n97  &  n_n82  &  n_n102 ) ;
 assign wire1450 = ( n_n100  &  n_n84  &  n_n82 ) ;
 assign wire1451 = ( (~ i_7_)  &  (~ i_6_)  &  n_n103  &  n_n92 ) ;
 assign wire1452 = ( n_n103  &  n_n82  &  n_n77 ) ;
 assign wire4952 = ( (~ i_7_)  &  (~ i_8_)  &  i_6_  &  (~ i_4_) ) ;
 assign wire1483 = ( (~ i_7_)  &  i_8_  &  n_n103  &  n_n96 ) ;
 assign wire1484 = ( i_7_  &  (~ i_8_)  &  n_n102  &  n_n85 ) ;
 assign wire1485 = ( i_7_  &  (~ i_6_)  &  n_n84  &  n_n90 ) ;
 assign wire1486 = ( (~ i_7_)  &  i_8_  &  n_n96  &  n_n94 ) ;
 assign wire1487 = ( (~ i_7_)  &  (~ i_6_)  &  n_n99  &  n_n83 ) ;
 assign wire1489 = ( n_n81  &  n_n91  &  n_n100 ) ;
 assign wire1490 = ( n_n91  &  n_n74  &  n_n83 ) ;
 assign wire1491 = ( n_n84  &  n_n63  &  n_n85 ) ;
 assign wire1499 = ( i_7_  &  i_8_  &  n_n84  &  n_n83 ) ;
 assign wire1507 = ( i_5_  &  (~ i_3_)  &  n_n93  &  n_n85 ) ;
 assign wire1508 = ( (~ i_7_)  &  i_8_  &  n_n83  &  n_n66 ) ;
 assign wire4931 = ( (~ i_7_)  &  i_8_  &  i_4_ ) ;
 assign wire1509 = ( (~ i_6_)  &  i_3_  &  n_n100  &  wire4931 ) ;
 assign wire1510 = ( i_1_  &  (~ i_0_)  &  n_n93  &  n_n102 ) ;
 assign wire1511 = ( (~ i_7_)  &  (~ i_8_)  &  n_n83  &  wire354 ) ;
 assign wire4930 = ( (~ i_3_)  &  i_1_  &  i_0_ ) ;
 assign wire1520 = ( i_8_  &  (~ i_6_)  &  n_n100  &  n_n102 ) ;
 assign wire1521 = ( n_n91  &  n_n92  &  n_n90 ) ;
 assign wire1522 = ( n_n100  &  n_n84  &  n_n63 ) ;
 assign wire1523 = ( n_n103  &  n_n92  &  n_n82 ) ;
 assign wire1524 = ( n_n81  &  n_n78  &  n_n103 ) ;
 assign wire1525 = ( n_n101  &  n_n99  &  n_n83 ) ;
 assign wire1527 = ( n_n92  &  n_n82  &  n_n94 ) ;
 assign wire4921 = ( i_3_  &  i_1_  &  i_2_ ) ;
 assign wire1533 = ( (~ i_7_)  &  i_8_  &  n_n79  &  wire4921 ) ;
 assign wire1534 = ( n_n78  &  n_n103  &  n_n102 ) ;
 assign wire1535 = ( n_n97  &  n_n102  &  n_n63 ) ;
 assign wire1536 = ( n_n81  &  n_n91  &  n_n97 ) ;
 assign wire1559 = ( n_n91  &  n_n71  &  n_n67 ) ;
 assign wire1560 = ( (~ i_5_)  &  (~ i_6_)  &  (~ i_4_)  &  _4857 ) ;
 assign wire1562 = ( i_7_  &  (~ i_6_)  &  n_n103  &  n_n84 ) ;
 assign wire1583 = ( (~ i_1_)  &  i_2_  &  i_0_  &  _4881 ) ;
 assign wire4841 = ( (~ i_7_)  &  i_8_  &  (~ i_1_)  &  i_2_ ) ;
 assign wire1589 = ( n_n81  &  (~ wire192)  &  wire4841 ) ;
 assign wire1590 = ( (~ i_7_)  &  i_8_  &  n_n80  &  n_n54 ) ;
 assign wire1591 = ( (~ i_6_)  &  i_3_  &  n_n100  &  wire172 ) ;
 assign wire1592 = ( i_7_  &  i_6_  &  n_n81  &  n_n85 ) ;
 assign wire1595 = ( i_7_  &  i_6_  &  n_n81  &  n_n83 ) ;
 assign wire1596 = ( n_n93  &  n_n100  &  n_n74 ) ;
 assign wire1599 = ( n_n101  &  n_n96  &  n_n94 ) ;
 assign wire1600 = ( n_n78  &  n_n97  &  n_n74 ) ;
 assign wire1601 = ( n_n58  &  n_n102  &  n_n94 ) ;
 assign wire1602 = ( n_n58  &  n_n103  &  n_n92 ) ;
 assign wire1617 = ( n_n91  &  n_n99  &  n_n97 ) ;
 assign wire1618 = ( n_n101  &  n_n97  &  n_n96 ) ;
 assign wire1619 = ( n_n103  &  n_n74  &  n_n95 ) ;
 assign wire1620 = ( n_n81  &  n_n93  &  n_n94 ) ;
 assign wire1621 = ( n_n99  &  n_n63  &  n_n85 ) ;
 assign wire1622 = ( n_n100  &  n_n84  &  n_n95 ) ;
 assign wire1623 = ( n_n93  &  n_n92  &  n_n83 ) ;
 assign wire1624 = ( n_n99  &  n_n97  &  n_n95 ) ;
 assign wire4840 = ( i_3_  &  (~ i_1_)  &  i_0_ ) ;
 assign wire1625 = ( (~ i_7_)  &  (~ i_8_)  &  n_n40  &  wire4840 ) ;
 assign wire1627 = ( n_n100  &  n_n92  &  n_n95 ) ;
 assign wire1628 = ( n_n91  &  n_n100  &  n_n77 ) ;
 assign wire1629 = ( (~ i_7_)  &  (~ i_6_)  &  n_n97  &  n_n77 ) ;
 assign wire1631 = ( i_7_  &  (~ i_8_)  &  n_n100  &  n_n54 ) ;
 assign wire4849 = ( n_n100  &  n_n84  &  wire192 ) | ( n_n100  &  wire192  &  n_n92 ) ;
 assign wire4851 = ( n_n101  &  n_n102  &  n_n83 ) | ( n_n91  &  n_n102  &  n_n83 ) ;
 assign wire4854 = ( n_n1217 ) | ( wire1627 ) | ( wire1628 ) | ( wire1629 ) ;
 assign wire4855 = ( wire357 ) | ( wire1623 ) | ( wire1624 ) | ( wire1625 ) ;
 assign wire4856 = ( wire1619 ) | ( wire1620 ) | ( wire1621 ) | ( wire1622 ) ;
 assign wire4857 = ( n_n1281 ) | ( n_n1185 ) | ( wire1617 ) | ( wire1618 ) ;
 assign wire4858 = ( n_n1174 ) | ( wire235 ) | ( wire252 ) | ( wire329 ) ;
 assign wire4859 = ( wire1589 ) | ( wire1590 ) | ( wire1591 ) | ( wire1592 ) ;
 assign wire4861 = ( wire1599 ) | ( wire1600 ) | ( wire4851 ) ;
 assign wire4875 = ( i_3_  &  i_1_  &  i_0_ ) ;
 assign wire4876 = ( i_7_  &  (~ i_8_)  &  (~ i_6_)  &  (~ i_4_) ) ;
 assign wire4877 = ( i_7_  &  (~ i_6_)  &  (~ i_3_)  &  i_4_ ) ;
 assign wire4878 = ( wire4875  &  wire4876 ) | ( n_n85  &  wire4877 ) ;
 assign wire4887 = ( n_n99  &  n_n95  &  n_n85 ) | ( n_n96  &  n_n95  &  n_n85 ) ;
 assign wire4890 = ( n_n1036 ) | ( n_n1035 ) | ( _4865 ) ;
 assign wire4891 = ( n_n1046 ) | ( n_n1026 ) | ( wire1583 ) | ( wire4878 ) ;
 assign wire4892 = ( n_n1022 ) | ( n_n1052 ) | ( (~ i_8_)  &  wire70 ) ;
 assign wire4893 = ( n_n1042 ) | ( n_n1043 ) | ( n_n1059 ) | ( n_n1048 ) ;
 assign wire4894 = ( n_n1009 ) | ( n_n1011 ) | ( n_n1025 ) | ( n_n1013 ) ;
 assign wire4895 = ( wire249 ) | ( wire1559 ) | ( wire4887 ) ;
 assign wire4899 = ( wire1560 ) | ( wire1562 ) | ( wire4890 ) | ( wire4895 ) ;
 assign wire4900 = ( wire4891 ) | ( wire4892 ) | ( wire4893 ) | ( wire4894 ) ;
 assign wire4904 = ( i_7_  &  i_3_  &  i_0_ ) | ( i_7_  &  i_2_  &  i_0_ ) ;
 assign wire4910 = ( n_n943 ) | ( n_n77  &  wire4904 ) ;
 assign wire4911 = ( n_n989 ) | ( n_n951 ) | ( n_n950 ) | ( n_n991 ) ;
 assign wire4912 = ( n_n982 ) | ( n_n967 ) | ( wire203 ) ;
 assign wire4913 = ( n_n961 ) | ( n_n952 ) | ( n_n986 ) | ( n_n976 ) ;
 assign wire4914 = ( n_n940 ) | ( n_n1006 ) | ( n_n984 ) | ( n_n978 ) ;
 assign wire4919 = ( wire298 ) | ( wire292 ) | ( n_n882 ) | ( wire4910 ) ;
 assign wire4920 = ( wire4911 ) | ( wire4912 ) | ( wire4913 ) | ( wire4914 ) ;
 assign wire4928 = ( n_n1330 ) | ( wire1520 ) | ( wire1521 ) | ( wire1527 ) ;
 assign wire4929 = ( wire1522 ) | ( wire1523 ) | ( wire1524 ) | ( wire1525 ) ;
 assign wire4954 = ( i_7_  &  i_6_  &  i_1_ ) ;
 assign wire4955 = ( i_8_  &  i_5_  &  i_3_  &  i_0_ ) ;
 assign wire4957 = ( (~ i_7_)  &  (~ i_8_)  &  i_5_  &  (~ i_4_) ) ;
 assign wire4960 = ( wire4954  &  wire4955 ) | ( n_n80  &  wire4957 ) ;
 assign wire4971 = ( wire1489 ) | ( wire1490 ) | ( wire4960 ) ;
 assign wire4972 = ( n_n1082 ) | ( wire1485 ) | ( wire1486 ) | ( wire1487 ) ;
 assign wire4973 = ( n_n1079 ) | ( n_n1070 ) | ( wire1483 ) | ( wire1484 ) ;
 assign wire4974 = ( n_n1077 ) | ( n_n1172 ) | ( n_n1078 ) | ( wire1445 ) ;
 assign wire4975 = ( n_n1081 ) | ( n_n1279 ) | ( n_n1153 ) | ( n_n1297 ) ;
 assign wire4976 = ( n_n1324 ) | ( n_n1092 ) | ( wire251 ) | ( wire321 ) ;
 assign wire4977 = ( wire1443 ) | ( wire1446 ) | ( wire1447 ) | ( wire1448 ) ;
 assign wire4978 = ( wire1449 ) | ( wire1450 ) | ( wire1451 ) | ( wire1452 ) ;
 assign wire4983 = ( wire232 ) | ( wire4928 ) | ( wire4929 ) ;
 assign wire4984 = ( wire4971 ) | ( wire4972 ) | ( wire4973 ) | ( wire4974 ) ;
 assign wire4985 = ( wire4975 ) | ( wire4976 ) | ( wire4977 ) | ( wire4978 ) ;
 assign wire4997 = ( n_n91  &  n_n103  &  n_n74 ) | ( n_n103  &  n_n74  &  n_n63 ) ;
 assign wire5001 = ( n_n1055 ) | ( n_n1085 ) | ( wire1421 ) ;
 assign wire5002 = ( n_n1158 ) | ( n_n1146 ) | ( n_n1163 ) | ( n_n1160 ) ;
 assign wire5003 = ( n_n1134 ) | ( n_n1132 ) | ( wire335 ) | ( wire1440 ) ;
 assign wire5004 = ( n_n1172 ) | ( n_n1022 ) | ( n_n1093 ) | ( n_n1128 ) ;
 assign wire5005 = ( n_n1164 ) | ( n_n1130 ) | ( wire4997 ) ;
 assign wire5006 = ( n_n1181 ) | ( wire356 ) | ( _5183 ) ;
 assign wire5010 = ( wire299 ) | ( wire5001 ) | ( wire5006 ) ;
 assign wire5011 = ( wire5002 ) | ( wire5003 ) | ( wire5004 ) | ( wire5005 ) ;
 assign wire5015 = ( n_n93  &  n_n100  &  n_n77 ) | ( n_n93  &  n_n83  &  n_n77 ) ;
 assign wire5020 = ( n_n951 ) | ( n_n950 ) | ( wire135 ) ;
 assign wire5021 = ( n_n942 ) | ( n_n973 ) | ( n_n938 ) | ( n_n975 ) ;
 assign wire5022 = ( n_n956 ) | ( n_n1014 ) | ( n_n1018 ) | ( n_n955 ) ;
 assign wire5023 = ( wire1557 ) | ( wire1558 ) | ( wire5015 ) ;
 assign wire5024 = ( n_n961 ) | ( n_n964 ) | ( n_n981 ) | ( n_n1004 ) ;
 assign wire5025 = ( n_n1021 ) | ( n_n991 ) | ( wire249 ) | ( n_n978 ) ;
 assign wire5029 = ( wire291 ) | ( wire5020 ) | ( wire5025 ) ;
 assign wire5030 = ( wire5021 ) | ( wire5022 ) | ( wire5023 ) | ( wire5024 ) ;
 assign wire5036 = ( n_n1217 ) | ( wire1535 ) | ( wire1536 ) | ( wire1629 ) ;
 assign wire5037 = ( n_n1281 ) | ( n_n1279 ) | ( n_n1188 ) | ( wire1417 ) ;
 assign wire5038 = ( wire346 ) | ( wire1413 ) | ( wire1414 ) | ( wire1415 ) ;
 assign wire5039 = ( n_n1185 ) | ( n_n1193 ) | ( wire343 ) | ( wire1411 ) ;
 assign wire5040 = ( n_n1254 ) | ( n_n1259 ) | ( n_n1204 ) | ( n_n1369 ) ;
 assign wire5041 = ( wire314 ) | ( wire349 ) | ( wire1388 ) | ( wire1389 ) ;
 assign wire5057 = ( n_n1217 ) | ( wire1535 ) | ( wire1536 ) | ( wire1629 ) ;
 assign wire5058 = ( wire1380 ) | ( wire1381 ) | ( wire1382 ) | ( wire1383 ) ;
 assign wire5059 = ( n_n1185 ) | ( n_n1172 ) | ( wire1361 ) ;
 assign wire5060 = ( n_n1153 ) | ( wire349 ) | ( n_n1267 ) | ( wire342 ) ;
 assign wire5061 = ( n_n1164 ) | ( n_n1184 ) | ( n_n1216 ) | ( n_n1146 ) ;
 assign wire5062 = ( n_n1170 ) | ( wire343 ) | ( wire1360 ) | ( wire1362 ) ;
 assign wire5072 = ( n_n978 ) | ( wire135 ) | ( n_n90  &  wire5012 ) ;
 assign wire5073 = ( n_n959 ) | ( n_n957 ) | ( n_n1001 ) | ( n_n1010 ) ;
 assign wire5074 = ( n_n971 ) | ( n_n976 ) | ( n_n1014 ) | ( n_n1018 ) ;
 assign wire5075 = ( n_n941 ) | ( n_n943 ) | ( n_n939 ) | ( n_n981 ) ;
 assign wire5076 = ( n_n983 ) | ( n_n940 ) | ( n_n999 ) | ( wire249 ) ;
 assign wire5080 = ( wire297 ) | ( wire305 ) | ( wire5076 ) ;
 assign wire5081 = ( wire5072 ) | ( wire5073 ) | ( wire5074 ) | ( wire5075 ) ;
 assign wire5093 = ( wire1320 ) | ( wire1358 ) | ( wire1359 ) ;
 assign wire5094 = ( n_n1058 ) | ( wire1354 ) | ( wire1356 ) | ( wire1357 ) ;
 assign wire5095 = ( wire323 ) | ( n_n1032 ) | ( n_n1040 ) | ( wire1352 ) ;
 assign wire5096 = ( n_n1036 ) | ( n_n1035 ) | ( n_n1055 ) | ( n_n1085 ) ;
 assign wire5097 = ( n_n1020 ) | ( n_n83  &  wire35 ) | ( n_n83  &  _4906 ) ;
 assign wire5098 = ( n_n1324 ) | ( n_n1092 ) | ( n_n1022 ) | ( n_n1134 ) ;
 assign wire5099 = ( n_n1039 ) | ( n_n1091 ) | ( n_n1093 ) | ( n_n1103 ) ;
 assign wire5100 = ( n_n1120 ) | ( n_n1052 ) | ( n_n1331 ) | ( wire1317 ) ;
 assign wire5101 = ( wire1318 ) | ( wire1319 ) | ( wire1350 ) | ( wire1351 ) ;
 assign wire5106 = ( wire5100 ) | ( wire5101 ) ;
 assign wire5107 = ( wire257 ) | ( wire5093 ) | ( wire5094 ) | ( wire5095 ) ;
 assign wire5117 = ( n_n944 ) | ( n_n939 ) | ( n_n1025 ) | ( n_n1020 ) ;
 assign wire5118 = ( n_n954 ) | ( n_n952 ) | ( n_n959 ) | ( n_n957 ) ;
 assign wire5119 = ( n_n971 ) | ( n_n1001 ) | ( n_n976 ) | ( n_n1010 ) ;
 assign wire5120 = ( wire189 ) | ( n_n958 ) | ( n_n989 ) | ( n_n1030 ) ;
 assign wire5121 = ( n_n961 ) | ( n_n949 ) | ( n_n969 ) | ( n_n966 ) ;
 assign wire5130 = ( _83 ) | ( n_n78  &  n_n103  &  n_n96 ) ;
 assign wire5131 = ( n_n1058 ) | ( wire1295 ) | ( wire1354 ) ;
 assign wire5132 = ( n_n1103 ) | ( n_n1095 ) | ( n_n1070 ) | ( wire1313 ) ;
 assign wire5133 = ( n_n1153 ) | ( n_n1092 ) | ( n_n1173 ) | ( n_n1170 ) ;
 assign wire5134 = ( n_n1120 ) | ( n_n1052 ) | ( n_n1082 ) | ( n_n1035 ) ;
 assign wire5139 = ( wire257 ) | ( wire306 ) | ( wire106 ) | ( wire5130 ) ;
 assign wire5140 = ( wire5131 ) | ( wire5132 ) | ( wire5133 ) | ( wire5134 ) ;
 assign wire5150 = ( wire357 ) | ( wire1621 ) | ( wire1622 ) | ( wire1625 ) ;
 assign wire5151 = ( wire1358 ) | ( wire1359 ) | ( wire1489 ) | ( wire1490 ) ;
 assign wire5152 = ( wire1291 ) | ( wire1292 ) | ( wire1356 ) | ( wire1357 ) ;
 assign wire5153 = ( wire1287 ) | ( wire1288 ) | ( wire1289 ) | ( wire1290 ) ;
 assign wire5154 = ( wire348 ) | ( wire1283 ) | ( wire1285 ) | ( wire1286 ) ;
 assign wire5155 = ( n_n1215 ) | ( wire1281 ) | ( wire1382 ) | ( wire1383 ) ;
 assign wire5156 = ( n_n1324 ) | ( wire1253 ) | ( wire4994  &  wire351 ) ;
 assign wire5157 = ( n_n1259 ) | ( n_n1193 ) | ( n_n1330 ) | ( n_n1267 ) ;
 assign wire5158 = ( wire342 ) | ( wire346 ) | ( wire1254 ) | ( wire1255 ) ;
 assign wire5159 = ( wire1256 ) | ( wire1257 ) | ( wire1350 ) | ( wire1351 ) ;
 assign wire5164 = ( wire5158 ) | ( wire5159 ) ;
 assign wire5165 = ( wire5150 ) | ( wire5151 ) | ( wire5152 ) | ( wire5153 ) ;
 assign wire5176 = ( n_n1082 ) | ( wire1235 ) | ( wire1487 ) ;
 assign wire5177 = ( n_n1188 ) | ( n_n1079 ) | ( n_n1070 ) | ( wire1417 ) ;
 assign wire5178 = ( n_n1163 ) | ( n_n1160 ) | ( n_n1215 ) | ( wire1281 ) ;
 assign wire5179 = ( n_n1204 ) | ( n_n1128 ) | ( wire236 ) | ( n_n1184 ) ;
 assign wire5180 = ( n_n1132 ) | ( n_n1130 ) | ( wire335 ) | ( n_n1173 ) ;
 assign wire5181 = ( n_n1181 ) | ( n_n1088 ) | ( n_n1216 ) | ( wire1234 ) ;
 assign wire5185 = ( wire306 ) | ( wire5176 ) | ( wire5181 ) ;
 assign wire5186 = ( wire5177 ) | ( wire5178 ) | ( wire5179 ) | ( wire5180 ) ;
 assign wire5191 = ( n_n93  &  n_n92  &  n_n94 ) | ( n_n92  &  n_n63  &  n_n94 ) ;
 assign wire5193 = ( n_n973 ) | ( n_n975 ) | ( wire1215 ) ;
 assign wire5194 = ( n_n967 ) | ( n_n966 ) | ( n_n987 ) | ( n_n984 ) ;
 assign wire5195 = ( n_n1021 ) | ( n_n956 ) | ( n_n1030 ) | ( n_n955 ) ;
 assign wire5196 = ( wire189 ) | ( n_n958 ) | ( n_n944 ) | ( n_n1060 ) ;
 assign wire5197 = ( n_n980 ) | ( n_n995 ) | ( n_n999 ) | ( n_n1004 ) ;
 assign wire5198 = ( n_n964 ) | ( n_n950 ) | ( wire5191 ) ;
 assign wire5202 = ( wire125 ) | ( wire5193 ) | ( wire5198 ) ;
 assign wire5203 = ( wire5194 ) | ( wire5195 ) | ( wire5196 ) | ( wire5197 ) ;
 assign wire5207 = ( n_n92  &  n_n82  &  n_n85 ) | ( n_n92  &  n_n95  &  n_n85 ) ;
 assign wire5208 = ( wire1197 ) | ( wire1489 ) | ( wire1490 ) ;
 assign wire5209 = ( n_n1281 ) | ( n_n1279 ) | ( wire1413 ) | ( wire1414 ) ;
 assign wire5210 = ( wire1287 ) | ( wire1288 ) | ( wire1291 ) | ( wire1292 ) ;
 assign wire5211 = ( wire348 ) | ( wire1283 ) | ( wire1285 ) | ( wire1286 ) ;
 assign wire5212 = ( n_n1254 ) | ( n_n1331 ) | ( wire1213 ) | ( wire1214 ) ;
 assign wire5213 = ( n_n1330 ) | ( wire323 ) | ( wire352 ) | ( wire357 ) ;
 assign wire5214 = ( wire1193 ) | ( wire1194 ) | ( wire5207 ) ;
 assign wire5227 = ( n_n1281 ) | ( n_n1279 ) | ( n_n1254 ) | ( n_n1331 ) ;
 assign wire5230 = ( n_n1074 ) | ( n_n1032 ) | ( n_n1294 ) | ( wire1179 ) ;
 assign wire5237 = ( n_n81  &  n_n78  &  n_n90 ) | ( n_n81  &  n_n82  &  n_n90 ) ;
 assign wire5239 = ( n_n1281 ) | ( n_n1279 ) | ( n_n1254 ) | ( n_n1331 ) ;
 assign wire5240 = ( n_n1109 ) | ( n_n1132 ) | ( n_n955 ) | ( wire135 ) ;
 assign wire5241 = ( n_n1330 ) | ( wire333 ) | ( _5553 ) ;
 assign wire5242 = ( n_n1324 ) | ( n_n1369 ) | ( n_n1286 ) | ( wire1175 ) ;
 assign wire5243 = ( n_n1259 ) | ( n_n1032 ) | ( n_n1169 ) | ( n_n942 ) ;
 assign wire5244 = ( n_n1128 ) | ( wire248 ) | ( wire5237 ) ;
 assign wire5257 = ( n_n1330 ) | ( wire189 ) | ( wire1527 ) ;
 assign wire5258 = ( n_n941 ) | ( wire333 ) | ( wire1173 ) | ( wire1177 ) ;
 assign wire5259 = ( n_n1324 ) | ( n_n1074 ) | ( wire1157 ) ;
 assign wire5295 = ( _69 ) | ( n_n91  &  n_n74  &  n_n83 ) ;
 assign wire5296 = ( wire1123 ) | ( wire1617 ) | ( wire1618 ) ;
 assign wire5297 = ( wire1485 ) | ( wire1486 ) | ( wire1535 ) | ( wire1536 ) ;
 assign wire5298 = ( wire323 ) | ( wire1142 ) | ( _5615 ) ;
 assign wire5299 = ( wire1144 ) | ( wire1145 ) | ( wire1533 ) | ( wire1534 ) ;
 assign wire5300 = ( wire252 ) | ( wire352 ) | ( n_n1176 ) | ( wire1106 ) ;
 assign wire5301 = ( wire246 ) | ( wire336 ) | ( n_n1217 ) | ( n_n1144 ) ;
 assign wire5302 = ( wire332 ) | ( wire333 ) | ( wire1107 ) | ( wire1108 ) ;
 assign wire5303 = ( wire1109 ) | ( wire1110 ) | ( wire1111 ) | ( wire1112 ) ;
 assign wire5304 = ( wire1113 ) | ( wire1114 ) | ( wire1115 ) | ( wire1116 ) ;
 assign wire5305 = ( wire1117 ) | ( wire1118 ) | ( wire1119 ) | ( wire1120 ) ;
 assign wire5326 = ( n_n1032 ) | ( n_n1040 ) | ( wire1085 ) ;
 assign wire5327 = ( n_n1036 ) | ( n_n1035 ) | ( _5724 ) ;
 assign wire5328 = ( wire203 ) | ( n_n1026 ) | ( wire4878 ) ;
 assign wire5329 = ( n_n1030 ) | ( n_n1060 ) | ( _5733 ) ;
 assign wire5330 = ( n_n1058 ) | ( n_n1048 ) | ( n_n999 ) | ( n_n1009 ) ;
 assign wire5331 = ( n_n1047 ) | ( n_n1001 ) | ( n_n1028 ) | ( n_n1018 ) ;
 assign wire5335 = ( wire286 ) | ( wire5326 ) | ( wire5331 ) ;
 assign wire5336 = ( wire5327 ) | ( wire5328 ) | ( wire5329 ) | ( wire5330 ) ;
 assign wire5340 = ( i_5_  &  (~ i_4_)  &  i_1_  &  i_2_ ) ;
 assign wire5342 = ( n_n97  &  n_n92 ) | ( n_n64  &  wire5340 ) ;
 assign wire5353 = ( n_n1125 ) | ( n_n1082 ) | ( wire1082 ) | ( wire1487 ) ;
 assign wire5354 = ( n_n1118 ) | ( n_n970 ) | ( n_n977 ) | ( wire1080 ) ;
 assign wire5355 = ( n_n990 ) | ( n_n993 ) | ( (~ i_8_)  &  wire70 ) ;
 assign wire5356 = ( n_n1081 ) | ( n_n1093 ) | ( n_n1074 ) | ( n_n1087 ) ;
 assign wire5357 = ( n_n968 ) | ( n_n958 ) | ( n_n974 ) | ( n_n973 ) ;
 assign wire5358 = ( n_n989 ) | ( n_n938 ) | ( n_n944 ) | ( n_n982 ) ;
 assign wire5359 = ( n_n967 ) | ( n_n956 ) | ( n_n1121 ) | ( wire236 ) ;
 assign wire5360 = ( wire319 ) | ( wire1046 ) | ( wire1048 ) | ( wire5342 ) ;
 assign wire5367 = ( wire232 ) | ( wire5360 ) ;
 assign wire5368 = ( wire257 ) | ( wire168 ) | ( wire291 ) | ( wire297 ) ;
 assign wire5379 = ( wire1024 ) | ( n_n83  &  _5783 ) ;
 assign wire5380 = ( n_n993 ) | ( wire1102 ) | ( _5786 ) ;
 assign wire5381 = ( n_n982 ) | ( n_n981 ) | ( wire1041 ) | ( wire1043 ) ;
 assign wire5382 = ( n_n969 ) | ( n_n1004 ) | ( n_n1001 ) | ( wire1039 ) ;
 assign wire5383 = ( n_n994 ) | ( n_n1025 ) | ( n_n976 ) | ( n_n987 ) ;
 assign wire5388 = ( wire292 ) | ( n_n882 ) | ( wire296 ) | ( wire5379 ) ;
 assign wire5389 = ( wire5380 ) | ( wire5381 ) | ( wire5382 ) | ( wire5383 ) ;
 assign wire5401 = ( n_n956 ) | ( n_n953 ) | ( n_n90  &  wire5012 ) ;
 assign wire5412 = ( _57 ) | ( n_n91  &  n_n92  &  n_n83 ) ;
 assign wire5413 = ( wire989 ) | ( wire1619 ) | ( wire1620 ) ;
 assign wire5414 = ( n_n1267 ) | ( wire1009 ) | ( wire1011 ) | ( wire1012 ) ;
 assign wire5415 = ( n_n1281 ) | ( wire346 ) | ( wire357 ) | ( wire248 ) ;
 assign wire5416 = ( wire326 ) | ( wire984 ) | ( wire985 ) | ( wire986 ) ;
 assign wire5421 = ( wire290 ) | ( wire289 ) | ( wire309 ) | ( wire5412 ) ;
 assign wire5422 = ( wire5413 ) | ( wire5414 ) | ( wire5415 ) | ( wire5416 ) ;
 assign wire5431 = ( wire963 ) | ( wire978 ) | ( wire979 ) ;
 assign wire5432 = ( wire1518 ) | ( wire1519 ) | ( wire982 ) | ( wire983 ) ;
 assign wire5433 = ( n_n1174 ) | ( n_n1177 ) | ( wire980 ) | ( wire981 ) ;
 assign wire5434 = ( wire252 ) | ( wire329 ) | ( n_n1176 ) | ( wire344 ) ;
 assign wire5435 = ( n_n1181 ) | ( wire243 ) | ( wire332 ) | ( n_n1170 ) ;
 assign wire5436 = ( wire959 ) | ( wire960 ) | ( wire961 ) | ( wire962 ) ;
 assign wire5440 = ( wire304 ) | ( wire5431 ) | ( wire5436 ) ;
 assign wire5441 = ( wire5432 ) | ( wire5433 ) | ( wire5434 ) | ( wire5435 ) ;
 assign wire5445 = ( i_7_  &  (~ i_8_)  &  (~ i_5_)  &  i_6_ ) ;
 assign wire5470 = ( wire334 ) | ( n_n1070 ) | ( wire946 ) | ( wire1313 ) ;
 assign wire5471 = ( n_n1105 ) | ( n_n1046 ) | ( n_n1047 ) | ( wire944 ) ;
 assign wire5472 = ( n_n1103 ) | ( n_n1095 ) | ( n_n1085 ) | ( wire942 ) ;
 assign wire5473 = ( n_n1077 ) | ( n_n1074 ) | ( n_n1048 ) | ( wire940 ) ;
 assign wire5474 = ( n_n1078 ) | ( n_n1032 ) | ( n_n1125 ) | ( wire906 ) ;
 assign wire5475 = ( wire319 ) | ( n_n1082 ) | ( n_n1045 ) | ( n_n1043 ) ;
 assign wire5476 = ( n_n1122 ) | ( n_n1036 ) | ( n_n1118 ) | ( n_n1030 ) ;
 assign wire5477 = ( n_n1083 ) | ( n_n1101 ) | ( wire355 ) | ( wire907 ) ;
 assign wire5478 = ( wire908 ) | ( wire909 ) | ( wire910 ) | ( wire911 ) ;
 assign wire5482 = ( wire5476 ) | ( wire5477 ) ;
 assign wire5483 = ( wire5470 ) | ( wire5471 ) | ( wire5478 ) ;
 assign wire5484 = ( wire5472 ) | ( wire5473 ) | ( wire5474 ) | ( wire5475 ) ;
 assign wire5502 = ( n_n1125 ) | ( n_n1163 ) | ( wire1082 ) ;
 assign wire5503 = ( n_n1118 ) | ( n_n1158 ) | ( n_n1146 ) | ( wire1080 ) ;
 assign wire5504 = ( n_n1108 ) | ( n_n1169 ) | ( wire897 ) | ( wire901 ) ;
 assign wire5505 = ( n_n1128 ) | ( wire356 ) | ( wire1386 ) | ( wire895 ) ;
 assign wire5506 = ( wire899 ) | ( wire900 ) | ( wire957 ) | ( wire958 ) ;
 assign wire5507 = ( n_n1153 ) | ( n_n1134 ) | ( n_n1132 ) | ( wire878 ) ;
 assign wire5508 = ( n_n1164 ) | ( n_n1145 ) | ( n_n1130 ) | ( wire246 ) ;
 assign wire5512 = ( wire5502 ) | ( wire5503 ) | ( wire5508 ) ;
 assign wire5513 = ( wire5504 ) | ( wire5505 ) | ( wire5506 ) | ( wire5507 ) ;
 assign wire5521 = ( n_n81  &  n_n83  &  n_n63 ) | ( n_n84  &  n_n83  &  n_n63 ) ;
 assign wire5523 = ( wire329 ) | ( n_n1286 ) | ( wire874 ) | ( wire1175 ) ;
 assign wire5524 = ( n_n1173 ) | ( n_n1170 ) | ( wire876 ) | ( wire877 ) ;
 assign wire5525 = ( wire872 ) | ( wire873 ) | ( wire982 ) | ( wire983 ) ;
 assign wire5526 = ( wire868 ) | ( wire869 ) | ( wire870 ) | ( wire871 ) ;
 assign wire5527 = ( n_n1172 ) | ( wire864 ) | ( wire866 ) | ( wire867 ) ;
 assign wire5528 = ( n_n1259 ) | ( wire314 ) | ( n_n1176 ) | ( n_n1184 ) ;
 assign wire5529 = ( wire326 ) | ( wire340 ) | ( _6026 ) ;
 assign wire5530 = ( wire833 ) | ( wire834 ) | ( wire835 ) | ( wire836 ) ;
 assign wire5537 = ( wire300 ) | ( wire5523 ) | ( wire5524 ) | ( wire5525 ) ;
 assign wire5538 = ( wire5526 ) | ( wire5527 ) | ( wire5528 ) | ( wire5529 ) ;
 assign wire5547 = ( _50 ) | ( n_n71  &  wire4873  &  _4879 ) ;
 assign wire5548 = ( n_n1001 ) | ( n_n1010 ) | ( wire812 ) ;
 assign wire5549 = ( n_n982 ) | ( n_n1019 ) | ( wire827 ) | ( wire1041 ) ;
 assign wire5550 = ( n_n1022 ) | ( n_n983 ) | ( n_n986 ) | ( wire825 ) ;
 assign wire5551 = ( n_n994 ) | ( n_n1025 ) | ( n_n1013 ) | ( n_n978 ) ;
 assign wire5556 = ( n_n882 ) | ( wire305 ) | ( wire286 ) | ( wire5547 ) ;
 assign wire5557 = ( wire5548 ) | ( wire5549 ) | ( wire5550 ) | ( wire5551 ) ;
 assign wire5569 = ( n_n1077 ) | ( n_n1074 ) | ( n_n1079 ) | ( n_n1070 ) ;
 assign wire5570 = ( wire809 ) | ( wire810 ) | ( wire807 ) | ( wire808 ) ;
 assign wire5571 = ( n_n1087 ) | ( n_n958 ) | ( n_n953 ) | ( wire805 ) ;
 assign wire5572 = ( n_n1052 ) | ( n_n951 ) | ( n_n950 ) | ( n_n1055 ) ;
 assign wire5573 = ( n_n1093 ) | ( n_n1057 ) | ( n_n956 ) | ( n_n1045 ) ;
 assign wire5574 = ( n_n1043 ) | ( n_n1101 ) | ( n_n1060 ) | ( n_n1100 ) ;
 assign wire5575 = ( n_n1046 ) | ( n_n954 ) | ( n_n969 ) | ( n_n939 ) ;
 assign wire5576 = ( n_n971 ) | ( n_n1035 ) | ( n_n1037 ) | ( n_n1058 ) ;
 assign wire5584 = ( wire168 ) | ( wire125 ) | ( _6088 ) ;
 assign wire5585 = ( wire298 ) | ( n_n421 ) | ( n_n241 ) | ( wire292 ) ;
 assign wire5586 = ( wire5569 ) | ( wire5570 ) | ( wire5571 ) | ( wire5572 ) ;
 assign wire5587 = ( wire5573 ) | ( wire5574 ) | ( wire5575 ) | ( wire5576 ) ;
 assign wire5597 = ( wire759 ) | ( wire1627 ) | ( wire1628 ) ;
 assign wire5598 = ( wire1155 ) | ( wire1156 ) | ( wire1289 ) | ( wire1290 ) ;
 assign wire5599 = ( wire1007 ) | ( wire1008 ) | ( wire980 ) | ( wire981 ) ;
 assign wire5600 = ( wire252 ) | ( n_n1279 ) | ( n_n1254 ) | ( wire348 ) ;
 assign wire5601 = ( wire755 ) | ( wire756 ) | ( wire757 ) | ( wire758 ) ;
 assign wire5605 = ( wire310 ) | ( wire309 ) | ( wire5601 ) ;
 assign wire5606 = ( wire5597 ) | ( wire5598 ) | ( wire5599 ) | ( wire5600 ) ;
 assign wire5613 = ( _41 ) | ( n_n97  &  n_n63  &  n_n77 ) ;
 assign wire5614 = ( n_n1036 ) | ( n_n1035 ) | ( wire736 ) ;
 assign wire5615 = ( n_n1020 ) | ( n_n993 ) | ( _6140 ) ;
 assign wire5616 = ( n_n982 ) | ( n_n1001 ) | ( n_n1019 ) | ( wire827 ) ;
 assign wire5617 = ( n_n1047 ) | ( n_n991 ) | ( n_n1013 ) | ( n_n1014 ) ;
 assign wire5622 = ( wire296 ) | ( wire167 ) | ( wire299 ) | ( wire5613 ) ;
 assign wire5623 = ( wire5614 ) | ( wire5615 ) | ( wire5616 ) | ( wire5617 ) ;
 assign wire5634 = ( _39 ) | ( n_n102  &  n_n85  &  _6161 ) ;
 assign wire5635 = ( n_n1103 ) | ( n_n1095 ) | ( wire1483 ) | ( wire1484 ) ;
 assign wire5636 = ( n_n958 ) | ( n_n951 ) | ( n_n950 ) | ( n_n953 ) ;
 assign wire5637 = ( n_n1057 ) | ( n_n944 ) | ( n_n939 ) | ( wire948 ) ;
 assign wire5638 = ( n_n947 ) | ( wire831 ) | ( n_n1068 ) | ( wire732 ) ;
 assign wire5639 = ( n_n956 ) | ( n_n1100 ) | ( n_n955 ) | ( wire1499 ) ;
 assign wire5640 = ( n_n969 ) | ( wire957 ) | ( wire958 ) | ( wire1039 ) ;
 assign wire5641 = ( n_n1134 ) | ( n_n962 ) | ( n_n964 ) | ( n_n1132 ) ;
 assign wire5642 = ( n_n1121 ) | ( wire236 ) | ( n_n1122 ) | ( wire734 ) ;
 assign wire5643 = ( n_n949 ) | ( n_n954 ) | ( n_n1101 ) | ( n_n1058 ) ;
 assign wire5644 = ( wire345 ) | ( n_n978 ) | ( n_n1079 ) | ( n_n977 ) ;
 assign wire5645 = ( n_n959 ) | ( n_n957 ) | ( wire696 ) | ( wire697 ) ;
 assign wire5652 = ( n_n941 ) | ( n_n943 ) | ( wire125 ) | ( wire5645 ) ;
 assign wire5653 = ( wire287 ) | ( wire5634 ) | ( wire5635 ) | ( wire5636 ) ;
 assign wire5654 = ( wire5637 ) | ( wire5638 ) | ( wire5639 ) | ( wire5640 ) ;
 assign wire5655 = ( wire5641 ) | ( wire5642 ) | ( wire5643 ) | ( wire5644 ) ;
 assign wire5662 = ( (~ i_5_)  &  i_3_ ) ;
 assign wire5668 = ( n_n91  &  n_n99  &  n_n94 ) | ( n_n91  &  n_n94  &  wire5662 ) ;
 assign wire5671 = ( n_n1204 ) | ( wire1531 ) | ( wire692 ) | ( wire693 ) ;
 assign wire5672 = ( n_n1163 ) | ( n_n1160 ) | ( wire1142 ) | ( wire1143 ) ;
 assign wire5673 = ( n_n1158 ) | ( n_n1216 ) | ( n_n1146 ) | ( wire690 ) ;
 assign wire5674 = ( wire235 ) | ( n_n1193 ) | ( wire342 ) | ( wire666 ) ;
 assign wire5675 = ( n_n1169 ) | ( n_n1184 ) | ( n_n1145 ) | ( n_n1188 ) ;
 assign wire5676 = ( wire668 ) | ( wire669 ) | ( wire5668 ) ;
 assign wire5681 = ( n_n554 ) | ( wire670 ) | ( wire671 ) | ( wire5676 ) ;
 assign wire5682 = ( n_n211 ) | ( wire5671 ) | ( wire5672 ) | ( wire5673 ) ;
 assign wire5698 = ( wire332 ) | ( wire664 ) | ( wire1627 ) | ( wire1628 ) ;
 assign wire5699 = ( wire1153 ) | ( wire1154 ) | ( wire662 ) | ( wire663 ) ;
 assign wire5700 = ( wire235 ) | ( n_n1259 ) | ( n_n1312 ) | ( wire344 ) ;
 assign wire5701 = ( wire343 ) | ( n_n1215 ) | ( wire350 ) | ( wire641 ) ;
 assign wire5702 = ( wire642 ) | ( wire643 ) | ( wire644 ) | ( wire645 ) ;
 assign wire5703 = ( wire646 ) | ( wire647 ) | ( wire648 ) | ( wire649 ) ;
 assign wire5707 = ( wire289 ) | ( wire5698 ) | ( wire5703 ) ;
 assign wire5708 = ( wire5699 ) | ( wire5700 ) | ( wire5701 ) | ( wire5702 ) ;
 assign wire5719 = ( n_n1185 ) | ( wire321 ) | ( n_n1193 ) | ( wire336 ) ;
 assign wire5720 = ( wire876 ) | ( wire877 ) | ( wire1144 ) | ( wire1145 ) ;
 assign wire5721 = ( wire870 ) | ( wire871 ) | ( wire872 ) | ( wire873 ) ;
 assign wire5722 = ( n_n1172 ) | ( wire864 ) | ( wire1507 ) | ( wire1508 ) ;
 assign wire5723 = ( n_n1134 ) | ( n_n1331 ) | ( wire248 ) | ( n_n1147 ) ;
 assign wire5724 = ( n_n1181 ) | ( wire246 ) | ( n_n1144 ) | ( wire333 ) ;
 assign wire5725 = ( n_n1160 ) | ( wire617 ) | ( wire618 ) | ( wire619 ) ;
 assign wire5730 = ( wire295 ) | ( wire620 ) | ( wire621 ) | ( wire5725 ) ;
 assign wire5731 = ( wire5719 ) | ( wire5720 ) | ( wire5721 ) | ( wire5722 ) ;
 assign wire5741 = ( n_n1014 ) | ( n_n1018 ) | ( n_n1019 ) | ( wire827 ) ;
 assign wire5742 = ( n_n1037 ) | ( n_n1009 ) | ( n_n1028 ) | ( wire611 ) ;
 assign wire5743 = ( n_n1021 ) | ( n_n1022 ) | ( n_n994 ) | ( n_n990 ) ;
 assign wire5744 = ( n_n1002 ) | ( n_n1006 ) | ( n_n1010 ) | ( wire596 ) ;
 assign wire5748 = ( wire302 ) | ( n_n296 ) | ( wire5744 ) ;
 assign wire5749 = ( wire305 ) | ( wire5741 ) | ( wire5742 ) | ( wire5743 ) ;
 assign wire5750 = ( (~ i_7_)  &  i_5_  &  i_6_  &  (~ i_4_) ) ;
 assign wire5756 = ( n_n58  &  n_n84  &  n_n85 ) | ( n_n84  &  n_n95  &  n_n85 ) ;
 assign wire5758 = ( wire562 ) | ( wire245  &  wire5750 ) ;
 assign wire5759 = ( n_n970 ) | ( n_n1055 ) | ( n_n1085 ) | ( n_n977 ) ;
 assign wire5760 = ( wire334 ) | ( n_n1070 ) | ( wire946 ) | ( wire1313 ) ;
 assign wire5761 = ( n_n942 ) | ( n_n1087 ) | ( n_n938 ) | ( wire805 ) ;
 assign wire5762 = ( n_n1057 ) | ( wire103 ) | ( wire948 ) ;
 assign wire5763 = ( n_n1108 ) | ( n_n944 ) | ( n_n939 ) | ( wire897 ) ;
 assign wire5764 = ( n_n947 ) | ( wire831 ) | ( n_n1068 ) | ( wire732 ) ;
 assign wire5765 = ( n_n1077 ) | ( n_n1081 ) | ( n_n1120 ) | ( n_n1122 ) ;
 assign wire5766 = ( n_n1091 ) | ( n_n982 ) | ( wire236 ) | ( n_n1083 ) ;
 assign wire5767 = ( n_n971 ) | ( n_n1132 ) | ( n_n1048 ) | ( n_n980 ) ;
 assign wire5768 = ( n_n983 ) | ( n_n1117 ) | ( wire5756 ) ;
 assign wire5775 = ( wire291 ) | ( wire5758 ) | ( wire5759 ) | ( wire5760 ) ;
 assign wire5776 = ( wire5761 ) | ( wire5762 ) | ( wire5763 ) | ( wire5764 ) ;
 assign wire5777 = ( wire5765 ) | ( wire5766 ) | ( wire5767 ) | ( wire5768 ) ;
 assign wire5787 = ( n_n1021 ) | ( n_n1030 ) | ( n_n1014 ) | ( n_n1018 ) ;
 assign wire5788 = ( n_n1046 ) | ( n_n1009 ) | ( _6353 ) ;
 assign wire5789 = ( _6358 ) | ( _6359 ) ;
 assign wire5790 = ( n_n1045 ) | ( n_n1037 ) | ( n_n1013 ) | ( n_n1028 ) ;
 assign wire5791 = ( n_n1010 ) | ( n_n1020 ) | ( wire249 ) | ( n_n1026 ) ;
 assign wire5795 = ( wire299 ) | ( wire286 ) | ( wire5791 ) ;
 assign wire5796 = ( wire5787 ) | ( wire5788 ) | ( wire5789 ) | ( wire5790 ) ;
 assign wire5803 = ( n_n959 ) | ( n_n970 ) | ( n_n977 ) ;
 assign wire5804 = ( n_n958 ) | ( wire103 ) | ( n_n953 ) ;
 assign wire5805 = ( n_n954 ) | ( n_n952 ) | ( n_n971 ) | ( n_n976 ) ;
 assign wire5806 = ( n_n973 ) | ( n_n975 ) | ( n_n987 ) | ( n_n984 ) ;
 assign wire5807 = ( n_n981 ) | ( n_n994 ) | ( n_n978 ) | ( wire1043 ) ;
 assign wire5808 = ( n_n968 ) | ( n_n989 ) | ( n_n956 ) | ( wire532 ) ;
 assign wire5809 = ( n_n969 ) | ( n_n995 ) | ( n_n999 ) | ( n_n1004 ) ;
 assign wire5815 = ( wire5807 ) | ( wire5808 ) ;
 assign wire5816 = ( wire168 ) | ( n_n990 ) | ( n_n993 ) | ( wire5809 ) ;
 assign wire5817 = ( wire303 ) | ( n_n652 ) | ( wire296 ) | ( wire167 ) ;
 assign wire5818 = ( wire5803 ) | ( wire5804 ) | ( wire5805 ) | ( wire5806 ) ;
 assign wire5833 = ( n_n91  &  n_n103  &  n_n92 ) | ( n_n91  &  n_n97  &  n_n92 ) ;
 assign wire5836 = ( n_n1077 ) | ( n_n1105 ) | ( n_n1074 ) | ( wire944 ) ;
 assign wire5837 = ( n_n1055 ) | ( wire805 ) | ( _6430 ) ;
 assign wire5838 = ( n_n1108 ) | ( wire897 ) | ( wire899 ) | ( wire900 ) ;
 assign wire5839 = ( n_n1092 ) | ( n_n1091 ) | ( n_n1109 ) | ( wire355 ) ;
 assign wire5840 = ( n_n1100 ) | ( n_n1117 ) | ( wire5833 ) ;
 assign wire5841 = ( n_n1047 ) | ( n_n1068 ) | ( wire507 ) | ( wire508 ) ;
 assign wire5845 = ( n_n421 ) | ( wire5836 ) | ( wire5841 ) ;
 assign wire5846 = ( wire5837 ) | ( wire5838 ) | ( wire5839 ) | ( wire5840 ) ;
 assign wire5848 = ( n_n78  &  n_n84  &  n_n90 ) | ( n_n78  &  n_n92  &  n_n90 ) ;
 assign wire5858 = ( n_n1188 ) | ( wire1417 ) | ( wire1623 ) | ( wire1624 ) ;
 assign wire5859 = ( wire343 ) | ( wire1213 ) | ( wire1214 ) | ( wire1411 ) ;
 assign wire5860 = ( n_n1169 ) | ( wire692 ) | ( wire693 ) | ( wire901 ) ;
 assign wire5861 = ( wire329 ) | ( wire874 ) | ( wire978 ) | ( wire979 ) ;
 assign wire5862 = ( n_n1286 ) | ( n_n1283 ) | ( wire5848 ) ;
 assign wire5863 = ( n_n1156 ) | ( n_n1177 ) | ( wire335 ) | ( wire340 ) ;
 assign wire5864 = ( wire344 ) | ( wire475 ) | ( wire476 ) | ( wire477 ) ;
 assign wire5865 = ( wire478 ) | ( wire479 ) | ( wire480 ) | ( wire481 ) ;
 assign wire5866 = ( wire482 ) | ( wire483 ) | ( wire484 ) | ( wire485 ) ;
 assign wire5871 = ( wire5865 ) | ( wire5866 ) ;
 assign wire5872 = ( wire301 ) | ( wire5858 ) | ( wire5859 ) | ( wire5860 ) ;
 assign wire5873 = ( wire5861 ) | ( wire5862 ) | ( wire5863 ) | ( wire5864 ) ;
 assign wire5886 = ( wire356 ) | ( n_n1085 ) | ( wire942 ) ;
 assign wire5887 = ( n_n1120 ) | ( n_n1122 ) | ( wire807 ) | ( wire808 ) ;
 assign wire5888 = ( n_n1014 ) | ( n_n1018 ) | ( n_n1019 ) | ( wire827 ) ;
 assign wire5889 = ( n_n1092 ) | ( n_n1074 ) | ( n_n1045 ) | ( n_n1060 ) ;
 assign wire5890 = ( n_n1145 ) | ( n_n1048 ) | ( n_n1147 ) | ( n_n1009 ) ;
 assign wire5891 = ( n_n1144 ) | ( n_n1013 ) | ( n_n1146 ) | ( n_n1010 ) ;
 assign wire5892 = ( n_n1108 ) | ( n_n1105 ) | ( wire334 ) | ( n_n1020 ) ;
 assign wire5896 = ( wire5886 ) | ( wire5887 ) | ( wire5892 ) ;
 assign wire5897 = ( wire5888 ) | ( wire5889 ) | ( wire5890 ) | ( wire5891 ) ;
 assign wire5901 = ( n_n980 ) | ( n_n981 ) | ( n_n999 ) | ( wire615 ) ;
 assign wire5902 = ( wire103 ) | ( n_n994 ) | ( n_n991 ) | ( n_n984 ) ;
 assign wire5905 = ( n_n78  &  n_n103  &  n_n84 ) | ( n_n78  &  n_n100  &  n_n84 ) ;
 assign wire5907 = ( n_n1174 ) | ( n_n1177 ) | ( wire876 ) | ( wire877 ) ;
 assign wire5908 = ( n_n1216 ) | ( wire469 ) | ( wire690 ) | ( wire5905 ) ;
 assign wire5919 = ( wire346 ) | ( n_n1163 ) | ( n_n1160 ) | ( wire1415 ) ;
 assign wire5920 = ( n_n1169 ) | ( wire467 ) | ( wire468 ) | ( wire901 ) ;
 assign wire5921 = ( wire332 ) | ( wire664 ) | ( wire1011 ) | ( wire1012 ) ;
 assign wire5922 = ( n_n1267 ) | ( wire662 ) | ( wire663 ) | ( wire1009 ) ;
 assign wire5923 = ( wire321 ) | ( n_n1173 ) | ( wire336 ) | ( n_n1170 ) ;
 assign wire5924 = ( wire235 ) | ( n_n1286 ) | ( n_n971 ) | ( n_n1158 ) ;
 assign wire5925 = ( n_n1312 ) | ( n_n970 ) | ( wire430 ) | ( wire431 ) ;
 assign wire5926 = ( wire432 ) | ( wire433 ) | ( wire434 ) | ( wire435 ) ;
 assign wire5927 = ( wire436 ) | ( wire437 ) | ( wire438 ) | ( wire439 ) ;
 assign wire5936 = ( wire5921 ) | ( wire5922 ) | ( wire5923 ) | ( wire5924 ) ;
 assign wire5937 = ( wire5901 ) | ( wire5902 ) | ( wire5925 ) | ( wire5926 ) ;
 assign wire5947 = ( _19 ) | ( n_n99  &  n_n95  &  n_n85 ) ;
 assign wire5948 = ( n_n1048 ) | ( n_n1085 ) | ( wire940 ) ;
 assign wire5949 = ( n_n1021 ) | ( n_n1030 ) | ( n_n1014 ) | ( n_n1018 ) ;
 assign wire5950 = ( n_n1043 ) | ( n_n1009 ) | ( wire559 ) | ( wire611 ) ;
 assign wire5951 = ( n_n1039 ) | ( n_n1037 ) | ( n_n1028 ) | ( wire413 ) ;
 assign wire5952 = ( n_n1057 ) | ( n_n1087 ) | ( n_n1083 ) | ( n_n1013 ) ;
 assign wire5957 = ( wire167 ) | ( wire287 ) | ( wire5947 ) | ( wire5948 ) ;
 assign wire5958 = ( wire5949 ) | ( wire5950 ) | ( wire5951 ) | ( wire5952 ) ;
 assign wire5971 = ( n_n1188 ) | ( wire395 ) | ( wire1417 ) ;
 assign wire5972 = ( n_n1185 ) | ( n_n1193 ) | ( wire1291 ) | ( wire1292 ) ;
 assign wire5973 = ( wire467 ) | ( wire468 ) | ( wire1380 ) | ( wire1381 ) ;
 assign wire5974 = ( n_n1297 ) | ( wire314 ) | ( wire866 ) | ( wire867 ) ;
 assign wire5975 = ( wire243 ) | ( wire323 ) | ( n_n1294 ) | ( n_n1283 ) ;
 assign wire5976 = ( n_n1215 ) | ( wire350 ) | ( wire348 ) | ( wire382 ) ;
 assign wire5977 = ( wire383 ) | ( wire384 ) | ( wire385 ) | ( wire386 ) ;
 assign wire5978 = ( wire387 ) | ( wire388 ) | ( wire389 ) | ( wire390 ) ;
 assign wire5979 = ( wire391 ) | ( wire392 ) | ( wire393 ) | ( wire394 ) ;
 assign wire5989 = ( n_n100  &  n_n74  &  n_n95 ) | ( n_n74  &  n_n95  &  n_n83 ) ;
 assign wire5995 = ( (~ i_7_)  &  (~ i_8_)  &  (~ i_6_)  &  i_2_ ) ;
 assign wire6006 = ( n_n77  &  wire5995 ) | ( n_n101  &  n_n77  &  n_n85 ) ;
 assign wire6007 = ( n_n970 ) | ( n_n977 ) | ( wire165 ) ;
 assign wire6008 = ( n_n1105 ) | ( n_n958 ) | ( n_n953 ) | ( wire944 ) ;
 assign wire6009 = ( n_n1120 ) | ( n_n944 ) | ( n_n1122 ) | ( n_n939 ) ;
 assign wire6010 = ( n_n1109 ) | ( wire1348 ) | ( n_n1100 ) | ( wire1499 ) ;
 assign wire6011 = ( n_n1092 ) | ( n_n1128 ) | ( wire60 ) | ( wire895 ) ;
 assign wire6012 = ( wire251 ) | ( wire321 ) | ( n_n1176 ) | ( n_n974 ) ;
 assign wire6013 = ( n_n1156 ) | ( n_n969 ) | ( n_n1184 ) | ( n_n1147 ) ;
 assign wire6014 = ( n_n1164 ) | ( n_n962 ) | ( n_n941 ) | ( n_n975 ) ;
 assign wire6015 = ( n_n966 ) | ( n_n1173 ) | ( n_n1088 ) | ( wire246 ) ;
 assign wire6016 = ( wire336 ) | ( wire69 ) | ( wire6006 ) ;
 assign wire6023 = ( wire125 ) | ( n_n652 ) | ( wire6007 ) | ( wire6008 ) ;
 assign _19 = ( n_n81  &  n_n93  &  n_n100 ) ;
 assign _39 = ( i_7_  &  (~ i_8_)  &  n_n84  &  n_n97 ) ;
 assign _41 = ( n_n96  &  n_n82  &  n_n85 ) ;
 assign _46 = ( i_8_  &  i_6_  &  n_n103  &  n_n77 ) ;
 assign _48 = ( n_n93  &  n_n96  &  n_n94 ) ;
 assign _50 = ( (~ i_7_)  &  (~ i_8_)  &  n_n85  &  n_n76 ) ;
 assign _57 = ( n_n93  &  n_n77  &  n_n94 ) ;
 assign _69 = ( n_n93  &  n_n100  &  n_n84 ) ;
 assign _83 = ( n_n81  &  n_n93  &  n_n100 ) ;
 assign _4857 = ( i_7_  &  i_8_  &  i_2_  &  i_0_ ) ;
 assign _4863 = ( i_7_  &  i_8_  &  (~ i_6_)  &  (~ i_3_) ) ;
 assign _4865 = ( n_n83  &  _4863 ) | ( n_n99  &  n_n95  &  n_n83 ) ;
 assign _4879 = ( (~ i_8_)  &  i_7_ ) ;
 assign _4881 = ( (~ i_7_)  &  (~ i_8_)  &  (~ i_5_)  &  i_6_ ) ;
 assign _4906 = ( i_7_  &  (~ i_8_)  &  (~ i_6_)  &  n_n74 ) ;
 assign _5158 = ( (~ i_3_)  &  (~ i_1_)  &  (~ i_0_) ) ;
 assign _5183 = ( n_n91  &  n_n103  &  n_n92 ) | ( n_n91  &  n_n97  &  n_n92 ) ;
 assign _5226 = ( (~ i_1_)  &  i_2_  &  (~ i_0_) ) ;
 assign _5523 = ( wire4994  &  _5158 ) | ( wire5012  &  _5226 ) ;
 assign _5553 = ( n_n92  &  n_n82  &  n_n90 ) | ( n_n92  &  n_n82  &  n_n94 ) ;
 assign _5615 = ( n_n58  &  n_n100  &  n_n84 ) | ( n_n100  &  n_n84  &  n_n95 ) ;
 assign _5644 = ( i_7_  &  (~ i_8_)  &  (~ i_1_)  &  i_2_ ) ;
 assign _5645 = ( i_5_  &  (~ i_6_)  &  (~ i_3_)  &  i_4_ ) ;
 assign _5668 = ( (~ i_7_)  &  i_8_  &  i_5_  &  (~ i_4_) ) ;
 assign _5724 = ( n_n83  &  _4863 ) | ( n_n99  &  n_n95  &  n_n83 ) ;
 assign _5729 = ( (~ i_5_)  &  (~ i_6_)  &  i_4_ ) ;
 assign _5732 = ( i_1_  &  (~ i_2_)  &  i_0_ ) ;
 assign _5733 = ( wire5318  &  _5729 ) | ( wire5319  &  _5732 ) ;
 assign _5783 = ( i_7_  &  i_8_  &  (~ i_6_)  &  i_3_ ) ;
 assign _5786 = ( n_n74  &  n_n95  &  n_n83 ) | ( n_n74  &  n_n95  &  n_n94 ) ;
 assign _5980 = ( wire839 ) | ( wire840 ) | ( wire5521 ) | ( wire5530 ) ;
 assign _6026 = ( n_n101  &  n_n103  &  n_n74 ) | ( n_n101  &  n_n100  &  n_n74 ) ;
 assign _6079 = ( (~ i_1_)  &  i_2_  &  i_0_ ) ;
 assign _6088 = ( n_n943 ) | ( n_n1059 ) | ( _46 ) | ( _48 ) ;
 assign _6101 = ( wire5537 ) | ( wire5586 ) | ( wire5587 ) | ( _5980 ) ;
 assign _6140 = ( n_n74  &  n_n82  &  n_n83 ) | ( n_n74  &  n_n95  &  n_n83 ) ;
 assign _6161 = ( (~ i_6_)  &  (~ i_7_) ) ;
 assign _6190 = ( wire5675 ) | ( wire5674 ) ;
 assign _6228 = ( wire5654 ) | ( wire5655 ) | ( wire5681 ) | ( _6190 ) ;
 assign _6248 = ( wire5724 ) | ( wire5723 ) ;
 assign _6319 = ( i_7_  &  i_8_  &  (~ i_6_)  &  i_3_ ) ;
 assign _6325 = ( i_6_  &  i_7_ ) ;
 assign _6345 = ( wire5730 ) | ( wire5776 ) | ( wire5777 ) | ( _6248 ) ;
 assign _6353 = ( n_n83  &  _4881 ) | ( n_n96  &  n_n83  &  _6325 ) ;
 assign _6357 = ( i_1_  &  i_2_  &  (~ i_0_) ) ;
 assign _6358 = ( wire5544  &  _6079 ) | ( wire5783  &  _6357 ) ;
 assign _6359 = ( n_n58  &  n_n102  &  n_n85 ) | ( n_n91  &  n_n102  &  n_n85 ) ;
 assign _6377 = ( i_7_  &  i_8_  &  (~ i_6_) ) ;
 assign _6430 = ( n_n81  &  n_n63  &  n_n94 ) | ( n_n74  &  n_n63  &  n_n94 ) ;


endmodule

